magic
tech sky130A
timestamp 1756577777
<< metal1 >>
rect 12410 10500 12430 10520
<< via1 >>
rect 13280 10055 13310 10085
<< metal2 >>
rect 11685 16840 11725 16845
rect 11685 16811 11690 16840
rect 11720 16811 11725 16840
rect 11685 16799 11725 16811
rect 11685 16770 11690 16799
rect 11720 16770 11725 16799
rect 11685 16765 11725 16770
rect 13275 10085 13315 10090
rect 13275 10055 13280 10085
rect 13310 10055 13315 10085
rect 13275 9765 13315 10055
rect 13255 9755 13335 9765
rect 13255 9725 13280 9755
rect 13310 9725 13335 9755
rect 13255 9715 13335 9725
<< via2 >>
rect 11690 16811 11720 16840
rect 11690 16770 11720 16799
rect 13280 9725 13310 9755
<< metal3 >>
rect 400 18210 11505 18215
rect 400 18170 405 18210
rect 445 18170 455 18210
rect 495 18170 505 18210
rect 545 18170 555 18210
rect 595 18170 11460 18210
rect 11500 18170 11505 18210
rect 400 18160 11505 18170
rect 400 18120 405 18160
rect 445 18120 455 18160
rect 495 18120 505 18160
rect 545 18120 555 18160
rect 595 18120 11460 18160
rect 11500 18120 11505 18160
rect 400 18110 11505 18120
rect 400 18070 405 18110
rect 445 18070 455 18110
rect 495 18070 505 18110
rect 545 18070 555 18110
rect 595 18070 11460 18110
rect 11500 18070 11505 18110
rect 400 18060 11505 18070
rect 400 18020 405 18060
rect 445 18020 455 18060
rect 495 18020 505 18060
rect 545 18020 555 18060
rect 595 18020 11460 18060
rect 11500 18020 11505 18060
rect 400 18015 11505 18020
rect 100 17795 12090 17800
rect 100 17755 105 17795
rect 145 17755 155 17795
rect 195 17755 205 17795
rect 245 17755 255 17795
rect 295 17755 12045 17795
rect 12085 17755 12090 17795
rect 100 17745 12090 17755
rect 100 17705 105 17745
rect 145 17705 155 17745
rect 195 17705 205 17745
rect 245 17705 255 17745
rect 295 17705 12045 17745
rect 12085 17705 12090 17745
rect 100 17695 12090 17705
rect 100 17655 105 17695
rect 145 17655 155 17695
rect 195 17655 205 17695
rect 245 17655 255 17695
rect 295 17655 12045 17695
rect 12085 17655 12090 17695
rect 100 17645 12090 17655
rect 100 17605 105 17645
rect 145 17605 155 17645
rect 195 17605 205 17645
rect 245 17605 255 17645
rect 295 17605 12045 17645
rect 12085 17605 12090 17645
rect 100 17600 12090 17605
rect 11685 16840 15265 16845
rect 11685 16811 11690 16840
rect 11720 16825 15265 16840
rect 11720 16811 15205 16825
rect 11685 16799 15205 16811
rect 11685 16770 11690 16799
rect 11720 16785 15205 16799
rect 15245 16785 15265 16825
rect 11720 16770 15265 16785
rect 11685 16765 15265 16770
rect 13255 9760 13335 9765
rect 13255 9720 13275 9760
rect 13315 9720 13335 9760
rect 13255 9715 13335 9720
<< via3 >>
rect 405 18170 445 18210
rect 455 18170 495 18210
rect 505 18170 545 18210
rect 555 18170 595 18210
rect 11460 18170 11500 18210
rect 405 18120 445 18160
rect 455 18120 495 18160
rect 505 18120 545 18160
rect 555 18120 595 18160
rect 11460 18120 11500 18160
rect 405 18070 445 18110
rect 455 18070 495 18110
rect 505 18070 545 18110
rect 555 18070 595 18110
rect 11460 18070 11500 18110
rect 405 18020 445 18060
rect 455 18020 495 18060
rect 505 18020 545 18060
rect 555 18020 595 18060
rect 11460 18020 11500 18060
rect 105 17755 145 17795
rect 155 17755 195 17795
rect 205 17755 245 17795
rect 255 17755 295 17795
rect 12045 17755 12085 17795
rect 105 17705 145 17745
rect 155 17705 195 17745
rect 205 17705 245 17745
rect 255 17705 295 17745
rect 12045 17705 12085 17745
rect 105 17655 145 17695
rect 155 17655 195 17695
rect 205 17655 245 17695
rect 255 17655 295 17695
rect 12045 17655 12085 17695
rect 105 17605 145 17645
rect 155 17605 195 17645
rect 205 17605 245 17645
rect 255 17605 295 17645
rect 12045 17605 12085 17645
rect 15205 16785 15245 16825
rect 13275 9755 13315 9760
rect 13275 9725 13280 9755
rect 13280 9725 13310 9755
rect 13310 9725 13315 9755
rect 13275 9720 13315 9725
<< metal4 >>
rect 100 17795 300 22076
rect 400 18210 600 22076
rect 400 18170 405 18210
rect 445 18170 455 18210
rect 495 18170 505 18210
rect 545 18170 555 18210
rect 595 18170 600 18210
rect 400 18160 600 18170
rect 400 18120 405 18160
rect 445 18120 455 18160
rect 495 18120 505 18160
rect 545 18120 555 18160
rect 595 18120 600 18160
rect 400 18110 600 18120
rect 400 18070 405 18110
rect 445 18070 455 18110
rect 495 18070 505 18110
rect 545 18070 555 18110
rect 595 18070 600 18110
rect 400 18060 600 18070
rect 400 18020 405 18060
rect 445 18020 455 18060
rect 495 18020 505 18060
rect 545 18020 555 18060
rect 595 18020 600 18060
rect 400 17800 600 18020
rect 11455 18210 11505 18215
rect 11455 18170 11460 18210
rect 11500 18170 11505 18210
rect 11455 18160 11505 18170
rect 11455 18120 11460 18160
rect 11500 18120 11505 18160
rect 11455 18110 11505 18120
rect 11455 18070 11460 18110
rect 11500 18070 11505 18110
rect 11455 18060 11505 18070
rect 11455 18020 11460 18060
rect 11500 18020 11505 18060
rect 100 17755 105 17795
rect 145 17755 155 17795
rect 195 17755 205 17795
rect 245 17755 255 17795
rect 295 17755 300 17795
rect 100 17745 300 17755
rect 100 17705 105 17745
rect 145 17705 155 17745
rect 195 17705 205 17745
rect 245 17705 255 17745
rect 295 17705 300 17745
rect 100 17695 300 17705
rect 100 17655 105 17695
rect 145 17655 155 17695
rect 195 17655 205 17695
rect 245 17655 255 17695
rect 295 17655 300 17695
rect 100 17645 300 17655
rect 100 17605 105 17645
rect 145 17605 155 17645
rect 195 17605 205 17645
rect 245 17605 255 17645
rect 295 17605 300 17645
rect 100 500 300 17605
rect 400 500 600 17600
rect 11455 16260 11505 18020
rect 12040 17795 12090 17800
rect 12040 17755 12045 17795
rect 12085 17755 12090 17795
rect 12040 17745 12090 17755
rect 12040 17705 12045 17745
rect 12085 17705 12090 17745
rect 12040 17695 12090 17705
rect 12040 17655 12045 17695
rect 12085 17655 12090 17695
rect 12040 17645 12090 17655
rect 12040 17605 12045 17645
rect 12085 17605 12090 17645
rect 12040 16410 12090 17605
rect 15185 16825 15265 16845
rect 15185 16785 15205 16825
rect 15245 16785 15265 16825
rect 13255 9760 13335 9765
rect 13255 9720 13275 9760
rect 13315 9720 13335 9760
rect 13255 100 13335 9720
rect 15185 100 15265 16785
rect 13249 0 13339 100
rect 15181 0 15271 100
use pll_bgr_magic_flat  pll_bgr_magic_flat_0
timestamp 1756577646
transform 0 -1 13930 -1 0 17120
box 0 0 15790 7605
<< labels >>
flabel metal4 s 15181 0 15271 100 0 FreeSans 480 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 13249 0 13339 100 0 FreeSans 480 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal1 12420 10500 12420 10500 5 FreeSans 800 0 0 -400 V_CONT
flabel metal4 100 500 300 22076 1 FreeSans 200 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 400 500 600 22076 1 FreeSans 200 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16100 22576
<< end >>
