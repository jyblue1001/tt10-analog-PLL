* PEX produced on Wed Sep  3 11:51:33 AM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from project_3.ext - technology: sky130A

.subckt project_3 ua[0] ua[1] VDPWR VGND
X0 a_13750_11850.t7 a_10354_16286.t6 a_14040_12560.t8 VGND.t212 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X1 VGND.t42 I_IN.t15 I_IN.t16 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X2 a_10710_11860.t11 a_8454_18026.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3 VGND.t176 VDPWR.t426 a_11880_10030.t9 VGND.t175 sky130_fd_pr__nfet_01v8 ad=1.01 pd=6.15 as=1 ps=5.8 w=2.5 l=5
X4 VDPWR.t114 a_21100_10960.t5 a_17450_6090.t7 VDPWR.t113 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X5 VDPWR.t23 ua[1].t2 a_21810_3370.t2 VDPWR.t22 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X6 a_17290_6090.t1 a_16900_6090.t2 VDPWR.t202 VDPWR.t186 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X7 a_16510_6090.t1 a_13440_6060.t3 VDPWR.t99 VDPWR.t98 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X8 a_16630_3080.t2 a_16740_3080.t3 VGND.t52 VGND.t51 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X9 a_19440_11540.t8 a_19440_11540.t7 a_19440_11540.t8 VDPWR.t373 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X10 a_10710_11860.t12 a_8454_18026.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X11 VDPWR.t31 a_18230_3320.t2 a_17820_3240.t0 VDPWR.t30 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X12 VDPWR.t80 PFET_GATE.t10 I_IN.t5 VDPWR.t79 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X13 a_20510_3370.t0 a_21210_3400.t2 VGND.t107 VGND.t106 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X14 a_11880_10030.t14 VDPWR.t376 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X15 a_19670_10930.t4 a_19670_10930.t3 VGND.t309 VGND.t308 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X16 PFET_GATE.t7 VDPWR.t427 VGND.t179 VGND.t178 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X17 a_10710_11860.t13 a_8454_18026.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X18 a_13360_6510.t0 ua[0].t0 VDPWR.t72 VDPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X19 VDPWR.t66 a_13880_11590.t14 a_13880_11590.t15 VDPWR.t65 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X20 VDPWR.t282 a_10710_11860.t14 PFET_GATE.t6 VDPWR.t281 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X21 ua[1].t0 a_23830_2840.t2 a_24238_3560.t0 VDPWR.t181 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.16
X22 a_10740_13170.t4 a_9573_16817.t7 a_10840_11590.t1 VGND.t117 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X23 a_13750_11850.t11 a_17574_18026.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X24 VDPWR.t125 PFET_GATE.t11 a_11431_12690.t9 VDPWR.t124 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X25 a_10710_11860.t15 a_8454_18026.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X26 a_17290_7270.t2 a_16900_7270.t2 VDPWR.t187 VDPWR.t186 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X27 VDPWR.t363 VDPWR.t360 VDPWR.t362 VDPWR.t361 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X28 VDPWR.t105 a_16270_3380.t2 a_13650_3080.t2 VDPWR.t104 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X29 a_16510_7270.t1 a_13440_7240.t3 VDPWR.t203 VDPWR.t98 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X30 VDPWR.t97 a_10840_11590.t17 a_10710_11860.t2 VDPWR.t96 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X31 a_13750_11850.t12 a_17574_18026.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X32 a_14120_3110.t2 a_14280_3560.t2 VGND.t65 VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X33 V_CONT.t3 a_17580_6090.t3 VDPWR.t232 VDPWR.t231 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X34 VDPWR.t270 VGND.t327 a_23718_3560.t2 VDPWR.t269 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=1.2 ps=6.8 w=3 l=0.15
X35 VDPWR.t101 a_13650_3080.t3 a_14280_3560.t0 VDPWR.t100 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X36 a_13360_7270.t1 a_12360_3440.t2 VDPWR.t178 VDPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X37 a_11880_10030.t15 VDPWR.t377 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 VGND.t214 VGND.t266 a_11580_15080.t8 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X39 I_IN.t14 I_IN.t13 VGND.t109 VGND.t108 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X40 VDPWR.t370 a_20810_11490.t6 a_21100_10960.t4 VDPWR.t369 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X41 a_11880_10030.t16 VDPWR.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X42 VDPWR.t264 a_13750_11850.t13 a_11880_10030.t8 VDPWR.t263 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X43 VGND.t63 a_14860_6060.t2 a_14340_6060.t0 VGND.t62 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X44 a_21130_3020.t0 a_20510_3370.t3 a_20830_3320.t0 VGND.t140 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X45 VGND.t181 VDPWR.t428 a_23718_2840.t2 VGND.t180 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.6 ps=3.8 w=1.5 l=0.15
X46 a_19210_3370.t2 a_19910_3400.t2 VDPWR.t134 VDPWR.t133 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X47 VDPWR.t165 PFET_GATE.t12 I_IN.t9 VDPWR.t164 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X48 a_11880_10030.t17 VDPWR.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X49 VDPWR.t180 a_10840_11590.t15 a_10840_11590.t16 VDPWR.t179 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X50 a_10710_11860.t16 a_8454_18026.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X51 a_16960_3370.t0 a_17400_3080.t2 VDPWR.t207 VDPWR.t206 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X52 VGND.t93 a_19210_3370.t3 a_19120_3150.t2 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X53 a_16900_7270.t1 VDPWR.t429 a_16510_7270.t3 VGND.t278 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X54 a_10740_13170.t3 a_9573_16817.t8 a_10840_11590.t2 VGND.t142 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X55 VGND.t218 VGND.t259 a_11580_15080.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X56 VDPWR.t396 a_19210_3370.t4 a_18610_3400.t0 VDPWR.t395 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X57 VGND.t218 VGND.t258 a_11580_15080.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X58 VDPWR.t129 PFET_GATE.t13 a_11431_12690.t8 VDPWR.t128 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X59 a_10710_11860.t17 a_8454_18026.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X60 VDPWR.t268 VGND.t328 a_23198_3560.t1 VDPWR.t267 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=1.2 ps=6.8 w=3 l=0.15
X61 a_12490_3240.t2 a_12620_3080.t2 VGND.t315 VGND.t314 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X62 VGND.t265 VGND.t263 VGND.t265 VGND.t264 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0 ps=0 w=1.25 l=0.5
X63 VGND.t262 VGND.t260 VGND.t262 VGND.t261 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X64 a_17820_3240.t3 a_16740_3080.t4 VGND.t13 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X65 a_14340_7240.t1 a_13960_7240.t3 VGND.t9 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X66 a_13540_3080.t2 a_13650_3080.t4 VGND.t61 VGND.t60 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X67 VGND.t157 I_IN.t18 a_19930_11490.t5 VGND.t156 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X68 a_10710_11860.t18 a_8454_18026.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X69 VDPWR.t252 a_13880_11590.t12 a_13880_11590.t13 VDPWR.t251 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X70 VDPWR.t359 VDPWR.t356 VDPWR.t358 VDPWR.t357 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X71 VGND.t55 a_18610_3400.t2 a_19830_3020.t0 VGND.t54 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X72 VGND.t126 a_19690_10220.t7 a_19690_10220.t8 VGND.t125 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X73 a_12520_10060.t7 a_11880_10030.t18 VDPWR.t211 VDPWR.t210 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X74 a_19440_11540.t12 V_CONT.t8 a_19670_10930.t5 VDPWR.t394 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X75 a_21720_3150.t2 a_21810_3370.t3 VGND.t207 VGND.t206 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X76 VGND.t257 VGND.t254 VGND.t256 VGND.t255 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X77 a_19244_9974.t8 a_19244_9974.t7 VDPWR.t131 VDPWR.t130 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X78 a_11431_12690.t7 PFET_GATE.t14 VDPWR.t391 VDPWR.t390 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X79 a_11880_10030.t13 VDPWR.t353 VDPWR.t355 VDPWR.t354 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.45 ps=2.9 w=1 l=0.15
X80 VGND.t279 VDPWR.t430 a_23198_2840.t2 VGND.t47 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.6 ps=3.8 w=1.5 l=0.15
X81 a_15300_6090.t0 a_13440_7240.t4 VGND.t311 VGND.t310 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X82 VDPWR.t413 a_23280_5000.t3 a_24238_3560.t2 VDPWR.t412 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X83 a_14260_6510.t1 a_13360_6090.t3 VDPWR.t159 VDPWR.t158 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X84 a_13750_11850.t14 a_17574_18026.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X85 a_15920_7240.t1 a_15740_6090.t2 VDPWR.t109 VDPWR.t108 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X86 VDPWR.t70 a_13880_11590.t17 a_13750_11850.t1 VDPWR.t69 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X87 VDPWR.t352 VDPWR.t350 VDPWR.t352 VDPWR.t351 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X88 VGND.t273 a_20510_3370.t4 a_20420_3150.t2 VGND.t272 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X89 a_19790_10270.t6 a_19790_10270.t4 a_19790_10270.t5 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X90 a_17450_6090.t10 a_23224_12716.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X91 VDPWR.t183 a_10840_11590.t18 a_10710_11860.t4 VDPWR.t182 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X92 VDPWR.t284 a_20510_3370.t5 a_19910_3400.t1 VDPWR.t283 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X93 VDPWR.t163 PFET_GATE.t15 I_IN.t8 VDPWR.t162 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X94 VDPWR.t195 a_19530_3320.t2 a_19120_3150.t3 VDPWR.t194 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X95 a_16630_3080.t3 a_16960_3370.t3 VDPWR.t398 VDPWR.t397 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X96 a_21810_3370.t0 ua[1].t3 VGND.t271 VGND.t270 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X97 VGND.t11 V_CONT.t9 a_24238_2840.t0 VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X98 VGND.t174 a_19120_3150.t4 a_18610_3400.t1 VGND.t173 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X99 a_17450_6090.t2 a_19960_10960.t5 VGND.t129 VGND.t128 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X100 VGND.t313 a_19690_10220.t9 a_19790_10270.t12 VGND.t312 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X101 a_13880_6510.t1 a_13360_6090.t4 a_13440_6060.t1 VDPWR.t171 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X102 VDPWR.t375 PFET_GATE.t16 a_11431_12690.t6 VDPWR.t374 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X103 a_14860_3240.t3 a_13650_3080.t5 VGND.t21 VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X104 VGND.t40 a_19670_10930.t6 a_19960_10960.t4 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X105 a_14860_3240.t2 a_13650_3080.t6 VGND.t131 VGND.t130 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X106 a_10840_11590.t14 a_10840_11590.t13 VDPWR.t217 VDPWR.t216 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X107 a_12490_3240.t1 a_12620_3080.t3 VGND.t114 VGND.t113 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X108 a_10740_13170.t10 a_11431_12690.t13 a_10710_11860.t10 VGND.t324 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X109 a_14260_7270.t0 a_13360_7890.t3 VDPWR.t172 VDPWR.t158 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X110 I_IN.t4 PFET_GATE.t17 VDPWR.t78 VDPWR.t77 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X111 VDPWR.t213 a_11880_10030.t19 a_9573_16817.t4 VDPWR.t212 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X112 a_13540_3080.t1 a_13650_3080.t7 VGND.t304 VGND.t303 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X113 a_19930_11490.t4 I_IN.t19 VGND.t184 VGND.t183 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X114 VDPWR.t262 a_13750_11850.t15 a_11880_10030.t7 VDPWR.t261 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X115 a_14040_12560.t3 a_12520_10060.t8 a_13880_11590.t3 VGND.t124 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X116 a_17450_6090.t6 a_21100_10960.t6 VDPWR.t17 VDPWR.t16 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X117 a_15490_3110.t1 a_13650_3080.t8 a_15380_3110.t1 VGND.t95 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X118 VDPWR.t39 a_15260_7240.t2 a_14860_6060.t0 VDPWR.t38 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X119 a_22130_3320.t0 a_21210_3400.t3 VDPWR.t76 VDPWR.t75 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X120 VDPWR.t103 a_18610_3400.t3 a_16740_3080.t0 VDPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X121 a_11880_10030.t20 VDPWR.t422 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X122 PFET_GATE.t5 a_10710_11860.t19 VDPWR.t280 VDPWR.t279 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X123 a_13880_7270.t0 a_13360_7890.t4 a_13440_7240.t1 VDPWR.t171 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X124 VGND.t286 a_13440_7240.t5 a_13360_7890.t1 VGND.t285 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X125 VDPWR.t5 a_20830_3320.t2 a_20420_3150.t3 VDPWR.t4 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X126 a_14040_12560.t10 a_12520_10060.t9 a_13880_11590.t16 VGND.t293 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X127 VDPWR.t349 VDPWR.t347 VDPWR.t349 VDPWR.t348 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X128 VGND.t24 a_20420_3150.t4 a_19910_3400.t0 VGND.t23 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X129 VDPWR.t278 a_10710_11860.t20 PFET_GATE.t4 VDPWR.t277 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X130 a_11880_10030.t21 VDPWR.t423 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X131 a_10740_13170.t5 a_11431_12690.t14 a_10710_11860.t3 VGND.t74 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X132 a_22430_3020.t1 a_21810_3370.t4 a_22130_3320.t1 VGND.t141 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X133 a_17580_6090.t4 a_17290_6090.t2 sky130_fd_pr__cap_mim_m3_1 l=6.3 w=5.2
X134 a_20510_3370.t2 a_21210_3400.t4 VDPWR.t74 VDPWR.t73 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X135 a_10710_11860.t21 a_8454_18026.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X136 a_17290_6090.t0 a_16900_6090.t3 VGND.t297 VGND.t296 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X137 a_16510_6090.t0 a_13440_6060.t4 VGND.t26 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X138 a_11160_14080.t5 a_11880_10030.t22 VDPWR.t367 VDPWR.t366 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X139 VGND.t38 a_10354_16286.t0 VGND.t37 sky130_fd_pr__res_xhigh_po_0p35 l=17.96
X140 VDPWR.t8 a_21100_10960.t7 a_17450_6090.t5 VDPWR.t7 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X141 VDPWR.t292 a_13880_11590.t18 a_13750_11850.t9 VDPWR.t291 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X142 a_10740_13170.t8 a_11431_12690.t15 a_10710_11860.t8 VGND.t269 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X143 a_13360_6090.t0 ua[0].t1 VGND.t149 VGND.t148 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X144 a_10710_11860.t22 a_8454_18026.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X145 a_16960_3370.t2 a_16740_3080.t5 a_17430_3110.t1 VGND.t118 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X146 VGND.t281 VDPWR.t431 a_10740_13170.t9 VGND.t280 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X147 a_13750_11850.t16 a_17574_18026.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X148 a_13240_14080.t0 a_11160_14080.t0 a_11160_14080.t1 VGND.t190 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X149 VGND.t301 a_12620_3080.t4 a_15570_3080.t0 VGND.t300 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X150 VGND.t253 VGND.t250 VGND.t252 VGND.t251 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X151 VGND.t34 a_19690_10220.t10 a_19790_10270.t11 VGND.t33 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X152 a_20810_11490.t3 a_20810_11490.t2 VDPWR.t243 VDPWR.t242 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X153 VGND.t214 VGND.t242 a_11580_15080.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X154 VDPWR.t346 VDPWR.t344 VDPWR.t346 VDPWR.t345 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0 ps=0 w=2.5 l=0.5
X155 VDPWR.t33 a_14280_3560.t3 a_14230_3430.t1 VDPWR.t32 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X156 a_13750_11850.t17 a_17574_18026.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X157 a_11880_10030.t6 a_13750_11850.t18 VDPWR.t260 VDPWR.t259 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X158 a_16900_6090.t1 a_16510_6090.t2 VDPWR.t230 VDPWR.t229 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X159 VGND.t116 a_15590_7240.t2 a_15260_7240.t0 VGND.t115 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X160 a_19690_10220.t6 a_19690_10220.t5 VGND.t167 VGND.t166 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X161 a_19960_10960.t2 a_19930_11490.t6 a_19440_11540.t0 VDPWR.t60 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X162 VDPWR.t177 a_13440_6060.t5 a_15300_6510.t2 VDPWR.t176 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X163 VDPWR.t89 a_19244_9974.t5 a_19244_9974.t6 VDPWR.t88 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X164 a_11880_10030.t23 VDPWR.t368 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X165 a_14992_19436.t0 V_CONT.t4 VGND.t46 sky130_fd_pr__res_xhigh_po_0p35 l=7.52
X166 a_17580_7270.t0 a_17290_7270.t3 I_IN.t7 VGND.t110 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X167 VDPWR.t387 a_11880_10030.t24 a_9573_16817.t3 VDPWR.t386 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X168 VDPWR.t121 a_23280_5000.t1 a_23280_5000.t2 VDPWR.t120 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X169 a_14780_6510.t0 a_13960_6060.t3 a_14340_6060.t2 VDPWR.t132 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X170 VGND.t73 a_21810_3370.t5 a_21720_3150.t1 VGND.t72 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X171 a_11880_10030.t25 VDPWR.t388 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X172 a_17580_7270.t3 a_17290_7270.t0 sky130_fd_pr__cap_mim_m3_1 l=3.8 w=2.7
X173 VDPWR.t62 a_21810_3370.t6 a_21210_3400.t0 VDPWR.t61 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X174 a_13880_11590.t11 a_13880_11590.t10 VDPWR.t127 VDPWR.t126 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X175 VGND.t218 VGND.t246 a_12520_10060.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X176 PFET_GATE.t3 a_10710_11860.t23 VDPWR.t276 VDPWR.t275 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X177 VDPWR.t343 VDPWR.t341 VDPWR.t343 VDPWR.t342 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X178 a_8454_18026.t0 PFET_GATE.t0 VGND.t155 sky130_fd_pr__res_high_po_0p35 l=2.05
X179 VGND.t159 a_19960_10960.t6 a_17450_6090.t3 VGND.t158 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X180 a_10710_11860.t24 a_8454_18026.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X181 a_19790_10270.t10 a_19690_10220.t11 VGND.t299 VGND.t298 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X182 a_14040_12560.t7 a_10354_16286.t7 a_13750_11850.t6 VGND.t211 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X183 a_16900_7270.t0 VGND.t329 a_16510_7270.t2 VDPWR.t229 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X184 a_17820_3240.t2 a_16740_3080.t6 VGND.t163 VGND.t162 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X185 a_9573_16817.t6 VDPWR.t338 VDPWR.t340 VDPWR.t339 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X186 VGND.t249 VGND.t247 VGND.t249 VGND.t248 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X187 VGND.t330 a_14992_19436.t1 sky130_fd_pr__cap_mim_m3_1 l=60 w=69.8
X188 a_10710_11860.t25 a_8454_18026.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X189 VGND.t245 VGND.t243 VGND.t245 VGND.t244 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X190 a_10710_11860.t9 a_10840_11590.t19 VDPWR.t286 VDPWR.t285 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X191 a_13750_11850.t19 a_17574_18026.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X192 a_14780_7270.t1 a_13960_7240.t4 a_14340_7240.t2 VDPWR.t132 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X193 VGND.t5 a_14340_7240.t3 a_13960_7240.t0 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X194 a_13540_3080.t3 a_13870_3370.t3 VDPWR.t405 VDPWR.t404 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X195 a_11431_12690.t5 PFET_GATE.t18 VDPWR.t223 VDPWR.t222 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X196 a_14040_12560.t5 a_10354_16286.t8 a_13750_11850.t5 VGND.t210 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X197 VDPWR.t119 a_19910_3400.t3 a_19210_3370.t1 VDPWR.t118 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X198 a_10710_11860.t0 a_10840_11590.t20 VDPWR.t1 VDPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X199 a_10354_16286.t5 a_11880_10030.t26 VDPWR.t417 VDPWR.t416 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X200 a_13750_11850.t20 a_17574_18026.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X201 a_16740_3080.t2 a_18610_3400.t4 VGND.t172 VGND.t171 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X202 VGND.t241 VGND.t238 VGND.t240 VGND.t239 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X203 VGND.t317 a_13960_7240.t5 a_13440_7240.t2 VGND.t316 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X204 VGND.t201 a_21720_3150.t4 a_21210_3400.t1 VGND.t200 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X205 a_13750_11850.t21 a_17574_18026.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X206 a_10840_11590.t12 a_10840_11590.t11 VDPWR.t95 VDPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X207 a_13960_6060.t2 a_13360_6090.t5 VGND.t292 VGND.t291 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X208 a_19440_11540.t6 a_19440_11540.t4 a_19440_11540.t5 VDPWR.t389 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X209 a_10710_11860.t6 a_11431_12690.t16 a_10740_13170.t7 VGND.t196 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X210 VGND.t89 a_15920_7240.t2 a_15590_7240.t0 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X211 VDPWR.t419 a_11880_10030.t27 a_12520_10060.t6 VDPWR.t418 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X212 a_11880_10030.t28 VDPWR.t196 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X213 a_15920_7240.t0 a_15740_6090.t3 VGND.t36 VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X214 a_21810_3370.t1 ua[1].t4 VDPWR.t381 VDPWR.t380 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X215 VDPWR.t19 a_17450_6090.t11 a_19930_11490.t3 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X216 a_15740_6090.t1 a_15300_6510.t3 VDPWR.t415 VDPWR.t414 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X217 a_19790_10270.t1 a_19930_11490.t7 a_21100_10960.t1 VGND.t53 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X218 VGND.t3 a_16740_3080.t7 a_16630_3080.t1 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X219 a_18230_3320.t1 a_13650_3080.t9 VDPWR.t168 VDPWR.t167 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X220 I_IN.t11 PFET_GATE.t19 VDPWR.t205 VDPWR.t204 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X221 a_13360_6090.t1 a_13440_6060.t6 a_13360_6510.t1 VDPWR.t11 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X222 a_17450_6090.t12 a_23224_9624.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X223 a_23310_2840.t1 ua[1].t5 a_23198_2840.t0 VGND.t94 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.16
X224 a_13120_3110.t1 a_12620_3080.t5 a_13010_3110.t1 VGND.t307 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X225 a_13440_6060.t0 a_13360_6090.t6 VGND.t15 VGND.t14 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X226 VDPWR.t198 a_11880_10030.t29 a_10354_16286.t4 VDPWR.t197 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X227 VGND.t331 V_CONT.t7 sky130_fd_pr__cap_mim_m3_1 l=60 w=13.8
X228 V_CONT.t6 a_17580_7270.t4 VGND.t194 VGND.t193 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X229 a_10710_11860.t26 a_8454_18026.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X230 a_11431_12690.t4 PFET_GATE.t20 VDPWR.t25 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X231 a_11431_12690.t11 VDPWR.t335 VDPWR.t337 VDPWR.t336 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X232 a_11880_10030.t2 a_11160_14080.t6 a_12520_10060.t2 VDPWR.t219 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X233 VDPWR.t193 a_20810_11490.t0 a_20810_11490.t1 VDPWR.t192 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X234 VDPWR.t45 a_15380_3110.t2 a_14860_3240.t0 VDPWR.t44 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X235 VDPWR.t334 VDPWR.t332 a_11880_10030.t12 VDPWR.t333 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X236 VDPWR.t136 a_19244_9974.t9 a_19440_11540.t3 VDPWR.t135 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X237 a_18530_3110.t0 a_16740_3080.t8 a_18230_3320.t0 VGND.t119 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X238 a_13750_11850.t2 a_13880_11590.t19 VDPWR.t185 VDPWR.t184 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X239 a_13750_11850.t22 a_17574_18026.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X240 a_14450_3110.t1 a_12620_3080.t6 a_14120_3110.t1 VGND.t127 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X241 a_10354_16286.t3 a_11880_10030.t30 VDPWR.t146 VDPWR.t145 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X242 a_19244_9974.t4 a_19244_9974.t3 VDPWR.t68 VDPWR.t67 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X243 a_13360_7890.t0 a_13440_7240.t6 a_13360_7270.t0 VDPWR.t11 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X244 VGND.t103 a_19670_10930.t1 a_19670_10930.t2 VGND.t102 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X245 a_14040_12560.t0 a_12520_10060.t10 a_13880_11590.t0 VGND.t44 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X246 a_13750_11850.t23 a_17574_18026.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X247 a_11160_14080.t4 a_11880_10030.t31 VDPWR.t148 VDPWR.t147 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X248 a_11880_10030.t5 a_13750_11850.t24 VDPWR.t258 VDPWR.t257 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X249 VGND.t105 a_16630_3080.t4 a_16270_3380.t1 VGND.t104 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X250 VGND.t80 a_19910_3400.t4 a_21130_3020.t1 VGND.t79 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X251 I_IN.t1 VDPWR.t329 VDPWR.t331 VDPWR.t330 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X252 I_IN.t3 PFET_GATE.t21 VDPWR.t64 VDPWR.t63 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X253 VGND.t237 VGND.t235 VGND.t237 VGND.t236 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X254 a_9573_16817.t2 a_11880_10030.t32 VDPWR.t91 VDPWR.t90 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X255 a_21100_10960.t0 a_20810_11490.t7 VDPWR.t29 VDPWR.t28 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X256 VGND.t234 VGND.t231 VGND.t233 VGND.t232 sky130_fd_pr__nfet_01v8 ad=0.625 pd=3.5 as=0 ps=0 w=1.25 l=0.5
X257 a_23310_2840.t0 ua[1].t6 a_23198_3560.t0 VDPWR.t166 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.16
X258 a_11880_10030.t4 a_13750_11850.t25 VDPWR.t256 VDPWR.t255 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X259 a_19120_3150.t1 a_19210_3370.t5 VGND.t99 VGND.t98 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X260 a_13750_11850.t4 a_10354_16286.t9 a_14040_12560.t4 VGND.t209 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X261 a_17580_6090.t2 a_17290_6090.t3 a_17450_6090.t0 VDPWR.t6 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X262 a_19440_11540.t10 a_19244_9974.t10 VDPWR.t170 VDPWR.t169 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X263 a_15570_3080.t2 a_12620_3080.t7 VDPWR.t59 VDPWR.t58 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X264 VGND.t288 a_11431_12690.t12 VGND.t287 sky130_fd_pr__res_xhigh_po_0p35 l=1
X265 a_13750_11850.t26 a_17574_18026.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X266 a_11431_12690.t3 PFET_GATE.t22 VDPWR.t156 VDPWR.t155 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X267 VGND.t218 VGND.t230 a_11580_15080.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X268 VDPWR.t266 VGND.t332 a_24238_3560.t1 VDPWR.t265 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=1.2 ps=6.8 w=3 l=0.15
X269 a_13650_3080.t1 a_16270_3380.t3 VDPWR.t49 VDPWR.t48 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X270 VGND.t86 a_14860_6060.t3 a_14340_7240.t0 VGND.t85 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X271 VDPWR.t93 a_11880_10030.t33 a_11160_14080.t3 VDPWR.t92 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X272 VDPWR.t189 a_16740_3080.t9 a_17400_3080.t1 VDPWR.t188 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X273 a_13880_11590.t9 a_13880_11590.t8 VDPWR.t141 VDPWR.t140 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X274 VGND.t84 a_12360_3440.t3 a_14120_3110.t0 VGND.t83 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X275 VDPWR.t161 a_15590_7240.t3 a_15260_7240.t1 VDPWR.t160 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X276 PFET_GATE.t2 a_10710_11860.t27 VDPWR.t274 VDPWR.t273 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X277 a_19790_10270.t9 a_19690_10220.t12 VGND.t306 VGND.t305 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X278 a_10840_11590.t0 a_9573_16817.t9 a_10740_13170.t2 VGND.t195 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X279 a_17450_6090.t8 a_19960_10960.t7 VGND.t277 VGND.t276 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X280 a_11880_10030.t34 VDPWR.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X281 a_16900_6090.t0 a_16510_6090.t3 VGND.t76 VGND.t75 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X282 VDPWR.t328 VDPWR.t326 a_11431_12690.t10 VDPWR.t327 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X283 a_17580_7270.t2 a_16900_7270.t3 I_IN.t10 VDPWR.t6 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X284 a_15300_6510.t1 a_13440_6060.t7 a_15300_6090.t1 VGND.t143 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X285 VGND.t282 VDPWR.t432 a_24238_2840.t2 VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.6 ps=3.8 w=1.5 l=0.15
X286 VGND.t32 a_9573_16817.t0 VGND.t31 sky130_fd_pr__res_xhigh_po_0p35 l=10.04
X287 a_13960_6060.t0 a_14340_6060.t3 a_14260_6510.t0 VDPWR.t117 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X288 a_11880_10030.t35 VDPWR.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X289 a_19670_10930.t0 V_CONT.t10 a_19440_11540.t9 VDPWR.t157 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X290 a_10710_11860.t1 a_10840_11590.t21 VDPWR.t53 VDPWR.t52 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X291 a_20420_3150.t1 a_20510_3370.t6 VGND.t203 VGND.t202 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X292 a_17320_3110.t1 a_16270_3380.t4 VGND.t187 VGND.t186 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X293 a_14340_6060.t1 a_13960_6060.t4 VGND.t71 VGND.t70 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X294 a_10840_11590.t4 a_9573_16817.t10 a_10740_13170.t1 VGND.t182 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X295 V_CONT.t2 a_17580_6090.t5 VDPWR.t239 VDPWR.t238 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X296 I_IN.t0 PFET_GATE.t23 VDPWR.t10 VDPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X297 VDPWR.t55 a_23280_5000.t4 a_23718_3560.t0 VDPWR.t54 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X298 a_19790_10270.t3 a_19790_10270.t2 a_19790_10270.t3 VGND.t170 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X299 a_19530_3320.t0 a_18610_3400.t5 VDPWR.t247 VDPWR.t246 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X300 a_13750_11850.t0 a_13880_11590.t20 VDPWR.t21 VDPWR.t20 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X301 a_10710_11860.t28 a_8454_18026.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X302 a_19120_3150.t0 a_19210_3370.t6 VGND.t123 VGND.t122 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X303 a_13750_11850.t27 a_17574_18026.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X304 VGND.t17 a_13240_14080.t1 a_13240_14080.t0 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X305 VGND.t229 VGND.t227 VGND.t229 VGND.t228 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X306 VDPWR.t43 a_13960_6060.t5 a_13880_6510.t0 VDPWR.t42 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X307 a_11580_15080.t0 a_10354_16286.t1 VGND.t45 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X308 a_10710_11860.t29 a_8454_18026.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X309 a_11431_12690.t2 PFET_GATE.t24 VDPWR.t27 VDPWR.t26 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X310 VGND.t197 V_CONT.t11 a_23718_2840.t1 VGND.t180 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X311 VDPWR.t325 VDPWR.t323 PFET_GATE.t9 VDPWR.t324 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X312 a_23830_2840.t0 a_23310_2840.t2 a_23718_2840.t0 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.16
X313 VGND.t30 a_12620_3080.t8 a_12490_3240.t0 VGND.t29 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X314 a_13750_11850.t28 a_17574_18026.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X315 VGND.t59 a_17820_3240.t4 a_17400_3080.t0 VGND.t58 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X316 a_17580_7270.t1 a_16900_7270.t4 VGND.t91 VGND.t90 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X317 a_13960_7240.t1 a_14340_7240.t4 a_14260_7270.t1 VDPWR.t117 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X318 VDPWR.t322 VDPWR.t320 I_IN.t2 VDPWR.t321 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X319 VGND.t67 a_19960_10960.t8 a_17450_6090.t1 VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X320 a_19440_11540.t11 a_19244_9974.t11 VDPWR.t379 VDPWR.t378 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X321 VGND.t152 a_13650_3080.t10 a_13540_3080.t0 VGND.t151 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X322 a_10840_11590.t10 a_10840_11590.t9 VDPWR.t150 VDPWR.t149 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X323 a_11880_10030.t36 VDPWR.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X324 VGND.t69 a_15570_3080.t3 a_15490_3110.t0 VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X325 a_10840_11590.t3 a_9573_16817.t11 a_10740_13170.t0 VGND.t274 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X326 a_19830_3020.t1 a_19210_3370.t7 a_19530_3320.t1 VGND.t43 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X327 a_13750_11850.t29 a_17574_18026.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 a_16740_3080.t1 a_18610_3400.t6 VDPWR.t209 VDPWR.t208 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X329 a_13750_11850.t30 a_17574_18026.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X330 VGND.t147 a_12360_3440.t4 a_13120_3110.t0 VGND.t146 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X331 a_20810_11490.t5 V_CONT.t12 a_19790_10270.t8 VGND.t7 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X332 a_19244_9974.t0 a_19690_10220.t0 sky130_fd_pr__res_generic_po w=0.33 l=2.4
X333 VDPWR.t407 PFET_GATE.t25 a_11431_12690.t1 VDPWR.t406 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X334 VDPWR.t87 a_19244_9974.t12 a_19440_11540.t2 VDPWR.t86 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X335 VDPWR.t383 a_23280_5000.t5 a_23198_3560.t2 VDPWR.t382 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X336 VDPWR.t199 a_13960_7240.t6 a_13880_7270.t1 VDPWR.t42 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X337 a_19960_10960.t3 a_19670_10930.t7 VGND.t268 VGND.t267 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X338 a_20830_3320.t1 a_19910_3400.t5 VDPWR.t411 VDPWR.t410 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X339 a_19960_10960.t0 a_23224_9624.t1 VGND.t19 sky130_fd_pr__res_xhigh_po_0p35 l=0.86
X340 a_20420_3150.t0 a_20510_3370.t7 VGND.t290 VGND.t289 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X341 a_13880_11590.t7 a_13880_11590.t6 VDPWR.t288 VDPWR.t287 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X342 a_10710_11860.t30 a_8454_18026.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X343 I_IN.t17 PFET_GATE.t26 VDPWR.t393 VDPWR.t392 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X344 VDPWR.t139 a_11880_10030.t37 a_10354_16286.t2 VDPWR.t138 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X345 VDPWR.t421 a_15920_7240.t3 a_15590_7240.t1 VDPWR.t420 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X346 a_11880_10030.t38 VDPWR.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X347 VGND.t48 V_CONT.t13 a_23198_2840.t1 VGND.t47 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X348 VDPWR.t228 a_16740_3080.t10 a_16270_3380.t0 VDPWR.t227 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X349 VGND.t1 a_21210_3400.t5 a_22430_3020.t0 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X350 a_23280_5000.t0 V_CONT.t14 VGND.t326 VGND.t325 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X351 a_19930_11490.t2 a_17450_6090.t13 VDPWR.t154 VDPWR.t153 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X352 a_11880_10030.t39 VDPWR.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X353 a_15740_6090.t0 a_15300_6510.t4 VGND.t135 VGND.t134 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X354 VGND.t161 a_17580_7270.t5 V_CONT.t5 VGND.t160 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X355 VGND.t319 a_14860_3240.t4 a_14280_3560.t1 VGND.t318 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X356 a_13750_11850.t10 a_13880_11590.t21 VDPWR.t365 VDPWR.t364 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X357 a_23830_2840.t1 a_23310_2840.t3 a_23718_3560.t1 VDPWR.t224 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.16
X358 VGND.t121 a_13650_3080.t11 a_14860_3240.t1 VGND.t120 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X359 VDPWR.t403 a_13010_3110.t2 a_12490_3240.t3 VDPWR.t402 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X360 VDPWR.t319 VDPWR.t316 VDPWR.t318 VDPWR.t317 sky130_fd_pr__pfet_01v8 ad=1.25 pd=6 as=0 ps=0 w=2.5 l=0.5
X361 VGND.t169 a_12490_3240.t4 a_12360_3440.t1 VGND.t168 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X362 VGND.t139 a_13440_6060.t8 a_13360_6090.t2 VGND.t138 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X363 a_10710_11860.t31 a_8454_18026.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X364 VDPWR.t215 PFET_GATE.t27 I_IN.t12 VDPWR.t214 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X365 a_13750_11850.t31 a_17574_18026.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X366 VGND.t295 a_13540_3080.t4 a_12620_3080.t1 VGND.t294 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X367 VGND.t101 a_12520_10060.t0 VGND.t100 sky130_fd_pr__res_xhigh_po_0p35 l=17.96
X368 VDPWR.t372 a_22130_3320.t2 a_21720_3150.t3 VDPWR.t371 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X369 VDPWR.t15 a_12620_3080.t9 a_15570_3080.t1 VDPWR.t14 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X370 a_17290_7270.t1 a_16900_7270.t5 VGND.t97 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X371 a_10710_11860.t32 a_8454_18026.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X372 VGND.t199 a_16270_3380.t5 a_13650_3080.t0 VGND.t198 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X373 a_16510_7270.t0 a_13440_7240.t7 VGND.t205 VGND.t204 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X374 a_13750_11850.t32 a_17574_18026.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X375 a_13870_3370.t2 a_12620_3080.t10 VDPWR.t35 VDPWR.t34 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X376 VDPWR.t51 a_13880_11590.t4 a_13880_11590.t5 VDPWR.t50 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X377 a_13750_11850.t33 a_17574_18026.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X378 VGND.t154 a_19690_10220.t3 a_19690_10220.t4 VGND.t153 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X379 VGND.t214 VGND.t213 a_11580_15080.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X380 VDPWR.t272 a_10710_11860.t33 PFET_GATE.t1 VDPWR.t271 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X381 a_12520_10060.t5 a_11880_10030.t40 VDPWR.t111 VDPWR.t110 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X382 a_17574_18026.t0 a_11880_10030.t0 VGND.t18 sky130_fd_pr__res_high_po_0p35 l=2.05
X383 a_19930_11490.t1 a_17450_6090.t14 VDPWR.t235 VDPWR.t234 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X384 a_13360_7890.t2 a_12360_3440.t5 VGND.t145 VGND.t144 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X385 VDPWR.t315 VDPWR.t312 VDPWR.t314 VDPWR.t313 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X386 a_11880_10030.t11 VDPWR.t309 VDPWR.t311 VDPWR.t310 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X387 a_11880_10030.t41 VDPWR.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X388 a_13880_11590.t2 a_12520_10060.t11 a_14040_12560.t2 VGND.t87 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X389 VDPWR.t308 VDPWR.t306 VDPWR.t308 VDPWR.t307 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X390 VDPWR.t107 a_14860_6060.t4 a_14780_6510.t1 VDPWR.t106 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X391 a_17450_6090.t4 a_21100_10960.t8 VDPWR.t13 VDPWR.t12 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X392 a_14040_12560.t9 VDPWR.t433 VGND.t284 VGND.t283 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1.01 ps=6.15 w=2.5 l=5
X393 VDPWR.t221 a_21210_3400.t6 a_20510_3370.t1 VDPWR.t220 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X394 a_11880_10030.t42 VDPWR.t173 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X395 VDPWR.t305 VDPWR.t302 VDPWR.t304 VDPWR.t303 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X396 VDPWR.t249 a_10840_11590.t22 a_10710_11860.t7 VDPWR.t248 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X397 VGND.t226 VGND.t223 VGND.t225 VGND.t224 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X398 a_19440_11540.t1 a_19930_11490.t8 a_19960_10960.t1 VDPWR.t85 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X399 a_12520_10060.t1 a_11160_14080.t7 a_11880_10030.t1 VDPWR.t218 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X400 a_19210_3370.t0 a_19910_3400.t6 VGND.t112 VGND.t111 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X401 VGND.t222 VGND.t219 VGND.t221 VGND.t220 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X402 VGND.t218 VGND.t217 a_11580_15080.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X403 a_13880_11590.t1 a_12520_10060.t12 a_14040_12560.t1 VGND.t81 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X404 a_10710_11860.t34 a_8454_18026.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X405 PFET_GATE.t8 VDPWR.t299 VDPWR.t301 VDPWR.t300 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X406 a_17430_3110.t0 a_17400_3080.t3 a_17320_3110.t0 VGND.t322 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X407 VDPWR.t175 a_11880_10030.t43 a_11160_14080.t2 VDPWR.t174 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X408 a_17580_6090.t0 a_16900_6090.t4 a_17450_6090.t9 VGND.t302 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X409 a_10710_11860.t35 a_8454_18026.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X410 VDPWR.t298 VDPWR.t296 a_9573_16817.t5 VDPWR.t297 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X411 VDPWR.t233 a_14860_6060.t5 a_14780_7270.t0 VDPWR.t106 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X412 VGND.t216 VGND.t215 a_11580_15080.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X413 a_14230_3430.t0 a_12360_3440.t6 a_13870_3370.t1 VDPWR.t250 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X414 VDPWR.t241 a_10840_11590.t7 a_10840_11590.t8 VDPWR.t240 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X415 a_10710_11860.t5 a_11431_12690.t17 a_10740_13170.t6 VGND.t177 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X416 a_19790_10270.t7 V_CONT.t15 a_20810_11490.t4 VGND.t275 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X417 VDPWR.t237 a_17450_6090.t15 a_19930_11490.t0 VDPWR.t236 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X418 a_15300_6510.t0 a_13440_7240.t8 VDPWR.t3 VDPWR.t2 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.805 ps=5 w=2 l=0.15
X419 VDPWR.t226 a_17580_6090.t6 V_CONT.t1 VDPWR.t225 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X420 a_17580_6090.t1 a_16900_6090.t5 VDPWR.t409 VDPWR.t408 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X421 a_11880_10030.t44 VDPWR.t142 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X422 a_21720_3150.t0 a_21810_3370.t7 VGND.t57 VGND.t56 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X423 VDPWR.t425 a_16270_3380.t6 a_16960_3370.t1 VDPWR.t424 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X424 VGND.t78 a_14340_6060.t4 a_13960_6060.t1 VGND.t77 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X425 a_9573_16817.t1 a_11880_10030.t45 VDPWR.t144 VDPWR.t143 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X426 a_13750_11850.t34 a_17574_18026.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X427 a_16630_3080.t0 a_16740_3080.t11 VGND.t165 VGND.t164 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X428 VDPWR.t116 PFET_GATE.t28 I_IN.t6 VDPWR.t115 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X429 VGND.t50 a_16740_3080.t12 a_17820_3240.t1 VGND.t49 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X430 a_10710_11860.t36 a_8454_18026.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X431 VDPWR.t290 a_13880_11590.t22 a_13750_11850.t8 VDPWR.t289 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X432 a_13750_11850.t35 a_17574_18026.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X433 VGND.t137 a_13960_6060.t6 a_13440_6060.t2 VGND.t136 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X434 a_21100_10960.t2 a_19930_11490.t9 a_19790_10270.t0 VGND.t82 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X435 ua[1].t1 a_23830_2840.t3 a_24238_2840.t1 VGND.t323 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.16
X436 a_13960_7240.t2 a_13360_7890.t5 VGND.t321 VGND.t320 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X437 VDPWR.t82 a_13650_3080.t12 a_12620_3080.t0 VDPWR.t81 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X438 VDPWR.t201 PFET_GATE.t29 a_11431_12690.t0 VDPWR.t200 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X439 a_15380_3110.t0 a_15570_3080.t4 VDPWR.t41 VDPWR.t40 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X440 a_13750_11850.t3 a_10354_16286.t10 a_14040_12560.t6 VGND.t208 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X441 a_11880_10030.t46 VDPWR.t384 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X442 a_13010_3110.t0 a_12360_3440.t7 VDPWR.t245 VDPWR.t244 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X443 VGND.t133 a_15260_7240.t3 a_14860_6060.t1 VGND.t132 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X444 VGND.t189 a_13650_3080.t13 a_18530_3110.t1 VGND.t188 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X445 a_19690_10220.t2 a_19690_10220.t1 VGND.t28 VGND.t27 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X446 VDPWR.t295 VDPWR.t293 a_11880_10030.t10 VDPWR.t294 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X447 a_11880_10030.t47 VDPWR.t385 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X448 VDPWR.t191 a_17580_6090.t7 V_CONT.t0 VDPWR.t190 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X449 a_13870_3370.t0 a_13650_3080.t14 a_14450_3110.t0 VGND.t150 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X450 VDPWR.t37 a_19244_9974.t1 a_19244_9974.t2 VDPWR.t36 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X451 VDPWR.t152 a_10840_11590.t5 a_10840_11590.t6 VDPWR.t151 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X452 a_11880_10030.t48 VDPWR.t399 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X453 a_13440_7240.t0 a_13360_7890.t6 VGND.t192 VGND.t191 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X454 VDPWR.t84 a_12620_3080.t11 a_12360_3440.t0 VDPWR.t83 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X455 VDPWR.t401 a_11880_10030.t49 a_12520_10060.t4 VDPWR.t400 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X456 a_23224_12716.t1 a_21100_10960.t3 VGND.t185 sky130_fd_pr__res_xhigh_po_0p35 l=1.14
X457 VDPWR.t254 a_13750_11850.t36 a_11880_10030.t3 VDPWR.t253 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
R0 a_10354_16286.n3 a_10354_16286.t10 291.502
R1 a_10354_16286.n3 a_10354_16286.t7 291.288
R2 a_10354_16286.n4 a_10354_16286.t6 291.288
R3 a_10354_16286.n5 a_10354_16286.t8 291.288
R4 a_10354_16286.n6 a_10354_16286.t9 291.288
R5 a_10354_16286.n8 a_10354_16286.t1 148.653
R6 a_10354_16286.n2 a_10354_16286.n0 105.609
R7 a_10354_16286.n2 a_10354_16286.n1 104.484
R8 a_10354_16286.t0 a_10354_16286.n8 60.2462
R9 a_10354_16286.n8 a_10354_16286.n7 21.4246
R10 a_10354_16286.n7 a_10354_16286.n2 14.2349
R11 a_10354_16286.n0 a_10354_16286.t2 13.1338
R12 a_10354_16286.n0 a_10354_16286.t5 13.1338
R13 a_10354_16286.n1 a_10354_16286.t4 13.1338
R14 a_10354_16286.n1 a_10354_16286.t3 13.1338
R15 a_10354_16286.n7 a_10354_16286.n6 6.43621
R16 a_10354_16286.n6 a_10354_16286.n5 0.643357
R17 a_10354_16286.n4 a_10354_16286.n3 0.643357
R18 a_10354_16286.n5 a_10354_16286.n4 0.214786
R19 a_14040_12560.n5 a_14040_12560.n0 199.935
R20 a_14040_12560.n0 a_14040_12560.n4 199.53
R21 a_14040_12560.n0 a_14040_12560.n3 199.53
R22 a_14040_12560.n0 a_14040_12560.n2 199.53
R23 a_14040_12560.n0 a_14040_12560.n1 199.53
R24 a_14040_12560.n0 a_14040_12560.t9 56.2681
R25 a_14040_12560.n4 a_14040_12560.t2 48.0005
R26 a_14040_12560.n4 a_14040_12560.t7 48.0005
R27 a_14040_12560.n3 a_14040_12560.t8 48.0005
R28 a_14040_12560.n3 a_14040_12560.t3 48.0005
R29 a_14040_12560.n2 a_14040_12560.t1 48.0005
R30 a_14040_12560.n2 a_14040_12560.t5 48.0005
R31 a_14040_12560.n1 a_14040_12560.t4 48.0005
R32 a_14040_12560.n1 a_14040_12560.t10 48.0005
R33 a_14040_12560.n5 a_14040_12560.t6 48.0005
R34 a_14040_12560.t0 a_14040_12560.n5 48.0005
R35 a_13750_11850.n6 a_13750_11850.t24 363.909
R36 a_13750_11850.n5 a_13750_11850.t15 351.974
R37 a_13750_11850.n5 a_13750_11850.n10 299.25
R38 a_13750_11850.n5 a_13750_11850.n12 299.25
R39 a_13750_11850.n6 a_13750_11850.n9 299.25
R40 a_13750_11850.n7 a_13750_11850.t4 242.968
R41 a_13750_11850.n14 a_13750_11850.n13 200.477
R42 a_13750_11850.n15 a_13750_11850.n14 199.727
R43 a_13750_11850.n11 a_13750_11850.t25 194.809
R44 a_13750_11850.n11 a_13750_11850.t36 194.809
R45 a_13750_11850.n8 a_13750_11850.t18 194.809
R46 a_13750_11850.n8 a_13750_11850.t13 194.809
R47 a_13750_11850.n5 a_13750_11850.n11 163.097
R48 a_13750_11850.n7 a_13750_11850.n8 161.653
R49 a_13750_11850.n13 a_13750_11850.t6 48.0005
R50 a_13750_11850.n13 a_13750_11850.t3 48.0005
R51 a_13750_11850.n15 a_13750_11850.t5 48.0005
R52 a_13750_11850.t7 a_13750_11850.n15 48.0005
R53 a_13750_11850.n10 a_13750_11850.t9 39.4005
R54 a_13750_11850.n10 a_13750_11850.t0 39.4005
R55 a_13750_11850.n12 a_13750_11850.t1 39.4005
R56 a_13750_11850.n12 a_13750_11850.t10 39.4005
R57 a_13750_11850.n9 a_13750_11850.t8 39.4005
R58 a_13750_11850.n9 a_13750_11850.t2 39.4005
R59 a_13750_11850.n6 a_13750_11850.n4 13.9592
R60 a_13750_11850.n14 a_13750_11850.n7 5.2505
R61 a_13750_11850.n2 a_13750_11850.t30 4.8248
R62 a_13750_11850.n0 a_13750_11850.t21 4.5005
R63 a_13750_11850.n0 a_13750_11850.t14 4.5005
R64 a_13750_11850.n0 a_13750_11850.t17 4.5005
R65 a_13750_11850.n3 a_13750_11850.t12 4.5005
R66 a_13750_11850.n3 a_13750_11850.t33 4.5005
R67 a_13750_11850.n3 a_13750_11850.t22 4.5005
R68 a_13750_11850.n3 a_13750_11850.t28 4.5005
R69 a_13750_11850.n2 a_13750_11850.t19 4.5005
R70 a_13750_11850.n2 a_13750_11850.t23 4.5005
R71 a_13750_11850.n0 a_13750_11850.t29 4.5005
R72 a_13750_11850.n0 a_13750_11850.t20 4.5005
R73 a_13750_11850.n1 a_13750_11850.t26 4.5005
R74 a_13750_11850.n1 a_13750_11850.t16 4.5005
R75 a_13750_11850.n1 a_13750_11850.t11 4.5005
R76 a_13750_11850.n1 a_13750_11850.t31 4.5005
R77 a_13750_11850.n4 a_13750_11850.t34 4.5005
R78 a_13750_11850.n4 a_13750_11850.t27 4.5005
R79 a_13750_11850.n4 a_13750_11850.t32 4.5005
R80 a_13750_11850.n4 a_13750_11850.t35 4.5005
R81 a_13750_11850.n1 a_13750_11850.n0 1.9275
R82 a_13750_11850.n7 a_13750_11850.n6 1.74149
R83 a_13750_11850.n0 a_13750_11850.n3 1.3165
R84 a_13750_11850.n3 a_13750_11850.n2 1.3165
R85 a_13750_11850.n4 a_13750_11850.n1 1.3118
R86 a_13750_11850.n6 a_13750_11850.n5 0.96925
R87 VGND.n1492 VGND.n845 2.15834e+06
R88 VGND.n843 VGND.n84 538609
R89 VGND.n1342 VGND.n845 462138
R90 VGND.n1355 VGND.n1342 132103
R91 VGND.n1492 VGND.n1491 132000
R92 VGND.n843 VGND.n842 74151.2
R93 VGND.n1378 VGND.n931 41071.3
R94 VGND.n1280 VGND.n83 30967.2
R95 VGND.n1439 VGND.n1438 24590
R96 VGND.n1440 VGND.n1439 17800
R97 VGND.n1363 VGND.n1338 17400
R98 VGND.n1491 VGND.t168 16643.9
R99 VGND.n2415 VGND.n2414 16025.7
R100 VGND.n1338 VGND.n840 15708.2
R101 VGND.n1369 VGND.n1280 14498.6
R102 VGND.n1015 VGND.n989 14177.8
R103 VGND.n1280 VGND.n1279 11369.3
R104 VGND.n1344 VGND.n846 11368.8
R105 VGND.n1491 VGND.n846 9777.78
R106 VGND.n1494 VGND.n840 9511.11
R107 VGND.n899 VGND.n887 8988.12
R108 VGND.n899 VGND.n885 8938.88
R109 VGND.n1494 VGND.n1493 8900
R110 VGND.n858 VGND.n846 8134.99
R111 VGND.n1438 VGND.n1437 7550
R112 VGND.n927 VGND.n887 7116.62
R113 VGND.n927 VGND.n885 7067.38
R114 VGND.t190 VGND.n784 7029.52
R115 VGND.n2414 VGND.n2413 6982.65
R116 VGND.n1437 VGND.n1436 6150.9
R117 VGND.n2465 VGND.n2464 5527.06
R118 VGND.n2467 VGND.n2461 5527.06
R119 VGND.n46 VGND.n44 5527.06
R120 VGND.n49 VGND.n43 5527.06
R121 VGND.n2507 VGND.n2501 5230.59
R122 VGND.n2505 VGND.n2504 5230.59
R123 VGND.n1439 VGND.n884 5000.6
R124 VGND.n844 VGND.n785 4952.55
R125 VGND.n929 VGND.n928 4855.96
R126 VGND.n1345 VGND.n845 4738.46
R127 VGND.n2477 VGND.n2475 4595.29
R128 VGND.n2480 VGND.n2474 4595.29
R129 VGND.n1015 VGND.n884 4410.82
R130 VGND.t218 VGND.n1494 4106.67
R131 VGND.n1341 VGND.n840 4106.67
R132 VGND.n1380 VGND.n1379 3944.94
R133 VGND.n1377 VGND.n1376 3572.31
R134 VGND.n2493 VGND.n2492 3300
R135 VGND.n2490 VGND.n2488 3300
R136 VGND.n25 VGND.n24 3300
R137 VGND.n22 VGND.n20 3300
R138 VGND.n1378 VGND.n1377 3125.57
R139 VGND.n1290 VGND.n1289 2978.82
R140 VGND.n1287 VGND.n1285 2978.82
R141 VGND.n2414 VGND.n83 2975.62
R142 VGND.n36 VGND.n30 2929.41
R143 VGND.n34 VGND.n33 2929.41
R144 VGND.n1007 VGND.n1005 2880
R145 VGND.n1010 VGND.n1004 2880
R146 VGND.n1436 VGND.n931 2645.5
R147 VGND.t280 VGND.n785 2478.56
R148 VGND.n1376 VGND.n929 2412.14
R149 VGND.n1493 VGND.n1492 2386.9
R150 VGND.n1338 VGND.t283 2350.42
R151 VGND.n1400 VGND.n1015 2236.98
R152 VGND.t190 VGND.n785 2042.86
R153 VGND.n2046 VGND.n97 1770.48
R154 VGND.t218 VGND.n361 1770.48
R155 VGND.n2504 VGND.n2503 1636.97
R156 VGND.n2507 VGND.n2506 1636.97
R157 VGND.t214 VGND.n1024 1410.87
R158 VGND.n1379 VGND.n1378 1394.75
R159 VGND.n1272 VGND.n1018 1365.52
R160 VGND.n1272 VGND.n1271 1365.52
R161 VGND.n1271 VGND.n1270 1365.52
R162 VGND.n1270 VGND.n1124 1365.52
R163 VGND.n1264 VGND.n1263 1365.52
R164 VGND.n1263 VGND.n1262 1365.52
R165 VGND.n1262 VGND.n1128 1365.52
R166 VGND.n1256 VGND.n1128 1365.52
R167 VGND.n1256 VGND.n1255 1365.52
R168 VGND.n1465 VGND.n1464 1217.93
R169 VGND.n1453 VGND.n1452 1217.93
R170 VGND.n1451 VGND.n1450 1217.93
R171 VGND.n192 VGND.n69 1214.72
R172 VGND.n198 VGND.n192 1214.72
R173 VGND.n199 VGND.n198 1214.72
R174 VGND.n199 VGND.n188 1214.72
R175 VGND.n205 VGND.n188 1214.72
R176 VGND.n207 VGND.n184 1214.72
R177 VGND.n213 VGND.n184 1214.72
R178 VGND.n213 VGND.n180 1214.72
R179 VGND.n219 VGND.n180 1214.72
R180 VGND.n220 VGND.n219 1214.72
R181 VGND.n1412 VGND.n1411 1186
R182 VGND.n993 VGND.n977 1186
R183 VGND.n939 VGND.n938 1186
R184 VGND.n1436 VGND.n1435 1186
R185 VGND.n1490 VGND.n1489 1182.8
R186 VGND.n1467 VGND.n1466 1182.8
R187 VGND.n2389 VGND.n97 1162.86
R188 VGND.t218 VGND.n362 1162.86
R189 VGND.n1279 VGND.n1018 1092.41
R190 VGND.n1400 VGND.n1016 1090.76
R191 VGND.t8 VGND.t4 1054.97
R192 VGND.t191 VGND.t285 1054.97
R193 VGND.n2407 VGND.n88 942.857
R194 VGND.n2407 VGND.n2406 942.857
R195 VGND.n2406 VGND.n2405 942.857
R196 VGND.n2405 VGND.n89 942.857
R197 VGND.n2399 VGND.n2398 942.857
R198 VGND.n2398 VGND.n2397 942.857
R199 VGND.n2397 VGND.n93 942.857
R200 VGND.n2391 VGND.n93 942.857
R201 VGND.n2391 VGND.n2390 942.857
R202 VGND.n2390 VGND.n2389 942.857
R203 VGND.n2046 VGND.n2045 942.857
R204 VGND.n2045 VGND.n2044 942.857
R205 VGND.n2044 VGND.n2035 942.857
R206 VGND.n2038 VGND.n2035 942.857
R207 VGND.n2038 VGND.n370 942.857
R208 VGND.n2331 VGND.n371 942.857
R209 VGND.n2325 VGND.n371 942.857
R210 VGND.n2325 VGND.n2324 942.857
R211 VGND.n2324 VGND.n2323 942.857
R212 VGND.n2323 VGND.n377 942.857
R213 VGND.n377 VGND.n362 942.857
R214 VGND.n1657 VGND.n361 942.857
R215 VGND.n1693 VGND.n1657 942.857
R216 VGND.n1694 VGND.n1693 942.857
R217 VGND.n1695 VGND.n1694 942.857
R218 VGND.n1695 VGND.n754 942.857
R219 VGND.n1652 VGND.n755 942.857
R220 VGND.n1703 VGND.n1652 942.857
R221 VGND.n1704 VGND.n1703 942.857
R222 VGND.n1706 VGND.n1704 942.857
R223 VGND.n1706 VGND.n1705 942.857
R224 VGND.n1705 VGND.n784 942.857
R225 VGND.n1124 VGND.t214 925.518
R226 VGND.n884 VGND.t302 912.245
R227 VGND.n205 VGND.t214 823.313
R228 VGND.t10 VGND.t325 790.419
R229 VGND.n1100 VGND.t214 764.684
R230 VGND.n2440 VGND.n2439 764.684
R231 VGND.n842 VGND.n88 754.287
R232 VGND.n1094 VGND.t214 748.327
R233 VGND.n2439 VGND.n2438 748.327
R234 VGND.n903 VGND.t328 741.635
R235 VGND.n892 VGND.t327 741.635
R236 VGND.n916 VGND.t332 741.635
R237 VGND.n1377 VGND.n83 736
R238 VGND.n1118 VGND.n1023 717.391
R239 VGND.n1118 VGND.n1117 717.391
R240 VGND.n1117 VGND.n1116 717.391
R241 VGND.n2467 VGND.n2466 690.328
R242 VGND.n2464 VGND.n2463 690.328
R243 VGND.n47 VGND.n43 690.328
R244 VGND.n48 VGND.n44 690.328
R245 VGND.n1312 VGND.n1311 686.717
R246 VGND.n1331 VGND.n1330 686.717
R247 VGND.n1336 VGND.n1335 686.717
R248 VGND.n1336 VGND.n1281 686.717
R249 VGND.n1323 VGND.n1322 686.717
R250 VGND.n1304 VGND.n1303 686.717
R251 VGND.t6 VGND.t47 683.713
R252 VGND.t218 VGND.t16 677.36
R253 VGND.n2478 VGND.n2474 672.937
R254 VGND.n2479 VGND.n2475 672.937
R255 VGND.n1398 VGND.n1397 669.307
R256 VGND.n1415 VGND.n1414 669.307
R257 VGND.n988 VGND.n979 669.307
R258 VGND.n1425 VGND.n1424 669.307
R259 VGND.n946 VGND.n940 669.307
R260 VGND.n965 VGND.n964 669.307
R261 VGND.n961 VGND.n955 669.307
R262 VGND.n1637 VGND.n1636 669.307
R263 VGND.n1623 VGND.n1622 669.307
R264 VGND.n2456 VGND.n2455 654.447
R265 VGND.t214 VGND.n89 639.048
R266 VGND.t218 VGND.n370 639.048
R267 VGND.t218 VGND.n754 639.048
R268 VGND.n886 VGND.t180 638.923
R269 VGND.t77 VGND.t70 628.572
R270 VGND.t14 VGND.t138 628.572
R271 VGND.n2468 VGND.n2460 589.553
R272 VGND.n2462 VGND.n2460 589.553
R273 VGND.n2462 VGND.n2459 589.553
R274 VGND.n50 VGND.n42 589.553
R275 VGND.n45 VGND.n42 589.553
R276 VGND.n45 VGND.n41 589.553
R277 VGND.n1364 VGND.n1363 585.003
R278 VGND.n861 VGND.n859 585.003
R279 VGND.n1354 VGND.n1353 585.003
R280 VGND.n1360 VGND.n1359 585.001
R281 VGND.n1362 VGND.n1361 585.001
R282 VGND.n1344 VGND.n1343 585.001
R283 VGND.n1356 VGND.n1355 585.001
R284 VGND.n1374 VGND.n1373 585.001
R285 VGND.n1371 VGND.n1370 585.001
R286 VGND.n1368 VGND.n1367 585.001
R287 VGND.n1402 VGND.n1401 585.001
R288 VGND.n1429 VGND.n1427 585.001
R289 VGND.n883 VGND.n882 585.001
R290 VGND.n880 VGND.n879 585.001
R291 VGND.n878 VGND.n877 585.001
R292 VGND.n876 VGND.n875 585.001
R293 VGND.n872 VGND.n871 585.001
R294 VGND.n870 VGND.n869 585.001
R295 VGND.n868 VGND.n867 585.001
R296 VGND.n858 VGND.n857 585.001
R297 VGND.n1115 VGND.n1114 585
R298 VGND.n1116 VGND.n1115 585
R299 VGND.n1022 VGND.n1021 585
R300 VGND.n1117 VGND.n1022 585
R301 VGND.n1120 VGND.n1119 585
R302 VGND.n1119 VGND.n1118 585
R303 VGND.n1121 VGND.n1019 585
R304 VGND.n1023 VGND.n1019 585
R305 VGND.n1275 VGND.n1020 585
R306 VGND.n1020 VGND.n1018 585
R307 VGND.n1274 VGND.n1273 585
R308 VGND.n1273 VGND.n1272 585
R309 VGND.n1123 VGND.n1122 585
R310 VGND.n1271 VGND.n1123 585
R311 VGND.n1269 VGND.n1268 585
R312 VGND.n1270 VGND.n1269 585
R313 VGND.n1267 VGND.n1125 585
R314 VGND.n1125 VGND.n1124 585
R315 VGND.n1266 VGND.n1265 585
R316 VGND.n1265 VGND.n1264 585
R317 VGND.n1127 VGND.n1126 585
R318 VGND.n1263 VGND.n1127 585
R319 VGND.n1261 VGND.n1260 585
R320 VGND.n1262 VGND.n1261 585
R321 VGND.n1259 VGND.n1129 585
R322 VGND.n1129 VGND.n1128 585
R323 VGND.n1258 VGND.n1257 585
R324 VGND.n1257 VGND.n1256 585
R325 VGND.n1255 VGND.n1254 585
R326 VGND.n1277 VGND.n1276 585
R327 VGND.n1278 VGND.n1277 585
R328 VGND.n1992 VGND.n1991 585
R329 VGND.n1990 VGND.n658 585
R330 VGND.n1989 VGND.n1988 585
R331 VGND.n1987 VGND.n1986 585
R332 VGND.n1985 VGND.n1984 585
R333 VGND.n1983 VGND.n1982 585
R334 VGND.n1981 VGND.n1980 585
R335 VGND.n1979 VGND.n1978 585
R336 VGND.n1977 VGND.n1976 585
R337 VGND.n1975 VGND.n1974 585
R338 VGND.n1973 VGND.n653 585
R339 VGND.n1994 VGND.n653 585
R340 VGND.n1972 VGND.n661 585
R341 VGND.n1972 VGND.n1971 585
R342 VGND.n2165 VGND.n1994 585
R343 VGND.n2143 VGND.n2142 585
R344 VGND.n2144 VGND.n1999 585
R345 VGND.n2146 VGND.n2145 585
R346 VGND.n2148 VGND.n1998 585
R347 VGND.n2151 VGND.n2150 585
R348 VGND.n2152 VGND.n1997 585
R349 VGND.n2154 VGND.n2153 585
R350 VGND.n2156 VGND.n1996 585
R351 VGND.n2159 VGND.n2158 585
R352 VGND.n2160 VGND.n1995 585
R353 VGND.n2162 VGND.n2161 585
R354 VGND.n2119 VGND.n350 585
R355 VGND.n2122 VGND.n2121 585
R356 VGND.n2124 VGND.n2123 585
R357 VGND.n2126 VGND.n2117 585
R358 VGND.n2128 VGND.n2127 585
R359 VGND.n2129 VGND.n2116 585
R360 VGND.n2131 VGND.n2130 585
R361 VGND.n2133 VGND.n2114 585
R362 VGND.n2135 VGND.n2134 585
R363 VGND.n2136 VGND.n2113 585
R364 VGND.n2138 VGND.n2137 585
R365 VGND.n2140 VGND.n2000 585
R366 VGND.n2110 VGND.n2109 585
R367 VGND.n2032 VGND.n2012 585
R368 VGND.n2031 VGND.n2030 585
R369 VGND.n2029 VGND.n2028 585
R370 VGND.n2027 VGND.n2026 585
R371 VGND.n2025 VGND.n2024 585
R372 VGND.n2023 VGND.n2022 585
R373 VGND.n2021 VGND.n2020 585
R374 VGND.n2019 VGND.n2018 585
R375 VGND.n2017 VGND.n2016 585
R376 VGND.n2015 VGND.n2014 585
R377 VGND.n353 VGND.n349 585
R378 VGND.n2049 VGND.n2048 585
R379 VGND.n2051 VGND.n2050 585
R380 VGND.n2053 VGND.n2052 585
R381 VGND.n2055 VGND.n2054 585
R382 VGND.n2057 VGND.n2056 585
R383 VGND.n2059 VGND.n2058 585
R384 VGND.n2061 VGND.n2060 585
R385 VGND.n2063 VGND.n2062 585
R386 VGND.n2065 VGND.n2064 585
R387 VGND.n2067 VGND.n2066 585
R388 VGND.n2069 VGND.n2068 585
R389 VGND.n2072 VGND.n2070 585
R390 VGND.n2339 VGND.n224 585
R391 VGND.n1251 VGND.n1250 585
R392 VGND.n1248 VGND.n1247 585
R393 VGND.n1132 VGND.n1131 585
R394 VGND.n1242 VGND.n1241 585
R395 VGND.n1239 VGND.n1238 585
R396 VGND.n1160 VGND.n1137 585
R397 VGND.n1163 VGND.n1162 585
R398 VGND.n1166 VGND.n1158 585
R399 VGND.n1172 VGND.n1171 585
R400 VGND.n1174 VGND.n1157 585
R401 VGND.n1179 VGND.n1178 585
R402 VGND.n1176 VGND.n1175 585
R403 VGND.n347 VGND.n226 585
R404 VGND.n345 VGND.n344 585
R405 VGND.n342 VGND.n341 585
R406 VGND.n257 VGND.n230 585
R407 VGND.n260 VGND.n259 585
R408 VGND.n263 VGND.n262 585
R409 VGND.n256 VGND.n252 585
R410 VGND.n268 VGND.n251 585
R411 VGND.n274 VGND.n273 585
R412 VGND.n276 VGND.n250 585
R413 VGND.n281 VGND.n280 585
R414 VGND.n278 VGND.n277 585
R415 VGND.n1686 VGND.n1659 585
R416 VGND.n1684 VGND.n1683 585
R417 VGND.n1682 VGND.n1660 585
R418 VGND.n1681 VGND.n1680 585
R419 VGND.n1678 VGND.n1661 585
R420 VGND.n1676 VGND.n1675 585
R421 VGND.n1674 VGND.n1662 585
R422 VGND.n1673 VGND.n1672 585
R423 VGND.n1670 VGND.n1663 585
R424 VGND.n1668 VGND.n1667 585
R425 VGND.n1666 VGND.n1665 585
R426 VGND.n747 VGND.n745 585
R427 VGND.n2168 VGND.n2167 585
R428 VGND.n2169 VGND.n588 585
R429 VGND.n2179 VGND.n2178 585
R430 VGND.n2181 VGND.n587 585
R431 VGND.n2184 VGND.n2183 585
R432 VGND.n2185 VGND.n583 585
R433 VGND.n2194 VGND.n2193 585
R434 VGND.n2196 VGND.n582 585
R435 VGND.n2199 VGND.n2198 585
R436 VGND.n2200 VGND.n576 585
R437 VGND.n2209 VGND.n2208 585
R438 VGND.n2211 VGND.n575 585
R439 VGND.n2219 VGND.n2218 585
R440 VGND.n2220 VGND.n476 585
R441 VGND.n2230 VGND.n2229 585
R442 VGND.n2232 VGND.n475 585
R443 VGND.n2235 VGND.n2234 585
R444 VGND.n2236 VGND.n471 585
R445 VGND.n2245 VGND.n2244 585
R446 VGND.n2247 VGND.n470 585
R447 VGND.n2250 VGND.n2249 585
R448 VGND.n2251 VGND.n464 585
R449 VGND.n2260 VGND.n2259 585
R450 VGND.n2262 VGND.n463 585
R451 VGND.n2274 VGND.n2273 585
R452 VGND.n2275 VGND.n393 585
R453 VGND.n2285 VGND.n2284 585
R454 VGND.n2287 VGND.n392 585
R455 VGND.n2290 VGND.n2289 585
R456 VGND.n2291 VGND.n388 585
R457 VGND.n2300 VGND.n2299 585
R458 VGND.n2302 VGND.n387 585
R459 VGND.n2305 VGND.n2304 585
R460 VGND.n2306 VGND.n381 585
R461 VGND.n2315 VGND.n2314 585
R462 VGND.n2317 VGND.n379 585
R463 VGND.n1813 VGND.n1812 585
R464 VGND.n1815 VGND.n743 585
R465 VGND.n1818 VGND.n1817 585
R466 VGND.n1819 VGND.n742 585
R467 VGND.n1821 VGND.n1820 585
R468 VGND.n1823 VGND.n741 585
R469 VGND.n1826 VGND.n1825 585
R470 VGND.n1827 VGND.n740 585
R471 VGND.n1829 VGND.n1828 585
R472 VGND.n1831 VGND.n739 585
R473 VGND.n1833 VGND.n1832 585
R474 VGND.n1835 VGND.n1834 585
R475 VGND.n736 VGND.n709 585
R476 VGND.n735 VGND.n734 585
R477 VGND.n732 VGND.n710 585
R478 VGND.n730 VGND.n729 585
R479 VGND.n728 VGND.n711 585
R480 VGND.n727 VGND.n726 585
R481 VGND.n724 VGND.n712 585
R482 VGND.n722 VGND.n721 585
R483 VGND.n720 VGND.n713 585
R484 VGND.n719 VGND.n718 585
R485 VGND.n716 VGND.n714 585
R486 VGND.n660 VGND.n659 585
R487 VGND.n697 VGND.n692 585
R488 VGND.n1868 VGND.n1867 585
R489 VGND.n1865 VGND.n700 585
R490 VGND.n1863 VGND.n1862 585
R491 VGND.n702 VGND.n701 585
R492 VGND.n1856 VGND.n1855 585
R493 VGND.n1853 VGND.n704 585
R494 VGND.n1851 VGND.n1850 585
R495 VGND.n706 VGND.n705 585
R496 VGND.n1844 VGND.n1843 585
R497 VGND.n1841 VGND.n708 585
R498 VGND.n1839 VGND.n1838 585
R499 VGND.n1838 VGND.n1837 585
R500 VGND.n708 VGND.n707 585
R501 VGND.n1845 VGND.n1844 585
R502 VGND.n1847 VGND.n706 585
R503 VGND.n1850 VGND.n1849 585
R504 VGND.n704 VGND.n703 585
R505 VGND.n1857 VGND.n1856 585
R506 VGND.n1859 VGND.n702 585
R507 VGND.n1862 VGND.n1861 585
R508 VGND.n700 VGND.n699 585
R509 VGND.n1869 VGND.n1868 585
R510 VGND.n1871 VGND.n697 585
R511 VGND.n2214 VGND.n2213 585
R512 VGND.n573 VGND.n541 585
R513 VGND.n572 VGND.n571 585
R514 VGND.n568 VGND.n565 585
R515 VGND.n564 VGND.n543 585
R516 VGND.n562 VGND.n561 585
R517 VGND.n558 VGND.n544 585
R518 VGND.n557 VGND.n554 585
R519 VGND.n552 VGND.n545 585
R520 VGND.n550 VGND.n549 585
R521 VGND.n547 VGND.n352 585
R522 VGND.n2335 VGND.n351 585
R523 VGND.n2212 VGND.n540 585
R524 VGND.n2212 VGND.n457 585
R525 VGND.n2335 VGND.n2334 585
R526 VGND.n354 VGND.n352 585
R527 VGND.n549 VGND.n548 585
R528 VGND.n555 VGND.n545 585
R529 VGND.n557 VGND.n556 585
R530 VGND.n559 VGND.n558 585
R531 VGND.n561 VGND.n560 585
R532 VGND.n566 VGND.n543 585
R533 VGND.n568 VGND.n567 585
R534 VGND.n571 VGND.n570 585
R535 VGND.n569 VGND.n541 585
R536 VGND.n2215 VGND.n2214 585
R537 VGND.n2216 VGND.n540 585
R538 VGND.n2216 VGND.n457 585
R539 VGND.n2337 VGND.n223 585
R540 VGND.n2339 VGND.n223 585
R541 VGND.n2338 VGND.n2337 585
R542 VGND.n2339 VGND.n2338 585
R543 VGND.n1061 VGND.n1060 585
R544 VGND.n1062 VGND.n1051 585
R545 VGND.n1065 VGND.n1050 585
R546 VGND.n1066 VGND.n1049 585
R547 VGND.n1069 VGND.n1048 585
R548 VGND.n1070 VGND.n1047 585
R549 VGND.n1073 VGND.n1046 585
R550 VGND.n1075 VGND.n1045 585
R551 VGND.n1076 VGND.n1044 585
R552 VGND.n1077 VGND.n1043 585
R553 VGND.n1052 VGND.n1042 585
R554 VGND.n1034 VGND.n1033 585
R555 VGND.n1082 VGND.n1034 585
R556 VGND.n1042 VGND.n1036 585
R557 VGND.n1078 VGND.n1077 585
R558 VGND.n1076 VGND.n1041 585
R559 VGND.n1075 VGND.n1074 585
R560 VGND.n1073 VGND.n1072 585
R561 VGND.n1071 VGND.n1070 585
R562 VGND.n1069 VGND.n1068 585
R563 VGND.n1067 VGND.n1066 585
R564 VGND.n1065 VGND.n1064 585
R565 VGND.n1063 VGND.n1062 585
R566 VGND.n1061 VGND.n225 585
R567 VGND.n1099 VGND.n1098 585
R568 VGND.n1100 VGND.n1099 585
R569 VGND.n1032 VGND.n1031 585
R570 VGND.n1101 VGND.n1032 585
R571 VGND.n1104 VGND.n1103 585
R572 VGND.n1103 VGND.n1102 585
R573 VGND.n1105 VGND.n1030 585
R574 VGND.n1030 VGND.n1029 585
R575 VGND.n1107 VGND.n1106 585
R576 VGND.n1108 VGND.n1107 585
R577 VGND.n1027 VGND.n1026 585
R578 VGND.n1109 VGND.n1027 585
R579 VGND.n1112 VGND.n1111 585
R580 VGND.n1111 VGND.n1110 585
R581 VGND.n1113 VGND.n1025 585
R582 VGND.n1028 VGND.n1025 585
R583 VGND.n57 VGND.n56 585
R584 VGND.n2454 VGND.n2453 585
R585 VGND.t214 VGND.n2454 585
R586 VGND.n1705 VGND.n1651 585
R587 VGND.n1708 VGND.n1707 585
R588 VGND.n1707 VGND.n1706 585
R589 VGND.n1650 VGND.n1649 585
R590 VGND.n1704 VGND.n1650 585
R591 VGND.n1702 VGND.n1701 585
R592 VGND.n1703 VGND.n1702 585
R593 VGND.n1700 VGND.n1653 585
R594 VGND.n1653 VGND.n1652 585
R595 VGND.n1699 VGND.n1698 585
R596 VGND.n1698 VGND.n755 585
R597 VGND.n1697 VGND.n1654 585
R598 VGND.n1697 VGND.n754 585
R599 VGND.n1696 VGND.n1656 585
R600 VGND.n1696 VGND.n1695 585
R601 VGND.n1690 VGND.n1655 585
R602 VGND.n1694 VGND.n1655 585
R603 VGND.n1692 VGND.n1691 585
R604 VGND.n1693 VGND.n1692 585
R605 VGND.n1689 VGND.n1658 585
R606 VGND.n1658 VGND.n1657 585
R607 VGND.n1688 VGND.n1687 585
R608 VGND.n1687 VGND.n361 585
R609 VGND.n1647 VGND.n784 585
R610 VGND.n378 VGND.n377 585
R611 VGND.n2322 VGND.n2321 585
R612 VGND.n2323 VGND.n2322 585
R613 VGND.n376 VGND.n375 585
R614 VGND.n2324 VGND.n376 585
R615 VGND.n2327 VGND.n2326 585
R616 VGND.n2326 VGND.n2325 585
R617 VGND.n2328 VGND.n373 585
R618 VGND.n373 VGND.n371 585
R619 VGND.n2330 VGND.n2329 585
R620 VGND.n2331 VGND.n2330 585
R621 VGND.n374 VGND.n372 585
R622 VGND.n372 VGND.n370 585
R623 VGND.n2040 VGND.n2039 585
R624 VGND.n2039 VGND.n2038 585
R625 VGND.n2041 VGND.n2036 585
R626 VGND.n2036 VGND.n2035 585
R627 VGND.n2043 VGND.n2042 585
R628 VGND.n2044 VGND.n2043 585
R629 VGND.n2037 VGND.n2034 585
R630 VGND.n2045 VGND.n2034 585
R631 VGND.n2047 VGND.n2033 585
R632 VGND.n2047 VGND.n2046 585
R633 VGND.n2318 VGND.n362 585
R634 VGND.n2390 VGND.n96 585
R635 VGND.n2389 VGND.n2388 585
R636 VGND.n2343 VGND.n2342 585
R637 VGND.n2344 VGND.n112 585
R638 VGND.n2354 VGND.n2353 585
R639 VGND.n2356 VGND.n111 585
R640 VGND.n2359 VGND.n2358 585
R641 VGND.n2360 VGND.n107 585
R642 VGND.n2369 VGND.n2368 585
R643 VGND.n2371 VGND.n106 585
R644 VGND.n2374 VGND.n2373 585
R645 VGND.n2375 VGND.n100 585
R646 VGND.n2384 VGND.n2383 585
R647 VGND.n2386 VGND.n98 585
R648 VGND.n2393 VGND.n2392 585
R649 VGND.n2392 VGND.n2391 585
R650 VGND.n2394 VGND.n94 585
R651 VGND.n94 VGND.n93 585
R652 VGND.n2396 VGND.n2395 585
R653 VGND.n2397 VGND.n2396 585
R654 VGND.n92 VGND.n91 585
R655 VGND.n2398 VGND.n92 585
R656 VGND.n2401 VGND.n2400 585
R657 VGND.n2400 VGND.n2399 585
R658 VGND.n2402 VGND.n90 585
R659 VGND.n90 VGND.n89 585
R660 VGND.n2404 VGND.n2403 585
R661 VGND.n2405 VGND.n2404 585
R662 VGND.n87 VGND.n86 585
R663 VGND.n2406 VGND.n87 585
R664 VGND.n2409 VGND.n2408 585
R665 VGND.n2408 VGND.n2407 585
R666 VGND.n2410 VGND.n85 585
R667 VGND.n88 VGND.n85 585
R668 VGND.n2412 VGND.n2411 585
R669 VGND.n2413 VGND.n2412 585
R670 VGND.n82 VGND.n81 585
R671 VGND.n2415 VGND.n82 585
R672 VGND.n2418 VGND.n2417 585
R673 VGND.n2417 VGND.n2416 585
R674 VGND.n2419 VGND.n80 585
R675 VGND.n80 VGND.n79 585
R676 VGND.n2421 VGND.n2420 585
R677 VGND.n2422 VGND.n2421 585
R678 VGND.n78 VGND.n77 585
R679 VGND.n2423 VGND.n78 585
R680 VGND.n2426 VGND.n2425 585
R681 VGND.n2425 VGND.n2424 585
R682 VGND.n2427 VGND.n76 585
R683 VGND.n76 VGND.n75 585
R684 VGND.n2429 VGND.n2428 585
R685 VGND.n2430 VGND.n2429 585
R686 VGND.n74 VGND.n73 585
R687 VGND.n2431 VGND.n74 585
R688 VGND.n2434 VGND.n2433 585
R689 VGND.n2433 VGND.n2432 585
R690 VGND.n2435 VGND.n72 585
R691 VGND.n72 VGND.n70 585
R692 VGND.n2437 VGND.n2436 585
R693 VGND.n2438 VGND.n2437 585
R694 VGND.n2442 VGND.n2441 585
R695 VGND.n2441 VGND.n2440 585
R696 VGND.n2443 VGND.n65 585
R697 VGND.n65 VGND.n64 585
R698 VGND.n2445 VGND.n2444 585
R699 VGND.n2446 VGND.n2445 585
R700 VGND.n66 VGND.n63 585
R701 VGND.n2447 VGND.n63 585
R702 VGND.n2449 VGND.n61 585
R703 VGND.n2449 VGND.n2448 585
R704 VGND.n2451 VGND.n2450 585
R705 VGND.n2450 VGND.n59 585
R706 VGND.n62 VGND.n60 585
R707 VGND.n62 VGND.n58 585
R708 VGND.n1088 VGND.n1087 585
R709 VGND.n1087 VGND.n1086 585
R710 VGND.n1089 VGND.n1085 585
R711 VGND.n1085 VGND.n1084 585
R712 VGND.n1091 VGND.n1090 585
R713 VGND.n1092 VGND.n1091 585
R714 VGND.n1083 VGND.n1035 585
R715 VGND.n1093 VGND.n1083 585
R716 VGND.n1096 VGND.n1095 585
R717 VGND.n1095 VGND.n1094 585
R718 VGND.n221 VGND.n179 585
R719 VGND.n221 VGND.n220 585
R720 VGND.n217 VGND.n178 585
R721 VGND.n219 VGND.n178 585
R722 VGND.n216 VGND.n215 585
R723 VGND.n215 VGND.n180 585
R724 VGND.n214 VGND.n182 585
R725 VGND.n214 VGND.n213 585
R726 VGND.n210 VGND.n183 585
R727 VGND.n184 VGND.n183 585
R728 VGND.n209 VGND.n208 585
R729 VGND.n208 VGND.n207 585
R730 VGND.n206 VGND.n186 585
R731 VGND.n206 VGND.n205 585
R732 VGND.n202 VGND.n187 585
R733 VGND.n188 VGND.n187 585
R734 VGND.n201 VGND.n200 585
R735 VGND.n200 VGND.n199 585
R736 VGND.n191 VGND.n190 585
R737 VGND.n198 VGND.n191 585
R738 VGND.n195 VGND.n194 585
R739 VGND.n194 VGND.n192 585
R740 VGND.n193 VGND.n68 585
R741 VGND.n69 VGND.n68 585
R742 VGND.n222 VGND.n177 585
R743 VGND.n2339 VGND.n222 585
R744 VGND.n193 VGND.n71 585
R745 VGND.n71 VGND.n69 585
R746 VGND.n196 VGND.n195 585
R747 VGND.n196 VGND.n192 585
R748 VGND.n197 VGND.n190 585
R749 VGND.n198 VGND.n197 585
R750 VGND.n201 VGND.n189 585
R751 VGND.n199 VGND.n189 585
R752 VGND.n203 VGND.n202 585
R753 VGND.n203 VGND.n188 585
R754 VGND.n204 VGND.n186 585
R755 VGND.n205 VGND.n204 585
R756 VGND.n209 VGND.n185 585
R757 VGND.n207 VGND.n185 585
R758 VGND.n211 VGND.n210 585
R759 VGND.n211 VGND.n184 585
R760 VGND.n212 VGND.n182 585
R761 VGND.n213 VGND.n212 585
R762 VGND.n216 VGND.n181 585
R763 VGND.n181 VGND.n180 585
R764 VGND.n218 VGND.n217 585
R765 VGND.n219 VGND.n218 585
R766 VGND.n179 VGND.n176 585
R767 VGND.n220 VGND.n176 585
R768 VGND.n2340 VGND.n177 585
R769 VGND.n2340 VGND.n2339 585
R770 VGND.n2264 VGND.n459 585
R771 VGND.n2267 VGND.n2266 585
R772 VGND.n462 VGND.n461 585
R773 VGND.n2089 VGND.n2088 585
R774 VGND.n2094 VGND.n2086 585
R775 VGND.n2095 VGND.n2084 585
R776 VGND.n2096 VGND.n2083 585
R777 VGND.n2081 VGND.n2079 585
R778 VGND.n2101 VGND.n2078 585
R779 VGND.n2102 VGND.n2076 585
R780 VGND.n2075 VGND.n2071 585
R781 VGND.n2107 VGND.n2013 585
R782 VGND.n2263 VGND.n458 585
R783 VGND.n2263 VGND.n457 585
R784 VGND.n2107 VGND.n2106 585
R785 VGND.n2104 VGND.n2071 585
R786 VGND.n2103 VGND.n2102 585
R787 VGND.n2101 VGND.n2100 585
R788 VGND.n2099 VGND.n2079 585
R789 VGND.n2097 VGND.n2096 585
R790 VGND.n2095 VGND.n2080 585
R791 VGND.n2094 VGND.n2093 585
R792 VGND.n2091 VGND.n2089 585
R793 VGND.n461 VGND.n460 585
R794 VGND.n2268 VGND.n2267 585
R795 VGND.n2270 VGND.n459 585
R796 VGND.n2271 VGND.n458 585
R797 VGND.n2271 VGND.n457 585
R798 VGND.n791 VGND.n790 585
R799 VGND.n1527 VGND.n1526 585
R800 VGND.n1523 VGND.n1500 585
R801 VGND.n1522 VGND.n1519 585
R802 VGND.n1518 VGND.n1517 585
R803 VGND.n1516 VGND.n1513 585
R804 VGND.n1512 VGND.n1511 585
R805 VGND.n1510 VGND.n1507 585
R806 VGND.n1506 VGND.n1505 585
R807 VGND.n1504 VGND.n1502 585
R808 VGND.n1501 VGND.n746 585
R809 VGND.n1810 VGND.n744 585
R810 VGND.n1810 VGND.n1809 585
R811 VGND.n748 VGND.n746 585
R812 VGND.n1504 VGND.n1503 585
R813 VGND.n1508 VGND.n1505 585
R814 VGND.n1510 VGND.n1509 585
R815 VGND.n1514 VGND.n1511 585
R816 VGND.n1516 VGND.n1515 585
R817 VGND.n1520 VGND.n1517 585
R818 VGND.n1522 VGND.n1521 585
R819 VGND.n1524 VGND.n1523 585
R820 VGND.n1526 VGND.n1525 585
R821 VGND.n790 VGND.n789 585
R822 VGND.n1635 VGND.n795 585
R823 VGND.n1634 VGND.n794 585
R824 VGND.n1638 VGND.n794 585
R825 VGND.n1329 VGND.n1318 585
R826 VGND.n1328 VGND.n1327 585
R827 VGND.n1328 VGND.t212 585
R828 VGND.n1325 VGND.n1321 585
R829 VGND.n1310 VGND.n1309 585
R830 VGND.n1307 VGND.n1299 585
R831 VGND.n1299 VGND.t269 585
R832 VGND.n1302 VGND.n1300 585
R833 VGND.n1874 VGND.n1873 585
R834 VGND.n1875 VGND.n1874 585
R835 VGND.n1970 VGND.n662 585
R836 VGND.n1970 VGND.n365 585
R837 VGND.n1969 VGND.n664 585
R838 VGND.n1969 VGND.n1968 585
R839 VGND.n1957 VGND.n663 585
R840 VGND.n1967 VGND.n663 585
R841 VGND.n1965 VGND.n1964 585
R842 VGND.n1966 VGND.n1965 585
R843 VGND.n668 VGND.n666 585
R844 VGND.n666 VGND.n665 585
R845 VGND.n1884 VGND.n1883 585
R846 VGND.n1883 VGND.n366 585
R847 VGND.n1881 VGND.n1880 585
R848 VGND.n1880 VGND.n1879 585
R849 VGND.n1893 VGND.n1892 585
R850 VGND.n1894 VGND.n1893 585
R851 VGND.n689 VGND.n688 585
R852 VGND.n1895 VGND.n689 585
R853 VGND.n1898 VGND.n1897 585
R854 VGND.n1897 VGND.n1896 585
R855 VGND.n1878 VGND.n691 585
R856 VGND.n1878 VGND.n1877 585
R857 VGND.n693 VGND.n690 585
R858 VGND.n1876 VGND.n690 585
R859 VGND.n1642 VGND.n1641 585
R860 VGND.n1641 VGND.n1640 585
R861 VGND.n1873 VGND.n1872 585
R862 VGND.n1872 VGND.n695 585
R863 VGND.n809 VGND.n696 585
R864 VGND.n806 VGND.n696 585
R865 VGND.n1617 VGND.n1616 585
R866 VGND.n1618 VGND.n1617 585
R867 VGND.n811 VGND.n808 585
R868 VGND.n808 VGND.n807 585
R869 VGND.n1611 VGND.n1610 585
R870 VGND.n1610 VGND.n1609 585
R871 VGND.n817 VGND.n815 585
R872 VGND.n1608 VGND.n815 585
R873 VGND.n1606 VGND.n1605 585
R874 VGND.n1607 VGND.n1606 585
R875 VGND.n819 VGND.n816 585
R876 VGND.n1530 VGND.n816 585
R877 VGND.n1538 VGND.n1537 585
R878 VGND.n1539 VGND.n1538 585
R879 VGND.n1532 VGND.n839 585
R880 VGND.n1540 VGND.n839 585
R881 VGND.n1542 VGND.n838 585
R882 VGND.n1542 VGND.n1541 585
R883 VGND.n1544 VGND.n1543 585
R884 VGND.n1543 VGND.n793 585
R885 VGND.n792 VGND.n788 585
R886 VGND.n1639 VGND.n792 585
R887 VGND.n1642 VGND.n787 585
R888 VGND.n787 VGND.n786 585
R889 VGND.n1781 VGND.n1780 585
R890 VGND.n1782 VGND.n1781 585
R891 VGND.n782 VGND.n780 585
R892 VGND.n1783 VGND.n782 585
R893 VGND.n1797 VGND.n1796 585
R894 VGND.n1796 VGND.n1795 585
R895 VGND.n1785 VGND.n783 585
R896 VGND.n1794 VGND.n783 585
R897 VGND.n1792 VGND.n1791 585
R898 VGND.n1793 VGND.n1792 585
R899 VGND.n1787 VGND.n756 585
R900 VGND.n1784 VGND.n756 585
R901 VGND.n1805 VGND.n1804 585
R902 VGND.n1806 VGND.n1805 585
R903 VGND.n759 VGND.n757 585
R904 VGND.n1712 VGND.n757 585
R905 VGND.n1717 VGND.n1716 585
R906 VGND.n1718 VGND.n1717 585
R907 VGND.n1646 VGND.n1645 585
R908 VGND.n1719 VGND.n1646 585
R909 VGND.n1723 VGND.n1722 585
R910 VGND.n1722 VGND.n1721 585
R911 VGND.n1711 VGND.n1710 585
R912 VGND.n1720 VGND.n1711 585
R913 VGND.n1620 VGND.n1619 585
R914 VGND.n1621 VGND.n1620 585
R915 VGND.n805 VGND.n804 585
R916 VGND.n963 VGND.n957 585
R917 VGND.n962 VGND.n960 585
R918 VGND.n944 VGND.n941 585
R919 VGND.n951 VGND.n947 585
R920 VGND.n983 VGND.n976 585
R921 VGND.n987 VGND.n986 585
R922 VGND.n1389 VGND.n1383 585
R923 VGND.n1391 VGND.n1382 585
R924 VGND.n1399 VGND.n1382 585
R925 VGND.n1395 VGND.n1394 585
R926 VGND.n1394 VGND.n1016 585
R927 VGND.n900 VGND.n888 580.801
R928 VGND.n1278 VGND.t214 580.557
R929 VGND.n1255 VGND.t214 576.553
R930 VGND.n1017 VGND.t329 572.105
R931 VGND.n2508 VGND.n2502 557.929
R932 VGND.n2502 VGND.n2500 557.929
R933 VGND.n2509 VGND.n2508 549.271
R934 VGND.n2509 VGND.n2500 549.271
R935 VGND.n1380 VGND.t90 544.597
R936 VGND.n1379 VGND.n1375 538.591
R937 VGND.n1438 VGND.n929 534.261
R938 VGND.n1279 VGND.n1278 527.083
R939 VGND.n2469 VGND.n2459 518.777
R940 VGND.n51 VGND.n50 518.777
R941 VGND.n220 VGND.t214 512.884
R942 VGND.n1399 VGND.n1381 497.053
R943 VGND.n2481 VGND.n2473 490.166
R944 VGND.n2476 VGND.n2473 490.166
R945 VGND.n2476 VGND.n2472 490.166
R946 VGND.t198 VGND.t300 467.257
R947 VGND.n926 VGND.n888 459.2
R948 VGND.t150 VGND.t318 454.277
R949 VGND.t302 VGND.t296 444.599
R950 VGND.t146 VGND.t294 441.298
R951 VGND.n1264 VGND.t214 440
R952 VGND.n878 VGND.t35 436.935
R953 VGND.t206 VGND.t141 428.32
R954 VGND.t202 VGND.t140 428.32
R955 VGND.t43 VGND.t98 428.32
R956 VGND.t162 VGND.t119 428.32
R957 VGND.t118 VGND.t58 428.32
R958 VGND.t60 VGND.t83 428.32
R959 VGND.n1376 VGND.n931 420.812
R960 VGND.n2482 VGND.n2481 420.519
R961 VGND.n1490 VGND.t300 408.851
R962 VGND.n1116 VGND.n1024 398.551
R963 VGND.n207 VGND.t214 391.411
R964 VGND.n1110 VGND.n1028 368.031
R965 VGND.n1109 VGND.n1108 368.031
R966 VGND.n1108 VGND.n1029 368.031
R967 VGND.n1102 VGND.n1029 368.031
R968 VGND.n1102 VGND.n1101 368.031
R969 VGND.n1101 VGND.n1100 368.031
R970 VGND.n1094 VGND.n1093 368.031
R971 VGND.n1093 VGND.n1092 368.031
R972 VGND.n1092 VGND.n1084 368.031
R973 VGND.n1086 VGND.n1084 368.031
R974 VGND.n1086 VGND.n58 368.031
R975 VGND.n2448 VGND.n59 368.031
R976 VGND.n2448 VGND.n2447 368.031
R977 VGND.n2447 VGND.n2446 368.031
R978 VGND.n2446 VGND.n64 368.031
R979 VGND.n2440 VGND.n64 368.031
R980 VGND.n2438 VGND.n70 368.031
R981 VGND.n2432 VGND.n70 368.031
R982 VGND.n2432 VGND.n2431 368.031
R983 VGND.n2431 VGND.n2430 368.031
R984 VGND.n2430 VGND.n75 368.031
R985 VGND.n2424 VGND.n2423 368.031
R986 VGND.n2423 VGND.n2422 368.031
R987 VGND.n2422 VGND.n79 368.031
R988 VGND.n2416 VGND.n79 368.031
R989 VGND.n2416 VGND.n2415 368.031
R990 VGND.n883 VGND.t75 360.279
R991 VGND.n879 VGND.t25 360.279
R992 VGND.t270 VGND.n1440 356.933
R993 VGND.n2489 VGND.n2486 352
R994 VGND.n2489 VGND.n2485 352
R995 VGND.n21 VGND.n18 352
R996 VGND.n21 VGND.n17 352
R997 VGND.n1355 VGND.t85 347.368
R998 VGND.t320 VGND.n1354 347.368
R999 VGND.n1354 VGND.t316 347.368
R1000 VGND.n2494 VGND.n2486 343.558
R1001 VGND.n26 VGND.n18 343.558
R1002 VGND.n2495 VGND.n2485 342.966
R1003 VGND.n27 VGND.n17 342.966
R1004 VGND.t88 VGND.n1362 341.834
R1005 VGND.t115 VGND.n1360 341.834
R1006 VGND.n978 VGND.t260 336.329
R1007 VGND.n978 VGND.t250 336.329
R1008 VGND.n945 VGND.t243 336.329
R1009 VGND.n945 VGND.t223 336.329
R1010 VGND.n953 VGND.t227 330
R1011 VGND.n1387 VGND.t254 330
R1012 VGND.t218 VGND.n360 172.876
R1013 VGND.t218 VGND.n367 172.876
R1014 VGND.t218 VGND.n369 172.876
R1015 VGND.t218 VGND.n1529 172.876
R1016 VGND.t104 VGND.t198 324.485
R1017 VGND.t130 VGND.t95 324.485
R1018 VGND.t314 VGND.t307 324.485
R1019 VGND.t218 VGND.n698 172.615
R1020 VGND.t218 VGND.n368 172.615
R1021 VGND.n2332 VGND.t218 172.615
R1022 VGND.n1807 VGND.t218 172.615
R1023 VGND.n1286 VGND.n1282 317.741
R1024 VGND.n1286 VGND.n1283 317.741
R1025 VGND.n1291 VGND.n1283 317.741
R1026 VGND.n37 VGND.n29 312.471
R1027 VGND.n31 VGND.n29 312.471
R1028 VGND.n1477 VGND.t147 309.733
R1029 VGND.n1474 VGND.t301 309.733
R1030 VGND.n1473 VGND.t199 309.733
R1031 VGND.n1006 VGND.n1002 307.2
R1032 VGND.n1006 VGND.n1003 307.2
R1033 VGND.n1011 VGND.n1003 307.2
R1034 VGND.n1410 VGND.t219 304.634
R1035 VGND.n994 VGND.t247 304.634
R1036 VGND.n937 VGND.t238 304.634
R1037 VGND.n1434 VGND.t235 304.634
R1038 VGND.n31 VGND.n28 304.245
R1039 VGND.n2399 VGND.t214 303.81
R1040 VGND.t218 VGND.n2331 303.81
R1041 VGND.t218 VGND.n755 303.81
R1042 VGND.n38 VGND.n37 303.06
R1043 VGND.n876 VGND.t134 298.955
R1044 VGND.n871 VGND.t143 298.955
R1045 VGND.n1403 VGND.t231 292.584
R1046 VGND.n1430 VGND.t263 292.584
R1047 VGND.n898 VGND.n887 292.5
R1048 VGND.n887 VGND.n886 292.5
R1049 VGND.n888 VGND.n885 292.5
R1050 VGND.n886 VGND.n885 292.5
R1051 VGND.t106 VGND.n1451 292.036
R1052 VGND.n1452 VGND.t111 292.036
R1053 VGND.t171 VGND.n1465 292.036
R1054 VGND.t85 VGND.t8 283.041
R1055 VGND.t4 VGND.t320 283.041
R1056 VGND.t316 VGND.t191 283.041
R1057 VGND.t285 VGND.t144 283.041
R1058 VGND.n910 VGND.n900 273.601
R1059 VGND.n926 VGND.n925 270.401
R1060 VGND.n1253 VGND.n1252 264.301
R1061 VGND.n1994 VGND.n652 264.301
R1062 VGND.n2164 VGND.n651 264.301
R1063 VGND.n1709 VGND.n1648 264.301
R1064 VGND.n2320 VGND.n2319 264.301
R1065 VGND.n2387 VGND.n95 264.301
R1066 VGND.n1342 VGND.n1341 262.949
R1067 VGND.n5 VGND.n4 261.733
R1068 VGND.n1476 VGND.n1475 261.733
R1069 VGND.n1479 VGND.n1478 261.733
R1070 VGND.n1481 VGND.n1480 261.733
R1071 VGND.n1483 VGND.n1482 261.733
R1072 VGND.n1485 VGND.n1484 261.733
R1073 VGND.n1487 VGND.n1486 261.733
R1074 VGND.n1472 VGND.n1471 261.733
R1075 VGND.n1470 VGND.n1469 261.733
R1076 VGND.n848 VGND.n847 261.733
R1077 VGND.n1461 VGND.n1460 261.733
R1078 VGND.n1440 VGND.n851 260.753
R1079 VGND.n1463 VGND.n1462 260.514
R1080 VGND.n1335 VGND.t17 260
R1081 VGND.t17 VGND.n1281 260
R1082 VGND.n2441 VGND.n68 259.416
R1083 VGND.n1687 VGND.n1686 259.416
R1084 VGND.n2048 VGND.n2047 259.416
R1085 VGND.n2110 VGND.n2013 259.416
R1086 VGND.n1839 VGND.n709 259.416
R1087 VGND.n1099 VGND.n1033 259.416
R1088 VGND.n2119 VGND.n351 259.416
R1089 VGND.n1813 VGND.n744 259.416
R1090 VGND.n2412 VGND.n82 259.416
R1091 VGND.n1581 VGND.n835 258.334
R1092 VGND.n524 VGND.n482 258.334
R1093 VGND.n1762 VGND.n1761 258.334
R1094 VGND.n320 VGND.n319 258.334
R1095 VGND.n441 VGND.n399 258.334
R1096 VGND.n1938 VGND.n674 258.334
R1097 VGND.n1216 VGND.n1154 258.334
R1098 VGND.n636 VGND.n594 258.334
R1099 VGND.n160 VGND.n118 258.334
R1100 VGND.n2455 VGND.t214 257.779
R1101 VGND.n1994 VGND.n1993 254.34
R1102 VGND.n1994 VGND.n657 254.34
R1103 VGND.n1994 VGND.n656 254.34
R1104 VGND.n1994 VGND.n655 254.34
R1105 VGND.n1994 VGND.n654 254.34
R1106 VGND.n2141 VGND.n1994 254.34
R1107 VGND.n2147 VGND.n1994 254.34
R1108 VGND.n2149 VGND.n1994 254.34
R1109 VGND.n2155 VGND.n1994 254.34
R1110 VGND.n2157 VGND.n1994 254.34
R1111 VGND.n2163 VGND.n1994 254.34
R1112 VGND.n2120 VGND.n2112 254.34
R1113 VGND.n2125 VGND.n2112 254.34
R1114 VGND.n2118 VGND.n2112 254.34
R1115 VGND.n2132 VGND.n2112 254.34
R1116 VGND.n2115 VGND.n2112 254.34
R1117 VGND.n2139 VGND.n2112 254.34
R1118 VGND.n2112 VGND.n2111 254.34
R1119 VGND.n2112 VGND.n2011 254.34
R1120 VGND.n2112 VGND.n2010 254.34
R1121 VGND.n2112 VGND.n2009 254.34
R1122 VGND.n2112 VGND.n2008 254.34
R1123 VGND.n2112 VGND.n2007 254.34
R1124 VGND.n2112 VGND.n2006 254.34
R1125 VGND.n2112 VGND.n2005 254.34
R1126 VGND.n2112 VGND.n2004 254.34
R1127 VGND.n2112 VGND.n2003 254.34
R1128 VGND.n2112 VGND.n2002 254.34
R1129 VGND.n2112 VGND.n2001 254.34
R1130 VGND.n1249 VGND.n99 254.34
R1131 VGND.n1240 VGND.n99 254.34
R1132 VGND.n1136 VGND.n99 254.34
R1133 VGND.n1161 VGND.n99 254.34
R1134 VGND.n1173 VGND.n99 254.34
R1135 VGND.n1177 VGND.n99 254.34
R1136 VGND.n343 VGND.n99 254.34
R1137 VGND.n229 VGND.n99 254.34
R1138 VGND.n261 VGND.n99 254.34
R1139 VGND.n255 VGND.n99 254.34
R1140 VGND.n275 VGND.n99 254.34
R1141 VGND.n279 VGND.n99 254.34
R1142 VGND.n1685 VGND.n363 254.34
R1143 VGND.n1679 VGND.n363 254.34
R1144 VGND.n1677 VGND.n363 254.34
R1145 VGND.n1671 VGND.n363 254.34
R1146 VGND.n1669 VGND.n363 254.34
R1147 VGND.n1664 VGND.n363 254.34
R1148 VGND.n2166 VGND.n380 254.34
R1149 VGND.n2180 VGND.n380 254.34
R1150 VGND.n2182 VGND.n380 254.34
R1151 VGND.n2195 VGND.n380 254.34
R1152 VGND.n2197 VGND.n380 254.34
R1153 VGND.n2210 VGND.n380 254.34
R1154 VGND.n2217 VGND.n380 254.34
R1155 VGND.n2231 VGND.n380 254.34
R1156 VGND.n2233 VGND.n380 254.34
R1157 VGND.n2246 VGND.n380 254.34
R1158 VGND.n2248 VGND.n380 254.34
R1159 VGND.n2261 VGND.n380 254.34
R1160 VGND.n2272 VGND.n380 254.34
R1161 VGND.n2286 VGND.n380 254.34
R1162 VGND.n2288 VGND.n380 254.34
R1163 VGND.n2301 VGND.n380 254.34
R1164 VGND.n2303 VGND.n380 254.34
R1165 VGND.n2316 VGND.n380 254.34
R1166 VGND.n1814 VGND.n363 254.34
R1167 VGND.n1816 VGND.n363 254.34
R1168 VGND.n1822 VGND.n363 254.34
R1169 VGND.n1824 VGND.n363 254.34
R1170 VGND.n1830 VGND.n363 254.34
R1171 VGND.n738 VGND.n363 254.34
R1172 VGND.n733 VGND.n363 254.34
R1173 VGND.n731 VGND.n363 254.34
R1174 VGND.n725 VGND.n363 254.34
R1175 VGND.n723 VGND.n363 254.34
R1176 VGND.n717 VGND.n363 254.34
R1177 VGND.n715 VGND.n363 254.34
R1178 VGND.n1866 VGND.n360 254.34
R1179 VGND.n1864 VGND.n360 254.34
R1180 VGND.n1854 VGND.n360 254.34
R1181 VGND.n1852 VGND.n360 254.34
R1182 VGND.n1842 VGND.n360 254.34
R1183 VGND.n1840 VGND.n360 254.34
R1184 VGND.n1836 VGND.n698 254.34
R1185 VGND.n1846 VGND.n698 254.34
R1186 VGND.n1848 VGND.n698 254.34
R1187 VGND.n1858 VGND.n698 254.34
R1188 VGND.n1860 VGND.n698 254.34
R1189 VGND.n1870 VGND.n698 254.34
R1190 VGND.n574 VGND.n369 254.34
R1191 VGND.n542 VGND.n369 254.34
R1192 VGND.n563 VGND.n369 254.34
R1193 VGND.n553 VGND.n369 254.34
R1194 VGND.n551 VGND.n369 254.34
R1195 VGND.n546 VGND.n369 254.34
R1196 VGND.n2333 VGND.n2332 254.34
R1197 VGND.n2332 VGND.n359 254.34
R1198 VGND.n2332 VGND.n358 254.34
R1199 VGND.n2332 VGND.n357 254.34
R1200 VGND.n2332 VGND.n356 254.34
R1201 VGND.n2332 VGND.n355 254.34
R1202 VGND.n1059 VGND.n1058 254.34
R1203 VGND.n1058 VGND.n1057 254.34
R1204 VGND.n1058 VGND.n1056 254.34
R1205 VGND.n1058 VGND.n1055 254.34
R1206 VGND.n1058 VGND.n1054 254.34
R1207 VGND.n1058 VGND.n1053 254.34
R1208 VGND.n1081 VGND.n1080 254.34
R1209 VGND.n1080 VGND.n1079 254.34
R1210 VGND.n1080 VGND.n1040 254.34
R1211 VGND.n1080 VGND.n1039 254.34
R1212 VGND.n1080 VGND.n1038 254.34
R1213 VGND.n1080 VGND.n1037 254.34
R1214 VGND.n2341 VGND.n99 254.34
R1215 VGND.n2355 VGND.n99 254.34
R1216 VGND.n2357 VGND.n99 254.34
R1217 VGND.n2370 VGND.n99 254.34
R1218 VGND.n2372 VGND.n99 254.34
R1219 VGND.n2385 VGND.n99 254.34
R1220 VGND.n2265 VGND.n367 254.34
R1221 VGND.n2087 VGND.n367 254.34
R1222 VGND.n2085 VGND.n367 254.34
R1223 VGND.n2082 VGND.n367 254.34
R1224 VGND.n2077 VGND.n367 254.34
R1225 VGND.n2074 VGND.n367 254.34
R1226 VGND.n2105 VGND.n368 254.34
R1227 VGND.n2073 VGND.n368 254.34
R1228 VGND.n2098 VGND.n368 254.34
R1229 VGND.n2092 VGND.n368 254.34
R1230 VGND.n2090 VGND.n368 254.34
R1231 VGND.n2269 VGND.n368 254.34
R1232 VGND.n1529 VGND.n1528 254.34
R1233 VGND.n1529 VGND.n1499 254.34
R1234 VGND.n1529 VGND.n1498 254.34
R1235 VGND.n1529 VGND.n1497 254.34
R1236 VGND.n1529 VGND.n1496 254.34
R1237 VGND.n1529 VGND.n1495 254.34
R1238 VGND.n1808 VGND.n1807 254.34
R1239 VGND.n1807 VGND.n753 254.34
R1240 VGND.n1807 VGND.n752 254.34
R1241 VGND.n1807 VGND.n751 254.34
R1242 VGND.n1807 VGND.n750 254.34
R1243 VGND.n1807 VGND.n749 254.34
R1244 VGND.n1451 VGND.t200 253.097
R1245 VGND.n1452 VGND.t23 253.097
R1246 VGND.n1465 VGND.t173 253.097
R1247 VGND.n1466 VGND.t164 253.097
R1248 VGND.n1638 VGND.n1637 250.349
R1249 VGND.n1622 VGND.n1621 250.349
R1250 VGND.n964 VGND.n930 250.349
R1251 VGND.n961 VGND.n930 250.349
R1252 VGND.n1426 VGND.n1425 250.349
R1253 VGND.n1426 VGND.n940 250.349
R1254 VGND.n1414 VGND.n1413 250.349
R1255 VGND.n1413 VGND.n988 250.349
R1256 VGND.n1399 VGND.n1398 250.349
R1257 VGND.n1095 VGND.n1082 249.663
R1258 VGND.n1809 VGND.n747 249.663
R1259 VGND.n2106 VGND.n2072 249.663
R1260 VGND.n2334 VGND.n353 249.663
R1261 VGND.n1992 VGND.n659 249.663
R1262 VGND.n1277 VGND.n1019 249.663
R1263 VGND.n2142 VGND.n2140 249.663
R1264 VGND.n1837 VGND.n1835 249.663
R1265 VGND.n2437 VGND.n71 249.663
R1266 VGND.n1310 VGND.n1299 246.25
R1267 VGND.n1302 VGND.n1299 246.25
R1268 VGND.n1329 VGND.n1328 246.25
R1269 VGND.n1328 VGND.n1321 246.25
R1270 VGND.n1411 VGND.t222 245
R1271 VGND.n993 VGND.t249 245
R1272 VGND.n938 VGND.t241 245
R1273 VGND.n1435 VGND.t237 245
R1274 VGND.t94 VGND.n851 242.395
R1275 VGND.n1337 VGND.n1336 241.643
R1276 VGND.n1330 VGND.t212 241.643
R1277 VGND.n1322 VGND.t212 241.643
R1278 VGND.n1311 VGND.t269 241.643
R1279 VGND.n1303 VGND.t269 241.643
R1280 VGND.t296 VGND.n883 237.631
R1281 VGND.n879 VGND.t75 237.631
R1282 VGND.t25 VGND.n878 237.631
R1283 VGND.n1363 VGND.t88 236.654
R1284 VGND.n1362 VGND.t115 236.654
R1285 VGND.n1360 VGND.t132 236.654
R1286 VGND.n1443 VGND.n1441 233.793
R1287 VGND.n1489 VGND.t69 233
R1288 VGND.n1467 VGND.t187 233
R1289 VGND.n1459 VGND.n1458 232.934
R1290 VGND.n1457 VGND.n1456 232.934
R1291 VGND.n1455 VGND.n1454 232.934
R1292 VGND.n850 VGND.n849 232.934
R1293 VGND.n1447 VGND.n1446 232.934
R1294 VGND.n1449 VGND.n1448 232.934
R1295 VGND.n1445 VGND.n1444 232.934
R1296 VGND.n1443 VGND.n1442 232.934
R1297 VGND.n928 VGND.t325 230.54
R1298 VGND.n870 VGND.n868 214.635
R1299 VGND.n854 VGND.t139 211.857
R1300 VGND.n855 VGND.t15 211.857
R1301 VGND.n864 VGND.t78 211.857
R1302 VGND.n865 VGND.t71 211.857
R1303 VGND.n1349 VGND.t286 211.857
R1304 VGND.n1350 VGND.t192 211.857
R1305 VGND.n1347 VGND.t5 211.857
R1306 VGND.n1340 VGND.t9 211.857
R1307 VGND.t35 VGND.n876 206.97
R1308 VGND.n871 VGND.t134 206.97
R1309 VGND.t310 VGND.n870 206.97
R1310 VGND.n868 VGND.t62 206.97
R1311 VGND.n859 VGND.t291 206.97
R1312 VGND.n859 VGND.t136 206.97
R1313 VGND.t148 VGND.n858 206.97
R1314 VGND.n1408 VGND.n991 204.201
R1315 VGND.n995 VGND.n992 204.201
R1316 VGND.n1409 VGND.n990 204.201
R1317 VGND.n1432 VGND.n933 204.201
R1318 VGND.n1433 VGND.n932 204.201
R1319 VGND.n935 VGND.n934 204.201
R1320 VGND.n1383 VGND.n1382 197
R1321 VGND.n1394 VGND.n1382 197
R1322 VGND.n987 VGND.n976 197
R1323 VGND.n947 VGND.n941 197
R1324 VGND.n963 VGND.n962 197
R1325 VGND.n795 VGND.n794 197
R1326 VGND.n1711 VGND.n1647 197
R1327 VGND.n278 VGND.n222 197
R1328 VGND.n2318 VGND.n2317 197
R1329 VGND.n2263 VGND.n2262 197
R1330 VGND.n1874 VGND.n690 197
R1331 VGND.n1176 VGND.n223 197
R1332 VGND.n2212 VGND.n2211 197
R1333 VGND.n1641 VGND.n792 197
R1334 VGND.n2388 VGND.n2386 197
R1335 VGND.n1620 VGND.n805 197
R1336 VGND.n900 VGND.n899 195
R1337 VGND.n899 VGND.n851 195
R1338 VGND.n927 VGND.n926 195
R1339 VGND.n928 VGND.n927 195
R1340 VGND.n1110 VGND.t214 192.194
R1341 VGND.t214 VGND.n58 192.194
R1342 VGND.t214 VGND.n75 192.194
R1343 VGND.n1292 VGND.n1291 191.625
R1344 VGND.n1781 VGND.n787 187.249
R1345 VGND.n2338 VGND.n226 187.249
R1346 VGND.n2273 VGND.n2271 187.249
R1347 VGND.n2218 VGND.n2216 187.249
R1348 VGND.n1971 VGND.n1970 187.249
R1349 VGND.n1250 VGND.n224 187.249
R1350 VGND.n2167 VGND.n2165 187.249
R1351 VGND.n1872 VGND.n696 187.249
R1352 VGND.n2342 VGND.n2340 187.249
R1353 VGND.n905 VGND.n904 185
R1354 VGND.n894 VGND.n893 185
R1355 VGND.n1397 VGND.n1396 185
R1356 VGND.n1396 VGND.n1395 185
R1357 VGND.n1415 VGND.n974 185
R1358 VGND.n979 VGND.n974 185
R1359 VGND.n1424 VGND.n943 185
R1360 VGND.n946 VGND.n943 185
R1361 VGND.n1312 VGND.n1298 185
R1362 VGND.n1305 VGND.n1304 185
R1363 VGND.n1331 VGND.n1320 185
R1364 VGND.n1327 VGND.n1320 185
R1365 VGND.n1331 VGND.n1317 185
R1366 VGND.n1323 VGND.n1317 185
R1367 VGND.n1583 VGND.n835 185
R1368 VGND.n1598 VGND.n1597 185
R1369 VGND.n1596 VGND.n836 185
R1370 VGND.n1595 VGND.n1594 185
R1371 VGND.n1593 VGND.n1592 185
R1372 VGND.n1591 VGND.n1590 185
R1373 VGND.n1589 VGND.n1588 185
R1374 VGND.n1587 VGND.n1586 185
R1375 VGND.n1585 VGND.n1584 185
R1376 VGND.n1566 VGND.n1565 185
R1377 VGND.n1568 VGND.n1567 185
R1378 VGND.n1570 VGND.n1569 185
R1379 VGND.n1572 VGND.n1571 185
R1380 VGND.n1574 VGND.n1573 185
R1381 VGND.n1576 VGND.n1575 185
R1382 VGND.n1578 VGND.n1577 185
R1383 VGND.n1580 VGND.n1579 185
R1384 VGND.n1582 VGND.n1581 185
R1385 VGND.n1548 VGND.n1547 185
R1386 VGND.n1550 VGND.n1549 185
R1387 VGND.n1552 VGND.n1551 185
R1388 VGND.n1554 VGND.n1553 185
R1389 VGND.n1556 VGND.n1555 185
R1390 VGND.n1558 VGND.n1557 185
R1391 VGND.n1560 VGND.n1559 185
R1392 VGND.n1562 VGND.n1561 185
R1393 VGND.n1564 VGND.n1563 185
R1394 VGND.n1546 VGND.n1545 185
R1395 VGND.n1534 VGND.n1533 185
R1396 VGND.n1536 VGND.n1535 185
R1397 VGND.n1531 VGND.n820 185
R1398 VGND.n1604 VGND.n1603 185
R1399 VGND.n1601 VGND.n818 185
R1400 VGND.n1600 VGND.n814 185
R1401 VGND.n1613 VGND.n1612 185
R1402 VGND.n1615 VGND.n1614 185
R1403 VGND.n524 VGND.n523 185
R1404 VGND.n526 VGND.n481 185
R1405 VGND.n529 VGND.n528 185
R1406 VGND.n530 VGND.n480 185
R1407 VGND.n532 VGND.n531 185
R1408 VGND.n534 VGND.n479 185
R1409 VGND.n537 VGND.n536 185
R1410 VGND.n538 VGND.n478 185
R1411 VGND.n2223 VGND.n2222 185
R1412 VGND.n506 VGND.n486 185
R1413 VGND.n508 VGND.n507 185
R1414 VGND.n510 VGND.n485 185
R1415 VGND.n513 VGND.n512 185
R1416 VGND.n514 VGND.n484 185
R1417 VGND.n516 VGND.n515 185
R1418 VGND.n518 VGND.n483 185
R1419 VGND.n521 VGND.n520 185
R1420 VGND.n522 VGND.n482 185
R1421 VGND.n2257 VGND.n2256 185
R1422 VGND.n491 VGND.n466 185
R1423 VGND.n493 VGND.n492 185
R1424 VGND.n495 VGND.n489 185
R1425 VGND.n497 VGND.n496 185
R1426 VGND.n498 VGND.n488 185
R1427 VGND.n500 VGND.n499 185
R1428 VGND.n502 VGND.n487 185
R1429 VGND.n505 VGND.n504 185
R1430 VGND.n2255 VGND.n465 185
R1431 VGND.n2253 VGND.n2252 185
R1432 VGND.n469 VGND.n468 185
R1433 VGND.n2243 VGND.n2242 185
R1434 VGND.n2240 VGND.n472 185
R1435 VGND.n2238 VGND.n2237 185
R1436 VGND.n474 VGND.n473 185
R1437 VGND.n2228 VGND.n2227 185
R1438 VGND.n2225 VGND.n477 185
R1439 VGND.n1763 VGND.n1762 185
R1440 VGND.n1765 VGND.n1764 185
R1441 VGND.n1767 VGND.n1766 185
R1442 VGND.n1769 VGND.n1768 185
R1443 VGND.n1771 VGND.n1770 185
R1444 VGND.n1773 VGND.n1772 185
R1445 VGND.n1775 VGND.n1774 185
R1446 VGND.n1777 VGND.n1776 185
R1447 VGND.n1778 VGND.n778 185
R1448 VGND.n1745 VGND.n1744 185
R1449 VGND.n1747 VGND.n1746 185
R1450 VGND.n1749 VGND.n1748 185
R1451 VGND.n1751 VGND.n1750 185
R1452 VGND.n1753 VGND.n1752 185
R1453 VGND.n1755 VGND.n1754 185
R1454 VGND.n1757 VGND.n1756 185
R1455 VGND.n1759 VGND.n1758 185
R1456 VGND.n1761 VGND.n1760 185
R1457 VGND.n1727 VGND.n1726 185
R1458 VGND.n1729 VGND.n1728 185
R1459 VGND.n1731 VGND.n1730 185
R1460 VGND.n1733 VGND.n1732 185
R1461 VGND.n1735 VGND.n1734 185
R1462 VGND.n1737 VGND.n1736 185
R1463 VGND.n1739 VGND.n1738 185
R1464 VGND.n1741 VGND.n1740 185
R1465 VGND.n1743 VGND.n1742 185
R1466 VGND.n1725 VGND.n1724 185
R1467 VGND.n1715 VGND.n1714 185
R1468 VGND.n1713 VGND.n761 185
R1469 VGND.n1803 VGND.n1802 185
R1470 VGND.n760 VGND.n758 185
R1471 VGND.n1790 VGND.n1789 185
R1472 VGND.n1788 VGND.n1786 185
R1473 VGND.n781 VGND.n779 185
R1474 VGND.n1799 VGND.n1798 185
R1475 VGND.n321 VGND.n320 185
R1476 VGND.n323 VGND.n322 185
R1477 VGND.n325 VGND.n324 185
R1478 VGND.n327 VGND.n326 185
R1479 VGND.n329 VGND.n328 185
R1480 VGND.n331 VGND.n330 185
R1481 VGND.n333 VGND.n332 185
R1482 VGND.n335 VGND.n334 185
R1483 VGND.n336 VGND.n227 185
R1484 VGND.n303 VGND.n302 185
R1485 VGND.n305 VGND.n304 185
R1486 VGND.n307 VGND.n306 185
R1487 VGND.n309 VGND.n308 185
R1488 VGND.n311 VGND.n310 185
R1489 VGND.n313 VGND.n312 185
R1490 VGND.n315 VGND.n314 185
R1491 VGND.n317 VGND.n316 185
R1492 VGND.n319 VGND.n318 185
R1493 VGND.n285 VGND.n284 185
R1494 VGND.n287 VGND.n286 185
R1495 VGND.n289 VGND.n288 185
R1496 VGND.n291 VGND.n290 185
R1497 VGND.n293 VGND.n292 185
R1498 VGND.n295 VGND.n294 185
R1499 VGND.n297 VGND.n296 185
R1500 VGND.n299 VGND.n298 185
R1501 VGND.n301 VGND.n300 185
R1502 VGND.n283 VGND.n282 185
R1503 VGND.n272 VGND.n271 185
R1504 VGND.n270 VGND.n269 185
R1505 VGND.n267 VGND.n266 185
R1506 VGND.n265 VGND.n264 185
R1507 VGND.n254 VGND.n253 185
R1508 VGND.n258 VGND.n232 185
R1509 VGND.n340 VGND.n339 185
R1510 VGND.n231 VGND.n228 185
R1511 VGND.n441 VGND.n440 185
R1512 VGND.n443 VGND.n398 185
R1513 VGND.n446 VGND.n445 185
R1514 VGND.n447 VGND.n397 185
R1515 VGND.n449 VGND.n448 185
R1516 VGND.n451 VGND.n396 185
R1517 VGND.n454 VGND.n453 185
R1518 VGND.n455 VGND.n395 185
R1519 VGND.n2278 VGND.n2277 185
R1520 VGND.n423 VGND.n403 185
R1521 VGND.n425 VGND.n424 185
R1522 VGND.n427 VGND.n402 185
R1523 VGND.n430 VGND.n429 185
R1524 VGND.n431 VGND.n401 185
R1525 VGND.n433 VGND.n432 185
R1526 VGND.n435 VGND.n400 185
R1527 VGND.n438 VGND.n437 185
R1528 VGND.n439 VGND.n399 185
R1529 VGND.n2312 VGND.n2311 185
R1530 VGND.n408 VGND.n383 185
R1531 VGND.n410 VGND.n409 185
R1532 VGND.n412 VGND.n406 185
R1533 VGND.n414 VGND.n413 185
R1534 VGND.n415 VGND.n405 185
R1535 VGND.n417 VGND.n416 185
R1536 VGND.n419 VGND.n404 185
R1537 VGND.n422 VGND.n421 185
R1538 VGND.n2310 VGND.n382 185
R1539 VGND.n2308 VGND.n2307 185
R1540 VGND.n386 VGND.n385 185
R1541 VGND.n2298 VGND.n2297 185
R1542 VGND.n2295 VGND.n389 185
R1543 VGND.n2293 VGND.n2292 185
R1544 VGND.n391 VGND.n390 185
R1545 VGND.n2283 VGND.n2282 185
R1546 VGND.n2280 VGND.n394 185
R1547 VGND.n1938 VGND.n1937 185
R1548 VGND.n1940 VGND.n673 185
R1549 VGND.n1943 VGND.n1942 185
R1550 VGND.n1944 VGND.n672 185
R1551 VGND.n1946 VGND.n1945 185
R1552 VGND.n1948 VGND.n671 185
R1553 VGND.n1951 VGND.n1950 185
R1554 VGND.n1952 VGND.n670 185
R1555 VGND.n1955 VGND.n1954 185
R1556 VGND.n1920 VGND.n678 185
R1557 VGND.n1922 VGND.n1921 185
R1558 VGND.n1924 VGND.n677 185
R1559 VGND.n1927 VGND.n1926 185
R1560 VGND.n1928 VGND.n676 185
R1561 VGND.n1930 VGND.n1929 185
R1562 VGND.n1932 VGND.n675 185
R1563 VGND.n1935 VGND.n1934 185
R1564 VGND.n1936 VGND.n674 185
R1565 VGND.n1904 VGND.n1903 185
R1566 VGND.n1905 VGND.n683 185
R1567 VGND.n1907 VGND.n1906 185
R1568 VGND.n1909 VGND.n681 185
R1569 VGND.n1911 VGND.n1910 185
R1570 VGND.n1912 VGND.n680 185
R1571 VGND.n1914 VGND.n1913 185
R1572 VGND.n1916 VGND.n679 185
R1573 VGND.n1919 VGND.n1918 185
R1574 VGND.n1902 VGND.n686 185
R1575 VGND.n1900 VGND.n1899 185
R1576 VGND.n1891 VGND.n687 185
R1577 VGND.n1890 VGND.n1889 185
R1578 VGND.n1887 VGND.n1885 185
R1579 VGND.n1882 VGND.n669 185
R1580 VGND.n1963 VGND.n1962 185
R1581 VGND.n1960 VGND.n667 185
R1582 VGND.n1959 VGND.n1958 185
R1583 VGND.n1218 VGND.n1154 185
R1584 VGND.n1233 VGND.n1232 185
R1585 VGND.n1231 VGND.n1155 185
R1586 VGND.n1230 VGND.n1229 185
R1587 VGND.n1228 VGND.n1227 185
R1588 VGND.n1226 VGND.n1225 185
R1589 VGND.n1224 VGND.n1223 185
R1590 VGND.n1222 VGND.n1221 185
R1591 VGND.n1220 VGND.n1219 185
R1592 VGND.n1201 VGND.n1200 185
R1593 VGND.n1203 VGND.n1202 185
R1594 VGND.n1205 VGND.n1204 185
R1595 VGND.n1207 VGND.n1206 185
R1596 VGND.n1209 VGND.n1208 185
R1597 VGND.n1211 VGND.n1210 185
R1598 VGND.n1213 VGND.n1212 185
R1599 VGND.n1215 VGND.n1214 185
R1600 VGND.n1217 VGND.n1216 185
R1601 VGND.n1183 VGND.n1182 185
R1602 VGND.n1185 VGND.n1184 185
R1603 VGND.n1187 VGND.n1186 185
R1604 VGND.n1189 VGND.n1188 185
R1605 VGND.n1191 VGND.n1190 185
R1606 VGND.n1193 VGND.n1192 185
R1607 VGND.n1195 VGND.n1194 185
R1608 VGND.n1197 VGND.n1196 185
R1609 VGND.n1199 VGND.n1198 185
R1610 VGND.n1181 VGND.n1180 185
R1611 VGND.n1170 VGND.n1169 185
R1612 VGND.n1168 VGND.n1167 185
R1613 VGND.n1165 VGND.n1164 185
R1614 VGND.n1159 VGND.n1139 185
R1615 VGND.n1237 VGND.n1236 185
R1616 VGND.n1138 VGND.n1135 185
R1617 VGND.n1244 VGND.n1243 185
R1618 VGND.n1246 VGND.n1245 185
R1619 VGND.n636 VGND.n635 185
R1620 VGND.n638 VGND.n593 185
R1621 VGND.n641 VGND.n640 185
R1622 VGND.n642 VGND.n592 185
R1623 VGND.n644 VGND.n643 185
R1624 VGND.n646 VGND.n591 185
R1625 VGND.n649 VGND.n648 185
R1626 VGND.n650 VGND.n590 185
R1627 VGND.n2172 VGND.n2171 185
R1628 VGND.n618 VGND.n598 185
R1629 VGND.n620 VGND.n619 185
R1630 VGND.n622 VGND.n597 185
R1631 VGND.n625 VGND.n624 185
R1632 VGND.n626 VGND.n596 185
R1633 VGND.n628 VGND.n627 185
R1634 VGND.n630 VGND.n595 185
R1635 VGND.n633 VGND.n632 185
R1636 VGND.n634 VGND.n594 185
R1637 VGND.n2206 VGND.n2205 185
R1638 VGND.n603 VGND.n578 185
R1639 VGND.n605 VGND.n604 185
R1640 VGND.n607 VGND.n601 185
R1641 VGND.n609 VGND.n608 185
R1642 VGND.n610 VGND.n600 185
R1643 VGND.n612 VGND.n611 185
R1644 VGND.n614 VGND.n599 185
R1645 VGND.n617 VGND.n616 185
R1646 VGND.n2204 VGND.n577 185
R1647 VGND.n2202 VGND.n2201 185
R1648 VGND.n581 VGND.n580 185
R1649 VGND.n2192 VGND.n2191 185
R1650 VGND.n2189 VGND.n584 185
R1651 VGND.n2187 VGND.n2186 185
R1652 VGND.n586 VGND.n585 185
R1653 VGND.n2177 VGND.n2176 185
R1654 VGND.n2174 VGND.n589 185
R1655 VGND.n160 VGND.n159 185
R1656 VGND.n162 VGND.n117 185
R1657 VGND.n165 VGND.n164 185
R1658 VGND.n166 VGND.n116 185
R1659 VGND.n168 VGND.n167 185
R1660 VGND.n170 VGND.n115 185
R1661 VGND.n173 VGND.n172 185
R1662 VGND.n174 VGND.n114 185
R1663 VGND.n2347 VGND.n2346 185
R1664 VGND.n142 VGND.n122 185
R1665 VGND.n144 VGND.n143 185
R1666 VGND.n146 VGND.n121 185
R1667 VGND.n149 VGND.n148 185
R1668 VGND.n150 VGND.n120 185
R1669 VGND.n152 VGND.n151 185
R1670 VGND.n154 VGND.n119 185
R1671 VGND.n157 VGND.n156 185
R1672 VGND.n158 VGND.n118 185
R1673 VGND.n2381 VGND.n2380 185
R1674 VGND.n127 VGND.n102 185
R1675 VGND.n129 VGND.n128 185
R1676 VGND.n131 VGND.n125 185
R1677 VGND.n133 VGND.n132 185
R1678 VGND.n134 VGND.n124 185
R1679 VGND.n136 VGND.n135 185
R1680 VGND.n138 VGND.n123 185
R1681 VGND.n141 VGND.n140 185
R1682 VGND.n2379 VGND.n101 185
R1683 VGND.n2377 VGND.n2376 185
R1684 VGND.n105 VGND.n104 185
R1685 VGND.n2367 VGND.n2366 185
R1686 VGND.n2364 VGND.n108 185
R1687 VGND.n2362 VGND.n2361 185
R1688 VGND.n110 VGND.n109 185
R1689 VGND.n2352 VGND.n2351 185
R1690 VGND.n2349 VGND.n113 185
R1691 VGND.n966 VGND.n965 185
R1692 VGND.n966 VGND.n955 185
R1693 VGND.n918 VGND.n917 185
R1694 VGND.n1012 VGND.n1002 181.835
R1695 VGND.n1345 VGND.n1344 180.118
R1696 VGND.t214 VGND.n1109 175.837
R1697 VGND.t214 VGND.n59 175.837
R1698 VGND.n2424 VGND.t214 175.837
R1699 VGND.n194 VGND.n68 175.546
R1700 VGND.n194 VGND.n191 175.546
R1701 VGND.n200 VGND.n191 175.546
R1702 VGND.n200 VGND.n187 175.546
R1703 VGND.n206 VGND.n187 175.546
R1704 VGND.n208 VGND.n206 175.546
R1705 VGND.n208 VGND.n183 175.546
R1706 VGND.n214 VGND.n183 175.546
R1707 VGND.n215 VGND.n214 175.546
R1708 VGND.n215 VGND.n178 175.546
R1709 VGND.n221 VGND.n178 175.546
R1710 VGND.n1095 VGND.n1083 175.546
R1711 VGND.n1091 VGND.n1083 175.546
R1712 VGND.n1091 VGND.n1085 175.546
R1713 VGND.n1087 VGND.n1085 175.546
R1714 VGND.n1087 VGND.n62 175.546
R1715 VGND.n2450 VGND.n62 175.546
R1716 VGND.n2450 VGND.n2449 175.546
R1717 VGND.n2449 VGND.n63 175.546
R1718 VGND.n2445 VGND.n63 175.546
R1719 VGND.n2445 VGND.n65 175.546
R1720 VGND.n2441 VGND.n65 175.546
R1721 VGND.n1078 VGND.n1036 175.546
R1722 VGND.n1074 VGND.n1041 175.546
R1723 VGND.n1072 VGND.n1071 175.546
R1724 VGND.n1068 VGND.n1067 175.546
R1725 VGND.n1064 VGND.n1063 175.546
R1726 VGND.n1687 VGND.n1658 175.546
R1727 VGND.n1692 VGND.n1658 175.546
R1728 VGND.n1692 VGND.n1655 175.546
R1729 VGND.n1696 VGND.n1655 175.546
R1730 VGND.n1697 VGND.n1696 175.546
R1731 VGND.n1698 VGND.n1697 175.546
R1732 VGND.n1698 VGND.n1653 175.546
R1733 VGND.n1702 VGND.n1653 175.546
R1734 VGND.n1702 VGND.n1650 175.546
R1735 VGND.n1707 VGND.n1650 175.546
R1736 VGND.n1707 VGND.n1651 175.546
R1737 VGND.n1781 VGND.n782 175.546
R1738 VGND.n1796 VGND.n782 175.546
R1739 VGND.n1796 VGND.n783 175.546
R1740 VGND.n1792 VGND.n783 175.546
R1741 VGND.n1792 VGND.n756 175.546
R1742 VGND.n1805 VGND.n756 175.546
R1743 VGND.n1805 VGND.n757 175.546
R1744 VGND.n1717 VGND.n757 175.546
R1745 VGND.n1717 VGND.n1646 175.546
R1746 VGND.n1722 VGND.n1646 175.546
R1747 VGND.n1722 VGND.n1711 175.546
R1748 VGND.n1503 VGND.n748 175.546
R1749 VGND.n1509 VGND.n1508 175.546
R1750 VGND.n1515 VGND.n1514 175.546
R1751 VGND.n1521 VGND.n1520 175.546
R1752 VGND.n1525 VGND.n1524 175.546
R1753 VGND.n1668 VGND.n1665 175.546
R1754 VGND.n1672 VGND.n1670 175.546
R1755 VGND.n1676 VGND.n1662 175.546
R1756 VGND.n1680 VGND.n1678 175.546
R1757 VGND.n1684 VGND.n1660 175.546
R1758 VGND.n344 VGND.n342 175.546
R1759 VGND.n260 VGND.n257 175.546
R1760 VGND.n262 VGND.n256 175.546
R1761 VGND.n274 VGND.n251 175.546
R1762 VGND.n280 VGND.n276 175.546
R1763 VGND.n2047 VGND.n2034 175.546
R1764 VGND.n2043 VGND.n2034 175.546
R1765 VGND.n2043 VGND.n2036 175.546
R1766 VGND.n2039 VGND.n2036 175.546
R1767 VGND.n2039 VGND.n372 175.546
R1768 VGND.n2330 VGND.n372 175.546
R1769 VGND.n2330 VGND.n373 175.546
R1770 VGND.n2326 VGND.n373 175.546
R1771 VGND.n2326 VGND.n376 175.546
R1772 VGND.n2322 VGND.n376 175.546
R1773 VGND.n2322 VGND.n378 175.546
R1774 VGND.n2285 VGND.n393 175.546
R1775 VGND.n2289 VGND.n2287 175.546
R1776 VGND.n2300 VGND.n388 175.546
R1777 VGND.n2304 VGND.n2302 175.546
R1778 VGND.n2315 VGND.n381 175.546
R1779 VGND.n2104 VGND.n2103 175.546
R1780 VGND.n2100 VGND.n2099 175.546
R1781 VGND.n2097 VGND.n2080 175.546
R1782 VGND.n2093 VGND.n2091 175.546
R1783 VGND.n2268 VGND.n460 175.546
R1784 VGND.n2068 VGND.n2067 175.546
R1785 VGND.n2064 VGND.n2063 175.546
R1786 VGND.n2060 VGND.n2059 175.546
R1787 VGND.n2056 VGND.n2055 175.546
R1788 VGND.n2052 VGND.n2051 175.546
R1789 VGND.n2076 VGND.n2075 175.546
R1790 VGND.n2081 VGND.n2078 175.546
R1791 VGND.n2084 VGND.n2083 175.546
R1792 VGND.n2088 VGND.n2086 175.546
R1793 VGND.n2266 VGND.n462 175.546
R1794 VGND.n2230 VGND.n476 175.546
R1795 VGND.n2234 VGND.n2232 175.546
R1796 VGND.n2245 VGND.n471 175.546
R1797 VGND.n2249 VGND.n2247 175.546
R1798 VGND.n2260 VGND.n464 175.546
R1799 VGND.n548 VGND.n354 175.546
R1800 VGND.n556 VGND.n555 175.546
R1801 VGND.n560 VGND.n559 175.546
R1802 VGND.n567 VGND.n566 175.546
R1803 VGND.n570 VGND.n569 175.546
R1804 VGND.n2016 VGND.n2015 175.546
R1805 VGND.n2020 VGND.n2019 175.546
R1806 VGND.n2024 VGND.n2023 175.546
R1807 VGND.n2028 VGND.n2027 175.546
R1808 VGND.n2030 VGND.n2012 175.546
R1809 VGND.n1843 VGND.n1841 175.546
R1810 VGND.n1851 VGND.n705 175.546
R1811 VGND.n1855 VGND.n1853 175.546
R1812 VGND.n1863 VGND.n701 175.546
R1813 VGND.n1867 VGND.n1865 175.546
R1814 VGND.n718 VGND.n716 175.546
R1815 VGND.n722 VGND.n713 175.546
R1816 VGND.n726 VGND.n724 175.546
R1817 VGND.n730 VGND.n711 175.546
R1818 VGND.n734 VGND.n732 175.546
R1819 VGND.n1970 VGND.n1969 175.546
R1820 VGND.n1969 VGND.n663 175.546
R1821 VGND.n1965 VGND.n663 175.546
R1822 VGND.n1965 VGND.n666 175.546
R1823 VGND.n1883 VGND.n666 175.546
R1824 VGND.n1883 VGND.n1880 175.546
R1825 VGND.n1893 VGND.n1880 175.546
R1826 VGND.n1893 VGND.n689 175.546
R1827 VGND.n1897 VGND.n689 175.546
R1828 VGND.n1897 VGND.n1878 175.546
R1829 VGND.n1878 VGND.n690 175.546
R1830 VGND.n1988 VGND.n658 175.546
R1831 VGND.n1986 VGND.n1985 175.546
R1832 VGND.n1982 VGND.n1981 175.546
R1833 VGND.n1978 VGND.n1977 175.546
R1834 VGND.n1974 VGND.n653 175.546
R1835 VGND.n661 VGND.n653 175.546
R1836 VGND.n1052 VGND.n1043 175.546
R1837 VGND.n1045 VGND.n1044 175.546
R1838 VGND.n1047 VGND.n1046 175.546
R1839 VGND.n1049 VGND.n1048 175.546
R1840 VGND.n1051 VGND.n1050 175.546
R1841 VGND.n1248 VGND.n1131 175.546
R1842 VGND.n1241 VGND.n1239 175.546
R1843 VGND.n1162 VGND.n1160 175.546
R1844 VGND.n1172 VGND.n1158 175.546
R1845 VGND.n1178 VGND.n1174 175.546
R1846 VGND.n1277 VGND.n1020 175.546
R1847 VGND.n1273 VGND.n1020 175.546
R1848 VGND.n1273 VGND.n1123 175.546
R1849 VGND.n1269 VGND.n1123 175.546
R1850 VGND.n1269 VGND.n1125 175.546
R1851 VGND.n1265 VGND.n1125 175.546
R1852 VGND.n1265 VGND.n1127 175.546
R1853 VGND.n1261 VGND.n1127 175.546
R1854 VGND.n1261 VGND.n1129 175.546
R1855 VGND.n1257 VGND.n1129 175.546
R1856 VGND.n1257 VGND.n1254 175.546
R1857 VGND.n1119 VGND.n1019 175.546
R1858 VGND.n1119 VGND.n1022 175.546
R1859 VGND.n1115 VGND.n1022 175.546
R1860 VGND.n1115 VGND.n1025 175.546
R1861 VGND.n1111 VGND.n1025 175.546
R1862 VGND.n1111 VGND.n1027 175.546
R1863 VGND.n1107 VGND.n1027 175.546
R1864 VGND.n1107 VGND.n1030 175.546
R1865 VGND.n1103 VGND.n1030 175.546
R1866 VGND.n1103 VGND.n1032 175.546
R1867 VGND.n1099 VGND.n1032 175.546
R1868 VGND.n550 VGND.n547 175.546
R1869 VGND.n554 VGND.n552 175.546
R1870 VGND.n562 VGND.n544 175.546
R1871 VGND.n565 VGND.n564 175.546
R1872 VGND.n573 VGND.n572 175.546
R1873 VGND.n2138 VGND.n2113 175.546
R1874 VGND.n2134 VGND.n2133 175.546
R1875 VGND.n2131 VGND.n2116 175.546
R1876 VGND.n2127 VGND.n2126 175.546
R1877 VGND.n2124 VGND.n2121 175.546
R1878 VGND.n2179 VGND.n588 175.546
R1879 VGND.n2183 VGND.n2181 175.546
R1880 VGND.n2194 VGND.n583 175.546
R1881 VGND.n2198 VGND.n2196 175.546
R1882 VGND.n2209 VGND.n576 175.546
R1883 VGND.n2146 VGND.n1999 175.546
R1884 VGND.n2150 VGND.n2148 175.546
R1885 VGND.n2154 VGND.n1997 175.546
R1886 VGND.n2158 VGND.n2156 175.546
R1887 VGND.n2162 VGND.n1995 175.546
R1888 VGND.n1502 VGND.n1501 175.546
R1889 VGND.n1507 VGND.n1506 175.546
R1890 VGND.n1513 VGND.n1512 175.546
R1891 VGND.n1519 VGND.n1518 175.546
R1892 VGND.n1527 VGND.n1500 175.546
R1893 VGND.n1617 VGND.n696 175.546
R1894 VGND.n1617 VGND.n808 175.546
R1895 VGND.n1610 VGND.n808 175.546
R1896 VGND.n1610 VGND.n815 175.546
R1897 VGND.n1606 VGND.n815 175.546
R1898 VGND.n1606 VGND.n816 175.546
R1899 VGND.n1538 VGND.n816 175.546
R1900 VGND.n1538 VGND.n839 175.546
R1901 VGND.n1542 VGND.n839 175.546
R1902 VGND.n1543 VGND.n1542 175.546
R1903 VGND.n1543 VGND.n792 175.546
R1904 VGND.n1845 VGND.n707 175.546
R1905 VGND.n1849 VGND.n1847 175.546
R1906 VGND.n1857 VGND.n703 175.546
R1907 VGND.n1861 VGND.n1859 175.546
R1908 VGND.n1869 VGND.n699 175.546
R1909 VGND.n1832 VGND.n1831 175.546
R1910 VGND.n1829 VGND.n740 175.546
R1911 VGND.n1825 VGND.n1823 175.546
R1912 VGND.n1821 VGND.n742 175.546
R1913 VGND.n1817 VGND.n1815 175.546
R1914 VGND.n196 VGND.n71 175.546
R1915 VGND.n197 VGND.n196 175.546
R1916 VGND.n197 VGND.n189 175.546
R1917 VGND.n203 VGND.n189 175.546
R1918 VGND.n204 VGND.n203 175.546
R1919 VGND.n204 VGND.n185 175.546
R1920 VGND.n211 VGND.n185 175.546
R1921 VGND.n212 VGND.n211 175.546
R1922 VGND.n212 VGND.n181 175.546
R1923 VGND.n218 VGND.n181 175.546
R1924 VGND.n218 VGND.n176 175.546
R1925 VGND.n2437 VGND.n72 175.546
R1926 VGND.n2433 VGND.n72 175.546
R1927 VGND.n2433 VGND.n74 175.546
R1928 VGND.n2429 VGND.n74 175.546
R1929 VGND.n2429 VGND.n76 175.546
R1930 VGND.n2425 VGND.n76 175.546
R1931 VGND.n2425 VGND.n78 175.546
R1932 VGND.n2421 VGND.n78 175.546
R1933 VGND.n2421 VGND.n80 175.546
R1934 VGND.n2417 VGND.n80 175.546
R1935 VGND.n2417 VGND.n82 175.546
R1936 VGND.n2354 VGND.n112 175.546
R1937 VGND.n2358 VGND.n2356 175.546
R1938 VGND.n2369 VGND.n107 175.546
R1939 VGND.n2373 VGND.n2371 175.546
R1940 VGND.n2384 VGND.n100 175.546
R1941 VGND.n2412 VGND.n85 175.546
R1942 VGND.n2408 VGND.n85 175.546
R1943 VGND.n2408 VGND.n87 175.546
R1944 VGND.n2404 VGND.n87 175.546
R1945 VGND.n2404 VGND.n90 175.546
R1946 VGND.n2400 VGND.n90 175.546
R1947 VGND.n2400 VGND.n92 175.546
R1948 VGND.n2396 VGND.n92 175.546
R1949 VGND.n2396 VGND.n94 175.546
R1950 VGND.n2392 VGND.n94 175.546
R1951 VGND.n2392 VGND.n96 175.546
R1952 VGND.n1466 VGND.t186 175.221
R1953 VGND.t68 VGND.n1490 175.221
R1954 VGND.n1058 VGND.t214 172.876
R1955 VGND.n1080 VGND.t214 172.615
R1956 VGND.n1493 VGND.n844 171.327
R1957 VGND.n841 VGND.t214 170.321
R1958 VGND.n977 VGND.t27 169.615
R1959 VGND.t143 VGND.t310 168.642
R1960 VGND.t70 VGND.t62 168.642
R1961 VGND.t291 VGND.t77 168.642
R1962 VGND.t136 VGND.t14 168.642
R1963 VGND.t138 VGND.t148 168.642
R1964 VGND.t144 VGND.n1345 167.251
R1965 VGND.n979 VGND.n978 166.63
R1966 VGND.n946 VGND.n945 166.63
R1967 VGND.n939 VGND.t239 164.626
R1968 VGND.n1028 VGND.n1024 163.57
R1969 VGND.n1547 VGND.n1546 163.333
R1970 VGND.n2256 VGND.n2255 163.333
R1971 VGND.n1726 VGND.n1725 163.333
R1972 VGND.n284 VGND.n283 163.333
R1973 VGND.n2311 VGND.n2310 163.333
R1974 VGND.n1903 VGND.n1902 163.333
R1975 VGND.n1182 VGND.n1181 163.333
R1976 VGND.n2205 VGND.n2204 163.333
R1977 VGND.n2380 VGND.n2379 163.333
R1978 VGND.n1023 VGND.t214 159.421
R1979 VGND.n2454 VGND.n57 157.601
R1980 VGND.n1369 VGND.t204 155.611
R1981 VGND.n911 VGND.n910 153.601
R1982 VGND.n1579 VGND.n1578 150
R1983 VGND.n1575 VGND.n1574 150
R1984 VGND.n1571 VGND.n1570 150
R1985 VGND.n1567 VGND.n1566 150
R1986 VGND.n1563 VGND.n1562 150
R1987 VGND.n1559 VGND.n1558 150
R1988 VGND.n1555 VGND.n1554 150
R1989 VGND.n1551 VGND.n1550 150
R1990 VGND.n1614 VGND.n1613 150
R1991 VGND.n1601 VGND.n1600 150
R1992 VGND.n1603 VGND.n820 150
R1993 VGND.n1535 VGND.n1534 150
R1994 VGND.n1598 VGND.n836 150
R1995 VGND.n1594 VGND.n1593 150
R1996 VGND.n1590 VGND.n1589 150
R1997 VGND.n1586 VGND.n1585 150
R1998 VGND.n520 VGND.n518 150
R1999 VGND.n516 VGND.n484 150
R2000 VGND.n512 VGND.n510 150
R2001 VGND.n508 VGND.n486 150
R2002 VGND.n504 VGND.n502 150
R2003 VGND.n500 VGND.n488 150
R2004 VGND.n496 VGND.n495 150
R2005 VGND.n493 VGND.n491 150
R2006 VGND.n2227 VGND.n2225 150
R2007 VGND.n2238 VGND.n473 150
R2008 VGND.n2242 VGND.n2240 150
R2009 VGND.n2253 VGND.n468 150
R2010 VGND.n528 VGND.n526 150
R2011 VGND.n532 VGND.n480 150
R2012 VGND.n536 VGND.n534 150
R2013 VGND.n2223 VGND.n478 150
R2014 VGND.n1758 VGND.n1757 150
R2015 VGND.n1754 VGND.n1753 150
R2016 VGND.n1750 VGND.n1749 150
R2017 VGND.n1746 VGND.n1745 150
R2018 VGND.n1742 VGND.n1741 150
R2019 VGND.n1738 VGND.n1737 150
R2020 VGND.n1734 VGND.n1733 150
R2021 VGND.n1730 VGND.n1729 150
R2022 VGND.n1799 VGND.n779 150
R2023 VGND.n1789 VGND.n1788 150
R2024 VGND.n1802 VGND.n760 150
R2025 VGND.n1714 VGND.n761 150
R2026 VGND.n1766 VGND.n1765 150
R2027 VGND.n1770 VGND.n1769 150
R2028 VGND.n1774 VGND.n1773 150
R2029 VGND.n1776 VGND.n778 150
R2030 VGND.n316 VGND.n315 150
R2031 VGND.n312 VGND.n311 150
R2032 VGND.n308 VGND.n307 150
R2033 VGND.n304 VGND.n303 150
R2034 VGND.n300 VGND.n299 150
R2035 VGND.n296 VGND.n295 150
R2036 VGND.n292 VGND.n291 150
R2037 VGND.n288 VGND.n287 150
R2038 VGND.n339 VGND.n231 150
R2039 VGND.n253 VGND.n232 150
R2040 VGND.n266 VGND.n265 150
R2041 VGND.n271 VGND.n270 150
R2042 VGND.n324 VGND.n323 150
R2043 VGND.n328 VGND.n327 150
R2044 VGND.n332 VGND.n331 150
R2045 VGND.n336 VGND.n335 150
R2046 VGND.n437 VGND.n435 150
R2047 VGND.n433 VGND.n401 150
R2048 VGND.n429 VGND.n427 150
R2049 VGND.n425 VGND.n403 150
R2050 VGND.n421 VGND.n419 150
R2051 VGND.n417 VGND.n405 150
R2052 VGND.n413 VGND.n412 150
R2053 VGND.n410 VGND.n408 150
R2054 VGND.n2282 VGND.n2280 150
R2055 VGND.n2293 VGND.n390 150
R2056 VGND.n2297 VGND.n2295 150
R2057 VGND.n2308 VGND.n385 150
R2058 VGND.n445 VGND.n443 150
R2059 VGND.n449 VGND.n397 150
R2060 VGND.n453 VGND.n451 150
R2061 VGND.n2278 VGND.n395 150
R2062 VGND.n1934 VGND.n1932 150
R2063 VGND.n1930 VGND.n676 150
R2064 VGND.n1926 VGND.n1924 150
R2065 VGND.n1922 VGND.n678 150
R2066 VGND.n1918 VGND.n1916 150
R2067 VGND.n1914 VGND.n680 150
R2068 VGND.n1910 VGND.n1909 150
R2069 VGND.n1907 VGND.n683 150
R2070 VGND.n1960 VGND.n1959 150
R2071 VGND.n1962 VGND.n669 150
R2072 VGND.n1889 VGND.n1887 150
R2073 VGND.n1900 VGND.n687 150
R2074 VGND.n1942 VGND.n1940 150
R2075 VGND.n1946 VGND.n672 150
R2076 VGND.n1950 VGND.n1948 150
R2077 VGND.n1955 VGND.n670 150
R2078 VGND.n1214 VGND.n1213 150
R2079 VGND.n1210 VGND.n1209 150
R2080 VGND.n1206 VGND.n1205 150
R2081 VGND.n1202 VGND.n1201 150
R2082 VGND.n1198 VGND.n1197 150
R2083 VGND.n1194 VGND.n1193 150
R2084 VGND.n1190 VGND.n1189 150
R2085 VGND.n1186 VGND.n1185 150
R2086 VGND.n1245 VGND.n1244 150
R2087 VGND.n1236 VGND.n1138 150
R2088 VGND.n1164 VGND.n1139 150
R2089 VGND.n1169 VGND.n1168 150
R2090 VGND.n1233 VGND.n1155 150
R2091 VGND.n1229 VGND.n1228 150
R2092 VGND.n1225 VGND.n1224 150
R2093 VGND.n1221 VGND.n1220 150
R2094 VGND.n632 VGND.n630 150
R2095 VGND.n628 VGND.n596 150
R2096 VGND.n624 VGND.n622 150
R2097 VGND.n620 VGND.n598 150
R2098 VGND.n616 VGND.n614 150
R2099 VGND.n612 VGND.n600 150
R2100 VGND.n608 VGND.n607 150
R2101 VGND.n605 VGND.n603 150
R2102 VGND.n2176 VGND.n2174 150
R2103 VGND.n2187 VGND.n585 150
R2104 VGND.n2191 VGND.n2189 150
R2105 VGND.n2202 VGND.n580 150
R2106 VGND.n640 VGND.n638 150
R2107 VGND.n644 VGND.n592 150
R2108 VGND.n648 VGND.n646 150
R2109 VGND.n2172 VGND.n590 150
R2110 VGND.n156 VGND.n154 150
R2111 VGND.n152 VGND.n120 150
R2112 VGND.n148 VGND.n146 150
R2113 VGND.n144 VGND.n122 150
R2114 VGND.n140 VGND.n138 150
R2115 VGND.n136 VGND.n124 150
R2116 VGND.n132 VGND.n131 150
R2117 VGND.n129 VGND.n127 150
R2118 VGND.n2351 VGND.n2349 150
R2119 VGND.n2362 VGND.n109 150
R2120 VGND.n2366 VGND.n2364 150
R2121 VGND.n2377 VGND.n104 150
R2122 VGND.n164 VGND.n162 150
R2123 VGND.n168 VGND.n116 150
R2124 VGND.n172 VGND.n170 150
R2125 VGND.n2347 VGND.n114 150
R2126 VGND.n1008 VGND.n1004 147.716
R2127 VGND.n1009 VGND.n1005 147.716
R2128 VGND.n1640 VGND.n1639 146.041
R2129 VGND.n33 VGND.n32 145.243
R2130 VGND.n36 VGND.n35 145.243
R2131 VGND.n925 VGND.n889 144
R2132 VGND.t0 VGND.t270 142.774
R2133 VGND.t141 VGND.t0 142.774
R2134 VGND.t72 VGND.t206 142.774
R2135 VGND.t56 VGND.t72 142.774
R2136 VGND.t200 VGND.t56 142.774
R2137 VGND.t79 VGND.t106 142.774
R2138 VGND.t140 VGND.t79 142.774
R2139 VGND.t272 VGND.t202 142.774
R2140 VGND.t289 VGND.t272 142.774
R2141 VGND.t23 VGND.t289 142.774
R2142 VGND.t111 VGND.t54 142.774
R2143 VGND.t54 VGND.t43 142.774
R2144 VGND.t98 VGND.t92 142.774
R2145 VGND.t92 VGND.t122 142.774
R2146 VGND.t122 VGND.t173 142.774
R2147 VGND.t188 VGND.t171 142.774
R2148 VGND.t119 VGND.t188 142.774
R2149 VGND.t49 VGND.t162 142.774
R2150 VGND.t12 VGND.t49 142.774
R2151 VGND.t58 VGND.t12 142.774
R2152 VGND.t322 VGND.t118 142.774
R2153 VGND.t186 VGND.t322 142.774
R2154 VGND.t164 VGND.t2 142.774
R2155 VGND.t2 VGND.t51 142.774
R2156 VGND.t51 VGND.t104 142.774
R2157 VGND.t95 VGND.t68 142.774
R2158 VGND.t120 VGND.t130 142.774
R2159 VGND.t20 VGND.t120 142.774
R2160 VGND.t318 VGND.t20 142.774
R2161 VGND.t127 VGND.t150 142.774
R2162 VGND.t64 VGND.t127 142.774
R2163 VGND.t83 VGND.t64 142.774
R2164 VGND.t151 VGND.t60 142.774
R2165 VGND.t303 VGND.t151 142.774
R2166 VGND.t294 VGND.t303 142.774
R2167 VGND.t307 VGND.t146 142.774
R2168 VGND.t29 VGND.t314 142.774
R2169 VGND.t113 VGND.t29 142.774
R2170 VGND.t168 VGND.t113 142.774
R2171 VGND.n1290 VGND.n1284 142.246
R2172 VGND.n1288 VGND.n1287 142.246
R2173 VGND.n806 VGND.n695 138.81
R2174 VGND.t96 VGND.t110 136.749
R2175 VGND.t208 VGND.n1875 135.919
R2176 VGND.n924 VGND.t326 134.954
R2177 VGND.t125 VGND.t248 134.695
R2178 VGND.n908 VGND.t48 134.62
R2179 VGND.n897 VGND.t197 134.62
R2180 VGND.n921 VGND.t11 134.62
R2181 VGND.n1402 VGND.t234 134.501
R2182 VGND.n1429 VGND.t265 134.501
R2183 VGND.n786 VGND.t324 134.474
R2184 VGND.n1320 VGND.n1319 134.268
R2185 VGND.n1319 VGND.n1317 134.268
R2186 VGND.n844 VGND.n843 133.04
R2187 VGND.n2164 VGND.n2163 132.721
R2188 VGND.n911 VGND.n898 131.201
R2189 VGND.n1352 VGND.t317 130.713
R2190 VGND.n1967 VGND.n1966 130.136
R2191 VGND.n1894 VGND.n1879 130.136
R2192 VGND.n1877 VGND.n1876 130.136
R2193 VGND.n1618 VGND.n807 130.136
R2194 VGND.n1609 VGND.n807 130.136
R2195 VGND.n1609 VGND.n1608 130.136
R2196 VGND.n1608 VGND.n1607 130.136
R2197 VGND.n1539 VGND.n1530 130.136
R2198 VGND.n1540 VGND.n1539 130.136
R2199 VGND.n1541 VGND.n1540 130.136
R2200 VGND.n1541 VGND.n793 130.136
R2201 VGND.n1783 VGND.n1782 130.136
R2202 VGND.n1793 VGND.n1784 130.136
R2203 VGND.n1719 VGND.n1718 130.136
R2204 VGND.n857 VGND.t149 130.001
R2205 VGND.n867 VGND.t63 130.001
R2206 VGND.n869 VGND.t311 130.001
R2207 VGND.n872 VGND.t135 130.001
R2208 VGND.n875 VGND.t36 130.001
R2209 VGND.n1359 VGND.t133 130.001
R2210 VGND.n1361 VGND.t116 130.001
R2211 VGND.n1343 VGND.t145 130.001
R2212 VGND.n1356 VGND.t86 130.001
R2213 VGND.n862 VGND.t292 130.001
R2214 VGND.n860 VGND.t137 130.001
R2215 VGND.n1346 VGND.t321 130.001
R2216 VGND.n1364 VGND.t89 130
R2217 VGND.t158 VGND.t236 129.706
R2218 VGND.t66 VGND.t128 129.706
R2219 VGND.t39 VGND.t267 129.706
R2220 VGND.t308 VGND.t220 129.706
R2221 VGND.n1720 VGND.t280 127.468
R2222 VGND.n2488 VGND.n2487 127.031
R2223 VGND.n2492 VGND.n2491 127.031
R2224 VGND.n20 VGND.n19 127.031
R2225 VGND.n24 VGND.n23 127.031
R2226 VGND.t218 VGND.n695 125.797
R2227 VGND.n1794 VGND.t195 125.797
R2228 VGND.t142 VGND.n1712 125.797
R2229 VGND.n222 VGND.n221 124.832
R2230 VGND.n2338 VGND.n225 124.832
R2231 VGND.n789 VGND.n787 124.832
R2232 VGND.n2271 VGND.n2270 124.832
R2233 VGND.n2264 VGND.n2263 124.832
R2234 VGND.n2216 VGND.n2215 124.832
R2235 VGND.n1874 VGND.n692 124.832
R2236 VGND.n1060 VGND.n223 124.832
R2237 VGND.n2213 VGND.n2212 124.832
R2238 VGND.n1641 VGND.n791 124.832
R2239 VGND.n1872 VGND.n1871 124.832
R2240 VGND.n2340 VGND.n176 124.832
R2241 VGND.t276 VGND.t160 124.718
R2242 VGND.t251 VGND.t22 124.718
R2243 VGND.n1640 VGND.t218 124.352
R2244 VGND.n877 VGND.t26 122.501
R2245 VGND.n880 VGND.t76 122.501
R2246 VGND.n882 VGND.t297 122.501
R2247 VGND.n1367 VGND.t205 122.501
R2248 VGND.n1371 VGND.t97 122.501
R2249 VGND.n1373 VGND.t91 122.501
R2250 VGND.n665 VGND.t81 120.013
R2251 VGND.n1895 VGND.t124 120.013
R2252 VGND.t7 VGND.t305 114.74
R2253 VGND.t41 VGND.t102 114.74
R2254 VGND.n1341 VGND.t132 113.945
R2255 VGND.n1337 VGND.t218 111.68
R2256 VGND.n1427 VGND.t224 109.751
R2257 VGND.t244 VGND.t264 109.751
R2258 VGND.n1292 VGND.n1282 108.8
R2259 VGND.n1012 VGND.n1011 108.047
R2260 VGND.n1374 VGND.t110 106.099
R2261 VGND.n1370 VGND.t278 106.099
R2262 VGND.n1381 VGND.n1380 103.734
R2263 VGND.n1406 VGND.n1405 102.136
R2264 VGND.n1001 VGND.n1000 102.136
R2265 VGND.n999 VGND.n998 102.136
R2266 VGND.n997 VGND.n996 102.136
R2267 VGND.n1428 VGND.n936 102.136
R2268 VGND.n1303 VGND.n1302 101.718
R2269 VGND.n1322 VGND.n1321 101.718
R2270 VGND.n1330 VGND.n1329 101.718
R2271 VGND.n1311 VGND.n1310 101.718
R2272 VGND.n1427 VGND.n1426 99.7737
R2273 VGND.t255 VGND.n1412 99.7737
R2274 VGND.t218 VGND.n363 47.6748
R2275 VGND.n1968 VGND.t293 96.8786
R2276 VGND.n99 VGND.n97 95.7473
R2277 VGND.t193 VGND.t276 94.7851
R2278 VGND.n1426 VGND.t170 94.7851
R2279 VGND.n2112 VGND.n97 92.4832
R2280 VGND.n984 VGND.n974 91.3721
R2281 VGND.n981 VGND.n975 91.3721
R2282 VGND.n982 VGND.n981 91.3721
R2283 VGND.n948 VGND.n943 91.3721
R2284 VGND.n1423 VGND.n1422 91.3721
R2285 VGND.n1422 VGND.n952 91.3721
R2286 VGND.n1721 VGND.t274 91.0948
R2287 VGND.n1308 VGND.n1298 91.069
R2288 VGND.n1301 VGND.n1298 91.069
R2289 VGND.n1305 VGND.n1297 91.069
R2290 VGND.n1306 VGND.n1305 91.069
R2291 VGND.n1324 VGND.n1320 91.069
R2292 VGND.n1326 VGND.n1317 91.069
R2293 VGND.n1396 VGND.n1390 90.7567
R2294 VGND.n966 VGND.n954 90.7567
R2295 VGND.n1437 VGND.n930 89.7964
R2296 VGND.n906 VGND.n905 87.4584
R2297 VGND.n895 VGND.n894 87.4584
R2298 VGND.n919 VGND.n918 87.4584
R2299 VGND.t211 VGND.t16 86.757
R2300 VGND.t190 VGND.t196 86.757
R2301 VGND.n2112 VGND.t218 84.867
R2302 VGND.t128 VGND.t228 84.8078
R2303 VGND.n1637 VGND.n795 84.306
R2304 VGND.n1622 VGND.n805 84.306
R2305 VGND.n964 VGND.n963 84.306
R2306 VGND.n962 VGND.n961 84.306
R2307 VGND.n1425 VGND.n941 84.306
R2308 VGND.n947 VGND.n940 84.306
R2309 VGND.n1414 VGND.n976 84.306
R2310 VGND.n988 VGND.n987 84.306
R2311 VGND.n1398 VGND.n1383 84.306
R2312 VGND.n1408 VGND.n995 83.2005
R2313 VGND.n1409 VGND.n1408 83.2005
R2314 VGND.n1621 VGND.n806 82.4192
R2315 VGND.n1795 VGND.t117 82.4192
R2316 VGND.n1806 VGND.t177 82.4192
R2317 VGND.n1721 VGND.t74 82.4192
R2318 VGND.n2439 VGND.n69 80.9821
R2319 VGND.n1370 VGND.t96 77.8057
R2320 VGND.t204 VGND.n1368 77.8057
R2321 VGND.n1968 VGND.t209 76.6354
R2322 VGND.t210 VGND.n366 76.6354
R2323 VGND.n1896 VGND.t87 76.6354
R2324 VGND.n1639 VGND.n1638 76.6354
R2325 VGND.n1082 VGND.n1081 76.3222
R2326 VGND.n1079 VGND.n1078 76.3222
R2327 VGND.n1074 VGND.n1040 76.3222
R2328 VGND.n1071 VGND.n1039 76.3222
R2329 VGND.n1067 VGND.n1038 76.3222
R2330 VGND.n1063 VGND.n1037 76.3222
R2331 VGND.n1809 VGND.n1808 76.3222
R2332 VGND.n1503 VGND.n753 76.3222
R2333 VGND.n1509 VGND.n752 76.3222
R2334 VGND.n1515 VGND.n751 76.3222
R2335 VGND.n1521 VGND.n750 76.3222
R2336 VGND.n1525 VGND.n749 76.3222
R2337 VGND.n1665 VGND.n1664 76.3222
R2338 VGND.n1670 VGND.n1669 76.3222
R2339 VGND.n1671 VGND.n1662 76.3222
R2340 VGND.n1678 VGND.n1677 76.3222
R2341 VGND.n1679 VGND.n1660 76.3222
R2342 VGND.n1686 VGND.n1685 76.3222
R2343 VGND.n343 VGND.n226 76.3222
R2344 VGND.n342 VGND.n229 76.3222
R2345 VGND.n261 VGND.n260 76.3222
R2346 VGND.n256 VGND.n255 76.3222
R2347 VGND.n275 VGND.n274 76.3222
R2348 VGND.n280 VGND.n279 76.3222
R2349 VGND.n2273 VGND.n2272 76.3222
R2350 VGND.n2286 VGND.n2285 76.3222
R2351 VGND.n2289 VGND.n2288 76.3222
R2352 VGND.n2301 VGND.n2300 76.3222
R2353 VGND.n2304 VGND.n2303 76.3222
R2354 VGND.n2316 VGND.n2315 76.3222
R2355 VGND.n2106 VGND.n2105 76.3222
R2356 VGND.n2103 VGND.n2073 76.3222
R2357 VGND.n2099 VGND.n2098 76.3222
R2358 VGND.n2092 VGND.n2080 76.3222
R2359 VGND.n2091 VGND.n2090 76.3222
R2360 VGND.n2269 VGND.n2268 76.3222
R2361 VGND.n2068 VGND.n2001 76.3222
R2362 VGND.n2064 VGND.n2002 76.3222
R2363 VGND.n2060 VGND.n2003 76.3222
R2364 VGND.n2056 VGND.n2004 76.3222
R2365 VGND.n2052 VGND.n2005 76.3222
R2366 VGND.n2048 VGND.n2006 76.3222
R2367 VGND.n2075 VGND.n2074 76.3222
R2368 VGND.n2078 VGND.n2077 76.3222
R2369 VGND.n2083 VGND.n2082 76.3222
R2370 VGND.n2086 VGND.n2085 76.3222
R2371 VGND.n2087 VGND.n462 76.3222
R2372 VGND.n2265 VGND.n2264 76.3222
R2373 VGND.n2218 VGND.n2217 76.3222
R2374 VGND.n2231 VGND.n2230 76.3222
R2375 VGND.n2234 VGND.n2233 76.3222
R2376 VGND.n2246 VGND.n2245 76.3222
R2377 VGND.n2249 VGND.n2248 76.3222
R2378 VGND.n2261 VGND.n2260 76.3222
R2379 VGND.n2334 VGND.n2333 76.3222
R2380 VGND.n548 VGND.n359 76.3222
R2381 VGND.n556 VGND.n358 76.3222
R2382 VGND.n560 VGND.n357 76.3222
R2383 VGND.n567 VGND.n356 76.3222
R2384 VGND.n569 VGND.n355 76.3222
R2385 VGND.n2015 VGND.n2007 76.3222
R2386 VGND.n2019 VGND.n2008 76.3222
R2387 VGND.n2023 VGND.n2009 76.3222
R2388 VGND.n2027 VGND.n2010 76.3222
R2389 VGND.n2030 VGND.n2011 76.3222
R2390 VGND.n2111 VGND.n2110 76.3222
R2391 VGND.n1840 VGND.n1839 76.3222
R2392 VGND.n1843 VGND.n1842 76.3222
R2393 VGND.n1852 VGND.n1851 76.3222
R2394 VGND.n1855 VGND.n1854 76.3222
R2395 VGND.n1864 VGND.n1863 76.3222
R2396 VGND.n1867 VGND.n1866 76.3222
R2397 VGND.n715 VGND.n659 76.3222
R2398 VGND.n718 VGND.n717 76.3222
R2399 VGND.n723 VGND.n722 76.3222
R2400 VGND.n726 VGND.n725 76.3222
R2401 VGND.n731 VGND.n730 76.3222
R2402 VGND.n734 VGND.n733 76.3222
R2403 VGND.n1993 VGND.n1992 76.3222
R2404 VGND.n1988 VGND.n657 76.3222
R2405 VGND.n1985 VGND.n656 76.3222
R2406 VGND.n1981 VGND.n655 76.3222
R2407 VGND.n1977 VGND.n654 76.3222
R2408 VGND.n1053 VGND.n1052 76.3222
R2409 VGND.n1054 VGND.n1044 76.3222
R2410 VGND.n1055 VGND.n1046 76.3222
R2411 VGND.n1056 VGND.n1048 76.3222
R2412 VGND.n1057 VGND.n1050 76.3222
R2413 VGND.n1060 VGND.n1059 76.3222
R2414 VGND.n1250 VGND.n1249 76.3222
R2415 VGND.n1240 VGND.n1131 76.3222
R2416 VGND.n1239 VGND.n1136 76.3222
R2417 VGND.n1162 VGND.n1161 76.3222
R2418 VGND.n1173 VGND.n1172 76.3222
R2419 VGND.n1178 VGND.n1177 76.3222
R2420 VGND.n1993 VGND.n658 76.3222
R2421 VGND.n1986 VGND.n657 76.3222
R2422 VGND.n1982 VGND.n656 76.3222
R2423 VGND.n1978 VGND.n655 76.3222
R2424 VGND.n1974 VGND.n654 76.3222
R2425 VGND.n547 VGND.n546 76.3222
R2426 VGND.n552 VGND.n551 76.3222
R2427 VGND.n553 VGND.n544 76.3222
R2428 VGND.n564 VGND.n563 76.3222
R2429 VGND.n572 VGND.n542 76.3222
R2430 VGND.n2213 VGND.n574 76.3222
R2431 VGND.n2139 VGND.n2138 76.3222
R2432 VGND.n2134 VGND.n2115 76.3222
R2433 VGND.n2132 VGND.n2131 76.3222
R2434 VGND.n2127 VGND.n2118 76.3222
R2435 VGND.n2125 VGND.n2124 76.3222
R2436 VGND.n2120 VGND.n2119 76.3222
R2437 VGND.n2167 VGND.n2166 76.3222
R2438 VGND.n2180 VGND.n2179 76.3222
R2439 VGND.n2183 VGND.n2182 76.3222
R2440 VGND.n2195 VGND.n2194 76.3222
R2441 VGND.n2198 VGND.n2197 76.3222
R2442 VGND.n2210 VGND.n2209 76.3222
R2443 VGND.n2142 VGND.n2141 76.3222
R2444 VGND.n2147 VGND.n2146 76.3222
R2445 VGND.n2150 VGND.n2149 76.3222
R2446 VGND.n2155 VGND.n2154 76.3222
R2447 VGND.n2158 VGND.n2157 76.3222
R2448 VGND.n2163 VGND.n2162 76.3222
R2449 VGND.n2141 VGND.n1999 76.3222
R2450 VGND.n2148 VGND.n2147 76.3222
R2451 VGND.n2149 VGND.n1997 76.3222
R2452 VGND.n2156 VGND.n2155 76.3222
R2453 VGND.n2157 VGND.n1995 76.3222
R2454 VGND.n2121 VGND.n2120 76.3222
R2455 VGND.n2126 VGND.n2125 76.3222
R2456 VGND.n2118 VGND.n2116 76.3222
R2457 VGND.n2133 VGND.n2132 76.3222
R2458 VGND.n2115 VGND.n2113 76.3222
R2459 VGND.n2140 VGND.n2139 76.3222
R2460 VGND.n2111 VGND.n2012 76.3222
R2461 VGND.n2028 VGND.n2011 76.3222
R2462 VGND.n2024 VGND.n2010 76.3222
R2463 VGND.n2020 VGND.n2009 76.3222
R2464 VGND.n2016 VGND.n2008 76.3222
R2465 VGND.n2007 VGND.n353 76.3222
R2466 VGND.n2051 VGND.n2006 76.3222
R2467 VGND.n2055 VGND.n2005 76.3222
R2468 VGND.n2059 VGND.n2004 76.3222
R2469 VGND.n2063 VGND.n2003 76.3222
R2470 VGND.n2067 VGND.n2002 76.3222
R2471 VGND.n2072 VGND.n2001 76.3222
R2472 VGND.n1249 VGND.n1248 76.3222
R2473 VGND.n1241 VGND.n1240 76.3222
R2474 VGND.n1160 VGND.n1136 76.3222
R2475 VGND.n1161 VGND.n1158 76.3222
R2476 VGND.n1174 VGND.n1173 76.3222
R2477 VGND.n1177 VGND.n1176 76.3222
R2478 VGND.n344 VGND.n343 76.3222
R2479 VGND.n257 VGND.n229 76.3222
R2480 VGND.n262 VGND.n261 76.3222
R2481 VGND.n255 VGND.n251 76.3222
R2482 VGND.n276 VGND.n275 76.3222
R2483 VGND.n279 VGND.n278 76.3222
R2484 VGND.n1685 VGND.n1684 76.3222
R2485 VGND.n1680 VGND.n1679 76.3222
R2486 VGND.n1677 VGND.n1676 76.3222
R2487 VGND.n1672 VGND.n1671 76.3222
R2488 VGND.n1669 VGND.n1668 76.3222
R2489 VGND.n1664 VGND.n747 76.3222
R2490 VGND.n2166 VGND.n588 76.3222
R2491 VGND.n2181 VGND.n2180 76.3222
R2492 VGND.n2182 VGND.n583 76.3222
R2493 VGND.n2196 VGND.n2195 76.3222
R2494 VGND.n2197 VGND.n576 76.3222
R2495 VGND.n2211 VGND.n2210 76.3222
R2496 VGND.n2217 VGND.n476 76.3222
R2497 VGND.n2232 VGND.n2231 76.3222
R2498 VGND.n2233 VGND.n471 76.3222
R2499 VGND.n2247 VGND.n2246 76.3222
R2500 VGND.n2248 VGND.n464 76.3222
R2501 VGND.n2262 VGND.n2261 76.3222
R2502 VGND.n2272 VGND.n393 76.3222
R2503 VGND.n2287 VGND.n2286 76.3222
R2504 VGND.n2288 VGND.n388 76.3222
R2505 VGND.n2302 VGND.n2301 76.3222
R2506 VGND.n2303 VGND.n381 76.3222
R2507 VGND.n2317 VGND.n2316 76.3222
R2508 VGND.n1501 VGND.n1495 76.3222
R2509 VGND.n1506 VGND.n1496 76.3222
R2510 VGND.n1512 VGND.n1497 76.3222
R2511 VGND.n1518 VGND.n1498 76.3222
R2512 VGND.n1500 VGND.n1499 76.3222
R2513 VGND.n1528 VGND.n791 76.3222
R2514 VGND.n1837 VGND.n1836 76.3222
R2515 VGND.n1846 VGND.n1845 76.3222
R2516 VGND.n1849 VGND.n1848 76.3222
R2517 VGND.n1858 VGND.n1857 76.3222
R2518 VGND.n1861 VGND.n1860 76.3222
R2519 VGND.n1870 VGND.n1869 76.3222
R2520 VGND.n1835 VGND.n738 76.3222
R2521 VGND.n1831 VGND.n1830 76.3222
R2522 VGND.n1824 VGND.n740 76.3222
R2523 VGND.n1823 VGND.n1822 76.3222
R2524 VGND.n1816 VGND.n742 76.3222
R2525 VGND.n1815 VGND.n1814 76.3222
R2526 VGND.n1814 VGND.n1813 76.3222
R2527 VGND.n1817 VGND.n1816 76.3222
R2528 VGND.n1822 VGND.n1821 76.3222
R2529 VGND.n1825 VGND.n1824 76.3222
R2530 VGND.n1830 VGND.n1829 76.3222
R2531 VGND.n1832 VGND.n738 76.3222
R2532 VGND.n733 VGND.n709 76.3222
R2533 VGND.n732 VGND.n731 76.3222
R2534 VGND.n725 VGND.n711 76.3222
R2535 VGND.n724 VGND.n723 76.3222
R2536 VGND.n717 VGND.n713 76.3222
R2537 VGND.n716 VGND.n715 76.3222
R2538 VGND.n1866 VGND.n692 76.3222
R2539 VGND.n1865 VGND.n1864 76.3222
R2540 VGND.n1854 VGND.n701 76.3222
R2541 VGND.n1853 VGND.n1852 76.3222
R2542 VGND.n1842 VGND.n705 76.3222
R2543 VGND.n1841 VGND.n1840 76.3222
R2544 VGND.n1836 VGND.n707 76.3222
R2545 VGND.n1847 VGND.n1846 76.3222
R2546 VGND.n1848 VGND.n703 76.3222
R2547 VGND.n1859 VGND.n1858 76.3222
R2548 VGND.n1860 VGND.n699 76.3222
R2549 VGND.n1871 VGND.n1870 76.3222
R2550 VGND.n574 VGND.n573 76.3222
R2551 VGND.n565 VGND.n542 76.3222
R2552 VGND.n563 VGND.n562 76.3222
R2553 VGND.n554 VGND.n553 76.3222
R2554 VGND.n551 VGND.n550 76.3222
R2555 VGND.n546 VGND.n351 76.3222
R2556 VGND.n2333 VGND.n354 76.3222
R2557 VGND.n555 VGND.n359 76.3222
R2558 VGND.n559 VGND.n358 76.3222
R2559 VGND.n566 VGND.n357 76.3222
R2560 VGND.n570 VGND.n356 76.3222
R2561 VGND.n2215 VGND.n355 76.3222
R2562 VGND.n1059 VGND.n1051 76.3222
R2563 VGND.n1057 VGND.n1049 76.3222
R2564 VGND.n1056 VGND.n1047 76.3222
R2565 VGND.n1055 VGND.n1045 76.3222
R2566 VGND.n1054 VGND.n1043 76.3222
R2567 VGND.n1053 VGND.n1033 76.3222
R2568 VGND.n1081 VGND.n1036 76.3222
R2569 VGND.n1079 VGND.n1041 76.3222
R2570 VGND.n1072 VGND.n1040 76.3222
R2571 VGND.n1068 VGND.n1039 76.3222
R2572 VGND.n1064 VGND.n1038 76.3222
R2573 VGND.n1037 VGND.n225 76.3222
R2574 VGND.n2342 VGND.n2341 76.3222
R2575 VGND.n2355 VGND.n2354 76.3222
R2576 VGND.n2358 VGND.n2357 76.3222
R2577 VGND.n2370 VGND.n2369 76.3222
R2578 VGND.n2373 VGND.n2372 76.3222
R2579 VGND.n2385 VGND.n2384 76.3222
R2580 VGND.n2341 VGND.n112 76.3222
R2581 VGND.n2356 VGND.n2355 76.3222
R2582 VGND.n2357 VGND.n107 76.3222
R2583 VGND.n2371 VGND.n2370 76.3222
R2584 VGND.n2372 VGND.n100 76.3222
R2585 VGND.n2386 VGND.n2385 76.3222
R2586 VGND.n2266 VGND.n2265 76.3222
R2587 VGND.n2088 VGND.n2087 76.3222
R2588 VGND.n2085 VGND.n2084 76.3222
R2589 VGND.n2082 VGND.n2081 76.3222
R2590 VGND.n2077 VGND.n2076 76.3222
R2591 VGND.n2074 VGND.n2013 76.3222
R2592 VGND.n2105 VGND.n2104 76.3222
R2593 VGND.n2100 VGND.n2073 76.3222
R2594 VGND.n2098 VGND.n2097 76.3222
R2595 VGND.n2093 VGND.n2092 76.3222
R2596 VGND.n2090 VGND.n460 76.3222
R2597 VGND.n2270 VGND.n2269 76.3222
R2598 VGND.n1528 VGND.n1527 76.3222
R2599 VGND.n1519 VGND.n1499 76.3222
R2600 VGND.n1513 VGND.n1498 76.3222
R2601 VGND.n1507 VGND.n1497 76.3222
R2602 VGND.n1502 VGND.n1496 76.3222
R2603 VGND.n1495 VGND.n744 76.3222
R2604 VGND.n1808 VGND.n748 76.3222
R2605 VGND.n1508 VGND.n753 76.3222
R2606 VGND.n1514 VGND.n752 76.3222
R2607 VGND.n1520 VGND.n751 76.3222
R2608 VGND.n1524 VGND.n750 76.3222
R2609 VGND.n789 VGND.n749 76.3222
R2610 VGND.t33 VGND.t53 74.8304
R2611 VGND.t156 VGND.t82 74.8304
R2612 VGND.t102 VGND.t298 74.8304
R2613 VGND.n1566 VGND.n825 74.5978
R2614 VGND.n1563 VGND.n825 74.5978
R2615 VGND.n503 VGND.n486 74.5978
R2616 VGND.n504 VGND.n503 74.5978
R2617 VGND.n1745 VGND.n767 74.5978
R2618 VGND.n1742 VGND.n767 74.5978
R2619 VGND.n303 VGND.n238 74.5978
R2620 VGND.n300 VGND.n238 74.5978
R2621 VGND.n420 VGND.n403 74.5978
R2622 VGND.n421 VGND.n420 74.5978
R2623 VGND.n1917 VGND.n678 74.5978
R2624 VGND.n1918 VGND.n1917 74.5978
R2625 VGND.n1201 VGND.n1144 74.5978
R2626 VGND.n1198 VGND.n1144 74.5978
R2627 VGND.n615 VGND.n598 74.5978
R2628 VGND.n616 VGND.n615 74.5978
R2629 VGND.n139 VGND.n122 74.5978
R2630 VGND.n140 VGND.n139 74.5978
R2631 VGND.n857 VGND.n8 74.09
R2632 VGND.n867 VGND.n866 74.09
R2633 VGND.n869 VGND.n853 74.09
R2634 VGND.n873 VGND.n872 74.09
R2635 VGND.n875 VGND.n874 74.09
R2636 VGND.n1359 VGND.n1358 74.09
R2637 VGND.n1361 VGND.n1339 74.09
R2638 VGND.n1343 VGND.n11 74.09
R2639 VGND.n1357 VGND.n1356 74.09
R2640 VGND.n1365 VGND.n1364 74.09
R2641 VGND.n882 VGND.n881 73.9572
R2642 VGND.n1381 VGND.n1016 73.9501
R2643 VGND.n1373 VGND.n1372 73.8434
R2644 VGND.n877 VGND.n852 73.3478
R2645 VGND.n881 VGND.n880 73.3478
R2646 VGND.n1367 VGND.n1366 72.7809
R2647 VGND.n1372 VGND.n1371 72.7809
R2648 VGND.n1375 VGND.t90 72.6135
R2649 VGND.n2455 VGND.n57 69.4466
R2650 VGND.n1614 VGND.n812 69.3109
R2651 VGND.n1585 VGND.n812 69.3109
R2652 VGND.n2225 VGND.n2224 69.3109
R2653 VGND.n2224 VGND.n2223 69.3109
R2654 VGND.n1800 VGND.n1799 69.3109
R2655 VGND.n1800 VGND.n778 69.3109
R2656 VGND.n337 VGND.n231 69.3109
R2657 VGND.n337 VGND.n336 69.3109
R2658 VGND.n2280 VGND.n2279 69.3109
R2659 VGND.n2279 VGND.n2278 69.3109
R2660 VGND.n1959 VGND.n1956 69.3109
R2661 VGND.n1956 VGND.n1955 69.3109
R2662 VGND.n1245 VGND.n1133 69.3109
R2663 VGND.n1220 VGND.n1133 69.3109
R2664 VGND.n2174 VGND.n2173 69.3109
R2665 VGND.n2173 VGND.n2172 69.3109
R2666 VGND.n2349 VGND.n2348 69.3109
R2667 VGND.n2348 VGND.n2347 69.3109
R2668 VGND.n1489 VGND.n1488 68.2005
R2669 VGND.n1468 VGND.n1467 68.2005
R2670 VGND.n863 VGND.n862 68.2005
R2671 VGND.n860 VGND.n856 68.2005
R2672 VGND.n1348 VGND.n1346 68.2005
R2673 VGND.n1352 VGND.n1351 68.2005
R2674 VGND.t218 VGND.n366 67.9598
R2675 VGND.n1433 VGND.n1432 66.5605
R2676 VGND.n1432 VGND.n935 66.5605
R2677 VGND.t259 VGND.n1599 65.8183
R2678 VGND.t259 VGND.n834 65.8183
R2679 VGND.t259 VGND.n833 65.8183
R2680 VGND.t259 VGND.n832 65.8183
R2681 VGND.t259 VGND.n823 65.8183
R2682 VGND.t259 VGND.n830 65.8183
R2683 VGND.t259 VGND.n821 65.8183
R2684 VGND.t259 VGND.n831 65.8183
R2685 VGND.t259 VGND.n829 65.8183
R2686 VGND.t259 VGND.n828 65.8183
R2687 VGND.t259 VGND.n827 65.8183
R2688 VGND.t259 VGND.n826 65.8183
R2689 VGND.t259 VGND.n824 65.8183
R2690 VGND.t259 VGND.n822 65.8183
R2691 VGND.n1602 VGND.t259 65.8183
R2692 VGND.t259 VGND.n813 65.8183
R2693 VGND.n525 VGND.t246 65.8183
R2694 VGND.n527 VGND.t246 65.8183
R2695 VGND.n533 VGND.t246 65.8183
R2696 VGND.n535 VGND.t246 65.8183
R2697 VGND.n509 VGND.t246 65.8183
R2698 VGND.n511 VGND.t246 65.8183
R2699 VGND.n517 VGND.t246 65.8183
R2700 VGND.n519 VGND.t246 65.8183
R2701 VGND.t246 VGND.n467 65.8183
R2702 VGND.n494 VGND.t246 65.8183
R2703 VGND.n490 VGND.t246 65.8183
R2704 VGND.n501 VGND.t246 65.8183
R2705 VGND.n2254 VGND.t246 65.8183
R2706 VGND.n2241 VGND.t246 65.8183
R2707 VGND.n2239 VGND.t246 65.8183
R2708 VGND.n2226 VGND.t246 65.8183
R2709 VGND.t215 VGND.n777 65.8183
R2710 VGND.t215 VGND.n776 65.8183
R2711 VGND.t215 VGND.n775 65.8183
R2712 VGND.t215 VGND.n774 65.8183
R2713 VGND.t215 VGND.n765 65.8183
R2714 VGND.t215 VGND.n772 65.8183
R2715 VGND.t215 VGND.n763 65.8183
R2716 VGND.t215 VGND.n773 65.8183
R2717 VGND.t215 VGND.n771 65.8183
R2718 VGND.t215 VGND.n770 65.8183
R2719 VGND.t215 VGND.n769 65.8183
R2720 VGND.t215 VGND.n768 65.8183
R2721 VGND.t215 VGND.n766 65.8183
R2722 VGND.n1801 VGND.t215 65.8183
R2723 VGND.t215 VGND.n764 65.8183
R2724 VGND.t215 VGND.n762 65.8183
R2725 VGND.t242 VGND.n248 65.8183
R2726 VGND.t242 VGND.n247 65.8183
R2727 VGND.t242 VGND.n246 65.8183
R2728 VGND.t242 VGND.n245 65.8183
R2729 VGND.t242 VGND.n236 65.8183
R2730 VGND.t242 VGND.n243 65.8183
R2731 VGND.t242 VGND.n233 65.8183
R2732 VGND.t242 VGND.n244 65.8183
R2733 VGND.t242 VGND.n242 65.8183
R2734 VGND.t242 VGND.n241 65.8183
R2735 VGND.t242 VGND.n240 65.8183
R2736 VGND.t242 VGND.n239 65.8183
R2737 VGND.t242 VGND.n237 65.8183
R2738 VGND.t242 VGND.n235 65.8183
R2739 VGND.t242 VGND.n234 65.8183
R2740 VGND.n338 VGND.t242 65.8183
R2741 VGND.n442 VGND.t258 65.8183
R2742 VGND.n444 VGND.t258 65.8183
R2743 VGND.n450 VGND.t258 65.8183
R2744 VGND.n452 VGND.t258 65.8183
R2745 VGND.n426 VGND.t258 65.8183
R2746 VGND.n428 VGND.t258 65.8183
R2747 VGND.n434 VGND.t258 65.8183
R2748 VGND.n436 VGND.t258 65.8183
R2749 VGND.t258 VGND.n384 65.8183
R2750 VGND.n411 VGND.t258 65.8183
R2751 VGND.n407 VGND.t258 65.8183
R2752 VGND.n418 VGND.t258 65.8183
R2753 VGND.n2309 VGND.t258 65.8183
R2754 VGND.n2296 VGND.t258 65.8183
R2755 VGND.n2294 VGND.t258 65.8183
R2756 VGND.n2281 VGND.t258 65.8183
R2757 VGND.n1939 VGND.t230 65.8183
R2758 VGND.n1941 VGND.t230 65.8183
R2759 VGND.n1947 VGND.t230 65.8183
R2760 VGND.n1949 VGND.t230 65.8183
R2761 VGND.n1923 VGND.t230 65.8183
R2762 VGND.n1925 VGND.t230 65.8183
R2763 VGND.n1931 VGND.t230 65.8183
R2764 VGND.n1933 VGND.t230 65.8183
R2765 VGND.n685 VGND.t230 65.8183
R2766 VGND.n1908 VGND.t230 65.8183
R2767 VGND.n682 VGND.t230 65.8183
R2768 VGND.n1915 VGND.t230 65.8183
R2769 VGND.n1901 VGND.t230 65.8183
R2770 VGND.n1888 VGND.t230 65.8183
R2771 VGND.n1886 VGND.t230 65.8183
R2772 VGND.n1961 VGND.t230 65.8183
R2773 VGND.t213 VGND.n1234 65.8183
R2774 VGND.t213 VGND.n1153 65.8183
R2775 VGND.t213 VGND.n1152 65.8183
R2776 VGND.t213 VGND.n1151 65.8183
R2777 VGND.t213 VGND.n1142 65.8183
R2778 VGND.t213 VGND.n1149 65.8183
R2779 VGND.t213 VGND.n1140 65.8183
R2780 VGND.t213 VGND.n1150 65.8183
R2781 VGND.t213 VGND.n1148 65.8183
R2782 VGND.t213 VGND.n1147 65.8183
R2783 VGND.t213 VGND.n1146 65.8183
R2784 VGND.t213 VGND.n1145 65.8183
R2785 VGND.t213 VGND.n1143 65.8183
R2786 VGND.t213 VGND.n1141 65.8183
R2787 VGND.n1235 VGND.t213 65.8183
R2788 VGND.t213 VGND.n1134 65.8183
R2789 VGND.n637 VGND.t217 65.8183
R2790 VGND.n639 VGND.t217 65.8183
R2791 VGND.n645 VGND.t217 65.8183
R2792 VGND.n647 VGND.t217 65.8183
R2793 VGND.n621 VGND.t217 65.8183
R2794 VGND.n623 VGND.t217 65.8183
R2795 VGND.n629 VGND.t217 65.8183
R2796 VGND.n631 VGND.t217 65.8183
R2797 VGND.t217 VGND.n579 65.8183
R2798 VGND.n606 VGND.t217 65.8183
R2799 VGND.n602 VGND.t217 65.8183
R2800 VGND.n613 VGND.t217 65.8183
R2801 VGND.n2203 VGND.t217 65.8183
R2802 VGND.n2190 VGND.t217 65.8183
R2803 VGND.n2188 VGND.t217 65.8183
R2804 VGND.n2175 VGND.t217 65.8183
R2805 VGND.n161 VGND.t266 65.8183
R2806 VGND.n163 VGND.t266 65.8183
R2807 VGND.n169 VGND.t266 65.8183
R2808 VGND.n171 VGND.t266 65.8183
R2809 VGND.n145 VGND.t266 65.8183
R2810 VGND.n147 VGND.t266 65.8183
R2811 VGND.n153 VGND.t266 65.8183
R2812 VGND.n155 VGND.t266 65.8183
R2813 VGND.t266 VGND.n103 65.8183
R2814 VGND.n130 VGND.t266 65.8183
R2815 VGND.n126 VGND.t266 65.8183
R2816 VGND.n137 VGND.t266 65.8183
R2817 VGND.n2378 VGND.t266 65.8183
R2818 VGND.n2365 VGND.t266 65.8183
R2819 VGND.n2363 VGND.t266 65.8183
R2820 VGND.n2350 VGND.t266 65.8183
R2821 VGND.t166 VGND.t39 64.8531
R2822 VGND.n1530 VGND.t218 62.176
R2823 VGND.t218 VGND.n1806 62.176
R2824 VGND.n991 VGND.t268 60.0005
R2825 VGND.n991 VGND.t103 60.0005
R2826 VGND.t249 VGND.n992 60.0005
R2827 VGND.n992 VGND.t40 60.0005
R2828 VGND.n990 VGND.t309 60.0005
R2829 VGND.n990 VGND.t221 60.0005
R2830 VGND.n933 VGND.t129 60.0005
R2831 VGND.n933 VGND.t67 60.0005
R2832 VGND.n932 VGND.t237 60.0005
R2833 VGND.n932 VGND.t159 60.0005
R2834 VGND.n934 VGND.t277 60.0005
R2835 VGND.n934 VGND.t240 60.0005
R2836 VGND.n1607 VGND.t45 59.2841
R2837 VGND.t259 VGND.n812 57.8461
R2838 VGND.n2224 VGND.t246 57.8461
R2839 VGND.t215 VGND.n1800 57.8461
R2840 VGND.t242 VGND.n337 57.8461
R2841 VGND.n2279 VGND.t258 57.8461
R2842 VGND.n1956 VGND.t230 57.8461
R2843 VGND.t213 VGND.n1133 57.8461
R2844 VGND.n2173 VGND.t217 57.8461
R2845 VGND.n2348 VGND.t266 57.8461
R2846 VGND.t218 VGND.t175 57.8382
R2847 VGND.t178 VGND.t218 57.8382
R2848 VGND.n2339 VGND.t214 56.5781
R2849 VGND.n1651 VGND.n1648 56.3995
R2850 VGND.n2319 VGND.n378 56.3995
R2851 VGND.n661 VGND.n652 56.3995
R2852 VGND.n1254 VGND.n1253 56.3995
R2853 VGND.n1971 VGND.n652 56.3995
R2854 VGND.n2165 VGND.n2164 56.3995
R2855 VGND.n1253 VGND.n224 56.3995
R2856 VGND.n1648 VGND.n1647 56.3995
R2857 VGND.n2319 VGND.n2318 56.3995
R2858 VGND.n2387 VGND.n96 56.3995
R2859 VGND.n2388 VGND.n2387 56.3995
R2860 VGND.n1408 VGND.n1407 55.4005
R2861 VGND.t259 VGND.n825 55.2026
R2862 VGND.n503 VGND.t246 55.2026
R2863 VGND.t215 VGND.n767 55.2026
R2864 VGND.t242 VGND.n238 55.2026
R2865 VGND.n420 VGND.t258 55.2026
R2866 VGND.n1917 VGND.t230 55.2026
R2867 VGND.t213 VGND.n1144 55.2026
R2868 VGND.n615 VGND.t217 55.2026
R2869 VGND.n139 VGND.t266 55.2026
R2870 VGND.t82 VGND.t33 54.8758
R2871 VGND.t275 VGND.t156 54.8758
R2872 VGND.t248 VGND.t261 54.8758
R2873 VGND.n1385 VGND.n1384 53.5422
R2874 VGND.n980 VGND.n972 53.5422
R2875 VGND.n1419 VGND.n1418 53.5422
R2876 VGND.n1421 VGND.n1420 53.5422
R2877 VGND.n970 VGND.n969 53.5422
R2878 VGND.n968 VGND.n967 53.5422
R2879 VGND.t209 VGND.n365 53.5003
R2880 VGND.n665 VGND.t210 53.5003
R2881 VGND.t87 VGND.n1895 53.5003
R2882 VGND.n1638 VGND.n793 53.5003
R2883 VGND.n2469 VGND.n2468 53.4593
R2884 VGND.n51 VGND.n41 53.4593
R2885 VGND.n1581 VGND.n831 53.3664
R2886 VGND.n1578 VGND.n821 53.3664
R2887 VGND.n1574 VGND.n830 53.3664
R2888 VGND.n1570 VGND.n823 53.3664
R2889 VGND.n1559 VGND.n826 53.3664
R2890 VGND.n1555 VGND.n827 53.3664
R2891 VGND.n1551 VGND.n828 53.3664
R2892 VGND.n1547 VGND.n829 53.3664
R2893 VGND.n1613 VGND.n813 53.3664
R2894 VGND.n1602 VGND.n1601 53.3664
R2895 VGND.n822 VGND.n820 53.3664
R2896 VGND.n1534 VGND.n824 53.3664
R2897 VGND.n1599 VGND.n1598 53.3664
R2898 VGND.n836 VGND.n834 53.3664
R2899 VGND.n1593 VGND.n833 53.3664
R2900 VGND.n1589 VGND.n832 53.3664
R2901 VGND.n1599 VGND.n835 53.3664
R2902 VGND.n1594 VGND.n834 53.3664
R2903 VGND.n1590 VGND.n833 53.3664
R2904 VGND.n1586 VGND.n832 53.3664
R2905 VGND.n1567 VGND.n823 53.3664
R2906 VGND.n1571 VGND.n830 53.3664
R2907 VGND.n1575 VGND.n821 53.3664
R2908 VGND.n1579 VGND.n831 53.3664
R2909 VGND.n1550 VGND.n829 53.3664
R2910 VGND.n1554 VGND.n828 53.3664
R2911 VGND.n1558 VGND.n827 53.3664
R2912 VGND.n1562 VGND.n826 53.3664
R2913 VGND.n1546 VGND.n824 53.3664
R2914 VGND.n1535 VGND.n822 53.3664
R2915 VGND.n1603 VGND.n1602 53.3664
R2916 VGND.n1600 VGND.n813 53.3664
R2917 VGND.n519 VGND.n482 53.3664
R2918 VGND.n518 VGND.n517 53.3664
R2919 VGND.n511 VGND.n484 53.3664
R2920 VGND.n510 VGND.n509 53.3664
R2921 VGND.n501 VGND.n500 53.3664
R2922 VGND.n496 VGND.n490 53.3664
R2923 VGND.n494 VGND.n493 53.3664
R2924 VGND.n2256 VGND.n467 53.3664
R2925 VGND.n2227 VGND.n2226 53.3664
R2926 VGND.n2239 VGND.n2238 53.3664
R2927 VGND.n2242 VGND.n2241 53.3664
R2928 VGND.n2254 VGND.n2253 53.3664
R2929 VGND.n526 VGND.n525 53.3664
R2930 VGND.n528 VGND.n527 53.3664
R2931 VGND.n533 VGND.n532 53.3664
R2932 VGND.n536 VGND.n535 53.3664
R2933 VGND.n525 VGND.n524 53.3664
R2934 VGND.n527 VGND.n480 53.3664
R2935 VGND.n534 VGND.n533 53.3664
R2936 VGND.n535 VGND.n478 53.3664
R2937 VGND.n509 VGND.n508 53.3664
R2938 VGND.n512 VGND.n511 53.3664
R2939 VGND.n517 VGND.n516 53.3664
R2940 VGND.n520 VGND.n519 53.3664
R2941 VGND.n491 VGND.n467 53.3664
R2942 VGND.n495 VGND.n494 53.3664
R2943 VGND.n490 VGND.n488 53.3664
R2944 VGND.n502 VGND.n501 53.3664
R2945 VGND.n2255 VGND.n2254 53.3664
R2946 VGND.n2241 VGND.n468 53.3664
R2947 VGND.n2240 VGND.n2239 53.3664
R2948 VGND.n2226 VGND.n473 53.3664
R2949 VGND.n1761 VGND.n773 53.3664
R2950 VGND.n1757 VGND.n763 53.3664
R2951 VGND.n1753 VGND.n772 53.3664
R2952 VGND.n1749 VGND.n765 53.3664
R2953 VGND.n1738 VGND.n768 53.3664
R2954 VGND.n1734 VGND.n769 53.3664
R2955 VGND.n1730 VGND.n770 53.3664
R2956 VGND.n1726 VGND.n771 53.3664
R2957 VGND.n779 VGND.n762 53.3664
R2958 VGND.n1789 VGND.n764 53.3664
R2959 VGND.n1802 VGND.n1801 53.3664
R2960 VGND.n1714 VGND.n766 53.3664
R2961 VGND.n1765 VGND.n777 53.3664
R2962 VGND.n1766 VGND.n776 53.3664
R2963 VGND.n1770 VGND.n775 53.3664
R2964 VGND.n1774 VGND.n774 53.3664
R2965 VGND.n1762 VGND.n777 53.3664
R2966 VGND.n1769 VGND.n776 53.3664
R2967 VGND.n1773 VGND.n775 53.3664
R2968 VGND.n1776 VGND.n774 53.3664
R2969 VGND.n1746 VGND.n765 53.3664
R2970 VGND.n1750 VGND.n772 53.3664
R2971 VGND.n1754 VGND.n763 53.3664
R2972 VGND.n1758 VGND.n773 53.3664
R2973 VGND.n1729 VGND.n771 53.3664
R2974 VGND.n1733 VGND.n770 53.3664
R2975 VGND.n1737 VGND.n769 53.3664
R2976 VGND.n1741 VGND.n768 53.3664
R2977 VGND.n1725 VGND.n766 53.3664
R2978 VGND.n1801 VGND.n761 53.3664
R2979 VGND.n764 VGND.n760 53.3664
R2980 VGND.n1788 VGND.n762 53.3664
R2981 VGND.n319 VGND.n244 53.3664
R2982 VGND.n315 VGND.n233 53.3664
R2983 VGND.n311 VGND.n243 53.3664
R2984 VGND.n307 VGND.n236 53.3664
R2985 VGND.n296 VGND.n239 53.3664
R2986 VGND.n292 VGND.n240 53.3664
R2987 VGND.n288 VGND.n241 53.3664
R2988 VGND.n284 VGND.n242 53.3664
R2989 VGND.n339 VGND.n338 53.3664
R2990 VGND.n253 VGND.n234 53.3664
R2991 VGND.n266 VGND.n235 53.3664
R2992 VGND.n271 VGND.n237 53.3664
R2993 VGND.n323 VGND.n248 53.3664
R2994 VGND.n324 VGND.n247 53.3664
R2995 VGND.n328 VGND.n246 53.3664
R2996 VGND.n332 VGND.n245 53.3664
R2997 VGND.n320 VGND.n248 53.3664
R2998 VGND.n327 VGND.n247 53.3664
R2999 VGND.n331 VGND.n246 53.3664
R3000 VGND.n335 VGND.n245 53.3664
R3001 VGND.n304 VGND.n236 53.3664
R3002 VGND.n308 VGND.n243 53.3664
R3003 VGND.n312 VGND.n233 53.3664
R3004 VGND.n316 VGND.n244 53.3664
R3005 VGND.n287 VGND.n242 53.3664
R3006 VGND.n291 VGND.n241 53.3664
R3007 VGND.n295 VGND.n240 53.3664
R3008 VGND.n299 VGND.n239 53.3664
R3009 VGND.n283 VGND.n237 53.3664
R3010 VGND.n270 VGND.n235 53.3664
R3011 VGND.n265 VGND.n234 53.3664
R3012 VGND.n338 VGND.n232 53.3664
R3013 VGND.n436 VGND.n399 53.3664
R3014 VGND.n435 VGND.n434 53.3664
R3015 VGND.n428 VGND.n401 53.3664
R3016 VGND.n427 VGND.n426 53.3664
R3017 VGND.n418 VGND.n417 53.3664
R3018 VGND.n413 VGND.n407 53.3664
R3019 VGND.n411 VGND.n410 53.3664
R3020 VGND.n2311 VGND.n384 53.3664
R3021 VGND.n2282 VGND.n2281 53.3664
R3022 VGND.n2294 VGND.n2293 53.3664
R3023 VGND.n2297 VGND.n2296 53.3664
R3024 VGND.n2309 VGND.n2308 53.3664
R3025 VGND.n443 VGND.n442 53.3664
R3026 VGND.n445 VGND.n444 53.3664
R3027 VGND.n450 VGND.n449 53.3664
R3028 VGND.n453 VGND.n452 53.3664
R3029 VGND.n442 VGND.n441 53.3664
R3030 VGND.n444 VGND.n397 53.3664
R3031 VGND.n451 VGND.n450 53.3664
R3032 VGND.n452 VGND.n395 53.3664
R3033 VGND.n426 VGND.n425 53.3664
R3034 VGND.n429 VGND.n428 53.3664
R3035 VGND.n434 VGND.n433 53.3664
R3036 VGND.n437 VGND.n436 53.3664
R3037 VGND.n408 VGND.n384 53.3664
R3038 VGND.n412 VGND.n411 53.3664
R3039 VGND.n407 VGND.n405 53.3664
R3040 VGND.n419 VGND.n418 53.3664
R3041 VGND.n2310 VGND.n2309 53.3664
R3042 VGND.n2296 VGND.n385 53.3664
R3043 VGND.n2295 VGND.n2294 53.3664
R3044 VGND.n2281 VGND.n390 53.3664
R3045 VGND.n1933 VGND.n674 53.3664
R3046 VGND.n1932 VGND.n1931 53.3664
R3047 VGND.n1925 VGND.n676 53.3664
R3048 VGND.n1924 VGND.n1923 53.3664
R3049 VGND.n1915 VGND.n1914 53.3664
R3050 VGND.n1910 VGND.n682 53.3664
R3051 VGND.n1908 VGND.n1907 53.3664
R3052 VGND.n1903 VGND.n685 53.3664
R3053 VGND.n1961 VGND.n1960 53.3664
R3054 VGND.n1886 VGND.n669 53.3664
R3055 VGND.n1889 VGND.n1888 53.3664
R3056 VGND.n1901 VGND.n1900 53.3664
R3057 VGND.n1940 VGND.n1939 53.3664
R3058 VGND.n1942 VGND.n1941 53.3664
R3059 VGND.n1947 VGND.n1946 53.3664
R3060 VGND.n1950 VGND.n1949 53.3664
R3061 VGND.n1939 VGND.n1938 53.3664
R3062 VGND.n1941 VGND.n672 53.3664
R3063 VGND.n1948 VGND.n1947 53.3664
R3064 VGND.n1949 VGND.n670 53.3664
R3065 VGND.n1923 VGND.n1922 53.3664
R3066 VGND.n1926 VGND.n1925 53.3664
R3067 VGND.n1931 VGND.n1930 53.3664
R3068 VGND.n1934 VGND.n1933 53.3664
R3069 VGND.n685 VGND.n683 53.3664
R3070 VGND.n1909 VGND.n1908 53.3664
R3071 VGND.n682 VGND.n680 53.3664
R3072 VGND.n1916 VGND.n1915 53.3664
R3073 VGND.n1902 VGND.n1901 53.3664
R3074 VGND.n1888 VGND.n687 53.3664
R3075 VGND.n1887 VGND.n1886 53.3664
R3076 VGND.n1962 VGND.n1961 53.3664
R3077 VGND.n1216 VGND.n1150 53.3664
R3078 VGND.n1213 VGND.n1140 53.3664
R3079 VGND.n1209 VGND.n1149 53.3664
R3080 VGND.n1205 VGND.n1142 53.3664
R3081 VGND.n1194 VGND.n1145 53.3664
R3082 VGND.n1190 VGND.n1146 53.3664
R3083 VGND.n1186 VGND.n1147 53.3664
R3084 VGND.n1182 VGND.n1148 53.3664
R3085 VGND.n1244 VGND.n1134 53.3664
R3086 VGND.n1236 VGND.n1235 53.3664
R3087 VGND.n1164 VGND.n1141 53.3664
R3088 VGND.n1169 VGND.n1143 53.3664
R3089 VGND.n1234 VGND.n1233 53.3664
R3090 VGND.n1155 VGND.n1153 53.3664
R3091 VGND.n1228 VGND.n1152 53.3664
R3092 VGND.n1224 VGND.n1151 53.3664
R3093 VGND.n1234 VGND.n1154 53.3664
R3094 VGND.n1229 VGND.n1153 53.3664
R3095 VGND.n1225 VGND.n1152 53.3664
R3096 VGND.n1221 VGND.n1151 53.3664
R3097 VGND.n1202 VGND.n1142 53.3664
R3098 VGND.n1206 VGND.n1149 53.3664
R3099 VGND.n1210 VGND.n1140 53.3664
R3100 VGND.n1214 VGND.n1150 53.3664
R3101 VGND.n1185 VGND.n1148 53.3664
R3102 VGND.n1189 VGND.n1147 53.3664
R3103 VGND.n1193 VGND.n1146 53.3664
R3104 VGND.n1197 VGND.n1145 53.3664
R3105 VGND.n1181 VGND.n1143 53.3664
R3106 VGND.n1168 VGND.n1141 53.3664
R3107 VGND.n1235 VGND.n1139 53.3664
R3108 VGND.n1138 VGND.n1134 53.3664
R3109 VGND.n631 VGND.n594 53.3664
R3110 VGND.n630 VGND.n629 53.3664
R3111 VGND.n623 VGND.n596 53.3664
R3112 VGND.n622 VGND.n621 53.3664
R3113 VGND.n613 VGND.n612 53.3664
R3114 VGND.n608 VGND.n602 53.3664
R3115 VGND.n606 VGND.n605 53.3664
R3116 VGND.n2205 VGND.n579 53.3664
R3117 VGND.n2176 VGND.n2175 53.3664
R3118 VGND.n2188 VGND.n2187 53.3664
R3119 VGND.n2191 VGND.n2190 53.3664
R3120 VGND.n2203 VGND.n2202 53.3664
R3121 VGND.n638 VGND.n637 53.3664
R3122 VGND.n640 VGND.n639 53.3664
R3123 VGND.n645 VGND.n644 53.3664
R3124 VGND.n648 VGND.n647 53.3664
R3125 VGND.n637 VGND.n636 53.3664
R3126 VGND.n639 VGND.n592 53.3664
R3127 VGND.n646 VGND.n645 53.3664
R3128 VGND.n647 VGND.n590 53.3664
R3129 VGND.n621 VGND.n620 53.3664
R3130 VGND.n624 VGND.n623 53.3664
R3131 VGND.n629 VGND.n628 53.3664
R3132 VGND.n632 VGND.n631 53.3664
R3133 VGND.n603 VGND.n579 53.3664
R3134 VGND.n607 VGND.n606 53.3664
R3135 VGND.n602 VGND.n600 53.3664
R3136 VGND.n614 VGND.n613 53.3664
R3137 VGND.n2204 VGND.n2203 53.3664
R3138 VGND.n2190 VGND.n580 53.3664
R3139 VGND.n2189 VGND.n2188 53.3664
R3140 VGND.n2175 VGND.n585 53.3664
R3141 VGND.n155 VGND.n118 53.3664
R3142 VGND.n154 VGND.n153 53.3664
R3143 VGND.n147 VGND.n120 53.3664
R3144 VGND.n146 VGND.n145 53.3664
R3145 VGND.n137 VGND.n136 53.3664
R3146 VGND.n132 VGND.n126 53.3664
R3147 VGND.n130 VGND.n129 53.3664
R3148 VGND.n2380 VGND.n103 53.3664
R3149 VGND.n2351 VGND.n2350 53.3664
R3150 VGND.n2363 VGND.n2362 53.3664
R3151 VGND.n2366 VGND.n2365 53.3664
R3152 VGND.n2378 VGND.n2377 53.3664
R3153 VGND.n162 VGND.n161 53.3664
R3154 VGND.n164 VGND.n163 53.3664
R3155 VGND.n169 VGND.n168 53.3664
R3156 VGND.n172 VGND.n171 53.3664
R3157 VGND.n161 VGND.n160 53.3664
R3158 VGND.n163 VGND.n116 53.3664
R3159 VGND.n170 VGND.n169 53.3664
R3160 VGND.n171 VGND.n114 53.3664
R3161 VGND.n145 VGND.n144 53.3664
R3162 VGND.n148 VGND.n147 53.3664
R3163 VGND.n153 VGND.n152 53.3664
R3164 VGND.n156 VGND.n155 53.3664
R3165 VGND.n127 VGND.n103 53.3664
R3166 VGND.n131 VGND.n130 53.3664
R3167 VGND.n126 VGND.n124 53.3664
R3168 VGND.n138 VGND.n137 53.3664
R3169 VGND.n2379 VGND.n2378 53.3664
R3170 VGND.n2365 VGND.n104 53.3664
R3171 VGND.n2364 VGND.n2363 53.3664
R3172 VGND.n2350 VGND.n109 53.3664
R3173 VGND.n1432 VGND.n1431 53.3255
R3174 VGND.n2482 VGND.n2472 52.3299
R3175 VGND.n0 VGND.t218 21.2213
R3176 VGND.t153 VGND.t183 49.8871
R3177 VGND.t232 VGND.t255 49.8871
R3178 VGND.n4 VGND.t114 48.0005
R3179 VGND.n4 VGND.t169 48.0005
R3180 VGND.n1475 VGND.t315 48.0005
R3181 VGND.n1475 VGND.t30 48.0005
R3182 VGND.n1478 VGND.t304 48.0005
R3183 VGND.n1478 VGND.t295 48.0005
R3184 VGND.n1480 VGND.t61 48.0005
R3185 VGND.n1480 VGND.t152 48.0005
R3186 VGND.n1482 VGND.t65 48.0005
R3187 VGND.n1482 VGND.t84 48.0005
R3188 VGND.n1484 VGND.t21 48.0005
R3189 VGND.n1484 VGND.t319 48.0005
R3190 VGND.n1486 VGND.t131 48.0005
R3191 VGND.n1486 VGND.t121 48.0005
R3192 VGND.n1471 VGND.t52 48.0005
R3193 VGND.n1471 VGND.t105 48.0005
R3194 VGND.n1469 VGND.t165 48.0005
R3195 VGND.n1469 VGND.t3 48.0005
R3196 VGND.n847 VGND.t13 48.0005
R3197 VGND.n847 VGND.t59 48.0005
R3198 VGND.n1460 VGND.t163 48.0005
R3199 VGND.n1460 VGND.t50 48.0005
R3200 VGND.n1462 VGND.t172 48.0005
R3201 VGND.n1462 VGND.t189 48.0005
R3202 VGND.n1458 VGND.t123 48.0005
R3203 VGND.n1458 VGND.t174 48.0005
R3204 VGND.n1456 VGND.t99 48.0005
R3205 VGND.n1456 VGND.t93 48.0005
R3206 VGND.n1454 VGND.t112 48.0005
R3207 VGND.n1454 VGND.t55 48.0005
R3208 VGND.n849 VGND.t290 48.0005
R3209 VGND.n849 VGND.t24 48.0005
R3210 VGND.n1446 VGND.t203 48.0005
R3211 VGND.n1446 VGND.t273 48.0005
R3212 VGND.n1448 VGND.t107 48.0005
R3213 VGND.n1448 VGND.t80 48.0005
R3214 VGND.n1444 VGND.t57 48.0005
R3215 VGND.n1444 VGND.t201 48.0005
R3216 VGND.n1442 VGND.t207 48.0005
R3217 VGND.n1442 VGND.t73 48.0005
R3218 VGND.n1441 VGND.t271 48.0005
R3219 VGND.n1441 VGND.t1 48.0005
R3220 VGND.n1621 VGND.n1618 47.7166
R3221 VGND.t117 VGND.n1794 47.7166
R3222 VGND.n1712 VGND.t177 47.7166
R3223 VGND.t74 VGND.n1720 47.7166
R3224 VGND.n2508 VGND.n2507 46.2505
R3225 VGND.n2504 VGND.n2500 46.2505
R3226 VGND.n2490 VGND.n2489 46.2505
R3227 VGND.n2494 VGND.n2493 46.2505
R3228 VGND.n34 VGND.n29 46.2505
R3229 VGND.n30 VGND.n28 46.2505
R3230 VGND.n22 VGND.n21 46.2505
R3231 VGND.n26 VGND.n25 46.2505
R3232 VGND.n1285 VGND.n1282 46.2505
R3233 VGND.n1289 VGND.n1283 46.2505
R3234 VGND.n1007 VGND.n1006 46.2505
R3235 VGND.n1011 VGND.n1010 46.2505
R3236 VGND.t228 VGND.t158 44.8985
R3237 VGND.t22 VGND.t153 44.8985
R3238 VGND.n1412 VGND.n989 44.8985
R3239 VGND.n886 VGND.t323 44.7909
R3240 VGND.n2493 VGND.n2487 43.856
R3241 VGND.n2491 VGND.n2490 43.856
R3242 VGND.n25 VGND.n19 43.856
R3243 VGND.n23 VGND.n22 43.856
R3244 VGND.n1285 VGND.n1284 43.3691
R3245 VGND.n1289 VGND.n1288 43.3691
R3246 VGND.n32 VGND.n30 43.2747
R3247 VGND.n35 VGND.n34 43.2747
R3248 VGND.n1008 VGND.n1007 43.1853
R3249 VGND.n1010 VGND.n1009 43.1853
R3250 VGND.n39 VGND.t288 42.9191
R3251 VGND.n1401 VGND.n1400 39.9098
R3252 VGND.n786 VGND.t182 39.0409
R3253 VGND.t196 VGND.n1783 39.0409
R3254 VGND.n1784 VGND.t269 39.0409
R3255 VGND.t274 VGND.n1719 39.0409
R3256 VGND.n1375 VGND.n1374 38.1958
R3257 VGND.n1875 VGND.t44 37.595
R3258 VGND.t236 VGND.n930 34.9211
R3259 VGND.t239 VGND.t193 34.9211
R3260 VGND.t183 VGND.t7 34.9211
R3261 VGND.t293 VGND.n1967 33.2572
R3262 VGND.n1879 VGND.t212 33.2572
R3263 VGND.n1877 VGND.t211 33.2572
R3264 VGND.n1313 VGND.n1312 33.0525
R3265 VGND.t218 VGND.n364 32.9056
R3266 VGND.n1332 VGND.n1331 32.3962
R3267 VGND.t27 VGND.t251 29.9325
R3268 VGND.t298 VGND.t108 29.9325
R3269 VGND.t218 VGND.n365 28.9193
R3270 VGND.t218 VGND.t212 28.9193
R3271 VGND.t175 VGND.t44 28.9193
R3272 VGND.t182 VGND.t178 28.9193
R3273 VGND.t218 VGND.t269 28.9193
R3274 VGND.t278 VGND.n1369 28.2933
R3275 VGND.n1583 VGND.n1582 27.5561
R3276 VGND.n523 VGND.n522 27.5561
R3277 VGND.n1763 VGND.n1760 27.5561
R3278 VGND.n321 VGND.n318 27.5561
R3279 VGND.n440 VGND.n439 27.5561
R3280 VGND.n1937 VGND.n1936 27.5561
R3281 VGND.n1218 VGND.n1217 27.5561
R3282 VGND.n635 VGND.n634 27.5561
R3283 VGND.n159 VGND.n158 27.5561
R3284 VGND.n938 VGND.n937 27.2005
R3285 VGND.n1435 VGND.n1434 27.2005
R3286 VGND.n1565 VGND.n1564 26.6672
R3287 VGND.n506 VGND.n505 26.6672
R3288 VGND.n1744 VGND.n1743 26.6672
R3289 VGND.n302 VGND.n301 26.6672
R3290 VGND.n423 VGND.n422 26.6672
R3291 VGND.n1920 VGND.n1919 26.6672
R3292 VGND.n1200 VGND.n1199 26.6672
R3293 VGND.n618 VGND.n617 26.6672
R3294 VGND.n142 VGND.n141 26.6672
R3295 VGND.n1411 VGND.n1410 25.6005
R3296 VGND.n994 VGND.n993 25.6005
R3297 VGND.n1319 VGND.n1318 25.3679
R3298 VGND.n2339 VGND.n99 25.0252
R3299 VGND.t108 VGND.t308 24.9438
R3300 VGND.n1403 VGND.n1402 24.8279
R3301 VGND.n1430 VGND.n1429 24.8279
R3302 VGND.n1405 VGND.t299 24.0005
R3303 VGND.n1405 VGND.t233 24.0005
R3304 VGND.n1000 VGND.t167 24.0005
R3305 VGND.n1000 VGND.t313 24.0005
R3306 VGND.n998 VGND.t28 24.0005
R3307 VGND.n998 VGND.t126 24.0005
R3308 VGND.n996 VGND.t306 24.0005
R3309 VGND.n996 VGND.t154 24.0005
R3310 VGND.t265 VGND.n1428 24.0005
R3311 VGND.n1428 VGND.t34 24.0005
R3312 VGND.n1293 VGND.n1292 22.6374
R3313 VGND.n1013 VGND.n1012 22.6374
R3314 VGND.n898 VGND.n889 22.4005
R3315 VGND.n904 VGND.n902 21.3338
R3316 VGND.n893 VGND.n891 21.3338
R3317 VGND.n917 VGND.n915 21.3338
R3318 VGND.n2474 VGND.n2473 20.5561
R3319 VGND.n2475 VGND.n2472 20.5561
R3320 VGND.n2468 VGND.n2467 20.5561
R3321 VGND.n2464 VGND.n2462 20.5561
R3322 VGND.n43 VGND.n42 20.5561
R3323 VGND.n44 VGND.n41 20.5561
R3324 VGND.t224 VGND.n939 19.9551
R3325 VGND.n1413 VGND.t125 19.9551
R3326 VGND.n907 VGND.n906 19.3862
R3327 VGND.n896 VGND.n895 19.3862
R3328 VGND.n920 VGND.n919 19.3862
R3329 VGND.n1688 VGND.n1659 17.5843
R3330 VGND.n2049 VGND.n2033 17.5843
R3331 VGND.n2411 VGND.n81 17.5843
R3332 VGND.n1400 VGND.n1399 17.2893
R3333 VGND.n2453 VGND.n2452 16.9605
R3334 VGND.n1991 VGND.n660 16.9379
R3335 VGND.n1276 VGND.n1121 16.9379
R3336 VGND.n2143 VGND.n2000 16.9379
R3337 VGND.n737 VGND.n540 16.7709
R3338 VGND.n2337 VGND.n2336 16.7709
R3339 VGND.n2108 VGND.n177 16.7709
R3340 VGND.n1811 VGND.n458 16.7709
R3341 VGND.n905 VGND.t279 16.0005
R3342 VGND.n894 VGND.t181 16.0005
R3343 VGND.n1597 VGND.n1583 16.0005
R3344 VGND.n1597 VGND.n1596 16.0005
R3345 VGND.n1596 VGND.n1595 16.0005
R3346 VGND.n1595 VGND.n1592 16.0005
R3347 VGND.n1592 VGND.n1591 16.0005
R3348 VGND.n1591 VGND.n1588 16.0005
R3349 VGND.n1588 VGND.n1587 16.0005
R3350 VGND.n1587 VGND.n1584 16.0005
R3351 VGND.n1582 VGND.n1580 16.0005
R3352 VGND.n1580 VGND.n1577 16.0005
R3353 VGND.n1577 VGND.n1576 16.0005
R3354 VGND.n1576 VGND.n1573 16.0005
R3355 VGND.n1573 VGND.n1572 16.0005
R3356 VGND.n1572 VGND.n1569 16.0005
R3357 VGND.n1569 VGND.n1568 16.0005
R3358 VGND.n1568 VGND.n1565 16.0005
R3359 VGND.n1564 VGND.n1561 16.0005
R3360 VGND.n1561 VGND.n1560 16.0005
R3361 VGND.n1560 VGND.n1557 16.0005
R3362 VGND.n1557 VGND.n1556 16.0005
R3363 VGND.n1556 VGND.n1553 16.0005
R3364 VGND.n1553 VGND.n1552 16.0005
R3365 VGND.n1552 VGND.n1549 16.0005
R3366 VGND.n1549 VGND.n1548 16.0005
R3367 VGND.n523 VGND.n481 16.0005
R3368 VGND.n529 VGND.n481 16.0005
R3369 VGND.n530 VGND.n529 16.0005
R3370 VGND.n531 VGND.n530 16.0005
R3371 VGND.n531 VGND.n479 16.0005
R3372 VGND.n537 VGND.n479 16.0005
R3373 VGND.n538 VGND.n537 16.0005
R3374 VGND.n2222 VGND.n538 16.0005
R3375 VGND.n522 VGND.n521 16.0005
R3376 VGND.n521 VGND.n483 16.0005
R3377 VGND.n515 VGND.n483 16.0005
R3378 VGND.n515 VGND.n514 16.0005
R3379 VGND.n514 VGND.n513 16.0005
R3380 VGND.n513 VGND.n485 16.0005
R3381 VGND.n507 VGND.n485 16.0005
R3382 VGND.n507 VGND.n506 16.0005
R3383 VGND.n505 VGND.n487 16.0005
R3384 VGND.n499 VGND.n487 16.0005
R3385 VGND.n499 VGND.n498 16.0005
R3386 VGND.n498 VGND.n497 16.0005
R3387 VGND.n497 VGND.n489 16.0005
R3388 VGND.n492 VGND.n489 16.0005
R3389 VGND.n492 VGND.n466 16.0005
R3390 VGND.n2257 VGND.n466 16.0005
R3391 VGND.n1764 VGND.n1763 16.0005
R3392 VGND.n1767 VGND.n1764 16.0005
R3393 VGND.n1768 VGND.n1767 16.0005
R3394 VGND.n1771 VGND.n1768 16.0005
R3395 VGND.n1772 VGND.n1771 16.0005
R3396 VGND.n1775 VGND.n1772 16.0005
R3397 VGND.n1777 VGND.n1775 16.0005
R3398 VGND.n1778 VGND.n1777 16.0005
R3399 VGND.n1760 VGND.n1759 16.0005
R3400 VGND.n1759 VGND.n1756 16.0005
R3401 VGND.n1756 VGND.n1755 16.0005
R3402 VGND.n1755 VGND.n1752 16.0005
R3403 VGND.n1752 VGND.n1751 16.0005
R3404 VGND.n1751 VGND.n1748 16.0005
R3405 VGND.n1748 VGND.n1747 16.0005
R3406 VGND.n1747 VGND.n1744 16.0005
R3407 VGND.n1743 VGND.n1740 16.0005
R3408 VGND.n1740 VGND.n1739 16.0005
R3409 VGND.n1739 VGND.n1736 16.0005
R3410 VGND.n1736 VGND.n1735 16.0005
R3411 VGND.n1735 VGND.n1732 16.0005
R3412 VGND.n1732 VGND.n1731 16.0005
R3413 VGND.n1731 VGND.n1728 16.0005
R3414 VGND.n1728 VGND.n1727 16.0005
R3415 VGND.n322 VGND.n321 16.0005
R3416 VGND.n325 VGND.n322 16.0005
R3417 VGND.n326 VGND.n325 16.0005
R3418 VGND.n329 VGND.n326 16.0005
R3419 VGND.n330 VGND.n329 16.0005
R3420 VGND.n333 VGND.n330 16.0005
R3421 VGND.n334 VGND.n333 16.0005
R3422 VGND.n334 VGND.n227 16.0005
R3423 VGND.n318 VGND.n317 16.0005
R3424 VGND.n317 VGND.n314 16.0005
R3425 VGND.n314 VGND.n313 16.0005
R3426 VGND.n313 VGND.n310 16.0005
R3427 VGND.n310 VGND.n309 16.0005
R3428 VGND.n309 VGND.n306 16.0005
R3429 VGND.n306 VGND.n305 16.0005
R3430 VGND.n305 VGND.n302 16.0005
R3431 VGND.n301 VGND.n298 16.0005
R3432 VGND.n298 VGND.n297 16.0005
R3433 VGND.n297 VGND.n294 16.0005
R3434 VGND.n294 VGND.n293 16.0005
R3435 VGND.n293 VGND.n290 16.0005
R3436 VGND.n290 VGND.n289 16.0005
R3437 VGND.n289 VGND.n286 16.0005
R3438 VGND.n286 VGND.n285 16.0005
R3439 VGND.n440 VGND.n398 16.0005
R3440 VGND.n446 VGND.n398 16.0005
R3441 VGND.n447 VGND.n446 16.0005
R3442 VGND.n448 VGND.n447 16.0005
R3443 VGND.n448 VGND.n396 16.0005
R3444 VGND.n454 VGND.n396 16.0005
R3445 VGND.n455 VGND.n454 16.0005
R3446 VGND.n2277 VGND.n455 16.0005
R3447 VGND.n439 VGND.n438 16.0005
R3448 VGND.n438 VGND.n400 16.0005
R3449 VGND.n432 VGND.n400 16.0005
R3450 VGND.n432 VGND.n431 16.0005
R3451 VGND.n431 VGND.n430 16.0005
R3452 VGND.n430 VGND.n402 16.0005
R3453 VGND.n424 VGND.n402 16.0005
R3454 VGND.n424 VGND.n423 16.0005
R3455 VGND.n422 VGND.n404 16.0005
R3456 VGND.n416 VGND.n404 16.0005
R3457 VGND.n416 VGND.n415 16.0005
R3458 VGND.n415 VGND.n414 16.0005
R3459 VGND.n414 VGND.n406 16.0005
R3460 VGND.n409 VGND.n406 16.0005
R3461 VGND.n409 VGND.n383 16.0005
R3462 VGND.n2312 VGND.n383 16.0005
R3463 VGND.n1937 VGND.n673 16.0005
R3464 VGND.n1943 VGND.n673 16.0005
R3465 VGND.n1944 VGND.n1943 16.0005
R3466 VGND.n1945 VGND.n1944 16.0005
R3467 VGND.n1945 VGND.n671 16.0005
R3468 VGND.n1951 VGND.n671 16.0005
R3469 VGND.n1952 VGND.n1951 16.0005
R3470 VGND.n1954 VGND.n1952 16.0005
R3471 VGND.n1936 VGND.n1935 16.0005
R3472 VGND.n1935 VGND.n675 16.0005
R3473 VGND.n1929 VGND.n675 16.0005
R3474 VGND.n1929 VGND.n1928 16.0005
R3475 VGND.n1928 VGND.n1927 16.0005
R3476 VGND.n1927 VGND.n677 16.0005
R3477 VGND.n1921 VGND.n677 16.0005
R3478 VGND.n1921 VGND.n1920 16.0005
R3479 VGND.n1919 VGND.n679 16.0005
R3480 VGND.n1913 VGND.n679 16.0005
R3481 VGND.n1913 VGND.n1912 16.0005
R3482 VGND.n1912 VGND.n1911 16.0005
R3483 VGND.n1911 VGND.n681 16.0005
R3484 VGND.n1906 VGND.n681 16.0005
R3485 VGND.n1906 VGND.n1905 16.0005
R3486 VGND.n1905 VGND.n1904 16.0005
R3487 VGND.n1232 VGND.n1218 16.0005
R3488 VGND.n1232 VGND.n1231 16.0005
R3489 VGND.n1231 VGND.n1230 16.0005
R3490 VGND.n1230 VGND.n1227 16.0005
R3491 VGND.n1227 VGND.n1226 16.0005
R3492 VGND.n1226 VGND.n1223 16.0005
R3493 VGND.n1223 VGND.n1222 16.0005
R3494 VGND.n1222 VGND.n1219 16.0005
R3495 VGND.n1217 VGND.n1215 16.0005
R3496 VGND.n1215 VGND.n1212 16.0005
R3497 VGND.n1212 VGND.n1211 16.0005
R3498 VGND.n1211 VGND.n1208 16.0005
R3499 VGND.n1208 VGND.n1207 16.0005
R3500 VGND.n1207 VGND.n1204 16.0005
R3501 VGND.n1204 VGND.n1203 16.0005
R3502 VGND.n1203 VGND.n1200 16.0005
R3503 VGND.n1199 VGND.n1196 16.0005
R3504 VGND.n1196 VGND.n1195 16.0005
R3505 VGND.n1195 VGND.n1192 16.0005
R3506 VGND.n1192 VGND.n1191 16.0005
R3507 VGND.n1191 VGND.n1188 16.0005
R3508 VGND.n1188 VGND.n1187 16.0005
R3509 VGND.n1187 VGND.n1184 16.0005
R3510 VGND.n1184 VGND.n1183 16.0005
R3511 VGND.n635 VGND.n593 16.0005
R3512 VGND.n641 VGND.n593 16.0005
R3513 VGND.n642 VGND.n641 16.0005
R3514 VGND.n643 VGND.n642 16.0005
R3515 VGND.n643 VGND.n591 16.0005
R3516 VGND.n649 VGND.n591 16.0005
R3517 VGND.n650 VGND.n649 16.0005
R3518 VGND.n2171 VGND.n650 16.0005
R3519 VGND.n634 VGND.n633 16.0005
R3520 VGND.n633 VGND.n595 16.0005
R3521 VGND.n627 VGND.n595 16.0005
R3522 VGND.n627 VGND.n626 16.0005
R3523 VGND.n626 VGND.n625 16.0005
R3524 VGND.n625 VGND.n597 16.0005
R3525 VGND.n619 VGND.n597 16.0005
R3526 VGND.n619 VGND.n618 16.0005
R3527 VGND.n617 VGND.n599 16.0005
R3528 VGND.n611 VGND.n599 16.0005
R3529 VGND.n611 VGND.n610 16.0005
R3530 VGND.n610 VGND.n609 16.0005
R3531 VGND.n609 VGND.n601 16.0005
R3532 VGND.n604 VGND.n601 16.0005
R3533 VGND.n604 VGND.n578 16.0005
R3534 VGND.n2206 VGND.n578 16.0005
R3535 VGND.n159 VGND.n117 16.0005
R3536 VGND.n165 VGND.n117 16.0005
R3537 VGND.n166 VGND.n165 16.0005
R3538 VGND.n167 VGND.n166 16.0005
R3539 VGND.n167 VGND.n115 16.0005
R3540 VGND.n173 VGND.n115 16.0005
R3541 VGND.n174 VGND.n173 16.0005
R3542 VGND.n2346 VGND.n174 16.0005
R3543 VGND.n158 VGND.n157 16.0005
R3544 VGND.n157 VGND.n119 16.0005
R3545 VGND.n151 VGND.n119 16.0005
R3546 VGND.n151 VGND.n150 16.0005
R3547 VGND.n150 VGND.n149 16.0005
R3548 VGND.n149 VGND.n121 16.0005
R3549 VGND.n143 VGND.n121 16.0005
R3550 VGND.n143 VGND.n142 16.0005
R3551 VGND.n141 VGND.n123 16.0005
R3552 VGND.n135 VGND.n123 16.0005
R3553 VGND.n135 VGND.n134 16.0005
R3554 VGND.n134 VGND.n133 16.0005
R3555 VGND.n133 VGND.n125 16.0005
R3556 VGND.n128 VGND.n125 16.0005
R3557 VGND.n128 VGND.n102 16.0005
R3558 VGND.n2381 VGND.n102 16.0005
R3559 VGND.n918 VGND.t282 16.0005
R3560 VGND.n1396 VGND.t257 15.0005
R3561 VGND.n1384 VGND.t109 15.0005
R3562 VGND.n1384 VGND.t256 15.0005
R3563 VGND.t262 VGND.n980 15.0005
R3564 VGND.n980 VGND.t42 15.0005
R3565 VGND.n981 VGND.t262 15.0005
R3566 VGND.n974 VGND.t253 15.0005
R3567 VGND.n1418 VGND.t184 15.0005
R3568 VGND.n1418 VGND.t252 15.0005
R3569 VGND.t245 VGND.n1421 15.0005
R3570 VGND.n1421 VGND.t157 15.0005
R3571 VGND.n1422 VGND.t245 15.0005
R3572 VGND.n943 VGND.t226 15.0005
R3573 VGND.n969 VGND.t194 15.0005
R3574 VGND.n969 VGND.t225 15.0005
R3575 VGND.n967 VGND.t229 15.0005
R3576 VGND.n967 VGND.t161 15.0005
R3577 VGND.t229 VGND.n966 15.0005
R3578 VGND.t53 VGND.t244 14.9665
R3579 VGND.t305 VGND.t275 14.9665
R3580 VGND.t220 VGND.t232 14.9665
R3581 VGND.n380 VGND.n364 14.555
R3582 VGND.n937 VGND.n935 14.0805
R3583 VGND.n1434 VGND.n1433 14.0805
R3584 VGND.n1404 VGND.n1403 14.0349
R3585 VGND.n1431 VGND.n1430 14.0349
R3586 VGND.n2511 VGND.n2509 13.863
R3587 VGND.n1636 VGND.n1635 12.8005
R3588 VGND.n1635 VGND.n1634 12.8005
R3589 VGND.n2456 VGND.n56 12.8005
R3590 VGND.n2453 VGND.n56 12.8005
R3591 VGND.n1619 VGND.n804 12.8005
R3592 VGND.n1623 VGND.n804 12.8005
R3593 VGND.n1410 VGND.n1409 12.8005
R3594 VGND.n995 VGND.n994 12.8005
R3595 VGND.n1368 VGND.n1338 12.7323
R3596 VGND.n2510 VGND.t331 12.051
R3597 VGND.n40 VGND.n27 11.7484
R3598 VGND.n1689 VGND.n1688 11.6369
R3599 VGND.n1691 VGND.n1689 11.6369
R3600 VGND.n1691 VGND.n1690 11.6369
R3601 VGND.n1690 VGND.n1656 11.6369
R3602 VGND.n1656 VGND.n1654 11.6369
R3603 VGND.n1699 VGND.n1654 11.6369
R3604 VGND.n1700 VGND.n1699 11.6369
R3605 VGND.n1701 VGND.n1700 11.6369
R3606 VGND.n1701 VGND.n1649 11.6369
R3607 VGND.n1708 VGND.n1649 11.6369
R3608 VGND.n1666 VGND.n745 11.6369
R3609 VGND.n1667 VGND.n1666 11.6369
R3610 VGND.n1667 VGND.n1663 11.6369
R3611 VGND.n1673 VGND.n1663 11.6369
R3612 VGND.n1674 VGND.n1673 11.6369
R3613 VGND.n1675 VGND.n1674 11.6369
R3614 VGND.n1675 VGND.n1661 11.6369
R3615 VGND.n1681 VGND.n1661 11.6369
R3616 VGND.n1682 VGND.n1681 11.6369
R3617 VGND.n1683 VGND.n1682 11.6369
R3618 VGND.n1683 VGND.n1659 11.6369
R3619 VGND.n2037 VGND.n2033 11.6369
R3620 VGND.n2042 VGND.n2037 11.6369
R3621 VGND.n2042 VGND.n2041 11.6369
R3622 VGND.n2041 VGND.n2040 11.6369
R3623 VGND.n2040 VGND.n374 11.6369
R3624 VGND.n2329 VGND.n374 11.6369
R3625 VGND.n2329 VGND.n2328 11.6369
R3626 VGND.n2328 VGND.n2327 11.6369
R3627 VGND.n2327 VGND.n375 11.6369
R3628 VGND.n2321 VGND.n375 11.6369
R3629 VGND.n2070 VGND.n2069 11.6369
R3630 VGND.n2069 VGND.n2066 11.6369
R3631 VGND.n2066 VGND.n2065 11.6369
R3632 VGND.n2065 VGND.n2062 11.6369
R3633 VGND.n2062 VGND.n2061 11.6369
R3634 VGND.n2061 VGND.n2058 11.6369
R3635 VGND.n2058 VGND.n2057 11.6369
R3636 VGND.n2057 VGND.n2054 11.6369
R3637 VGND.n2054 VGND.n2053 11.6369
R3638 VGND.n2053 VGND.n2050 11.6369
R3639 VGND.n2050 VGND.n2049 11.6369
R3640 VGND.n2014 VGND.n349 11.6369
R3641 VGND.n2017 VGND.n2014 11.6369
R3642 VGND.n2018 VGND.n2017 11.6369
R3643 VGND.n2021 VGND.n2018 11.6369
R3644 VGND.n2022 VGND.n2021 11.6369
R3645 VGND.n2025 VGND.n2022 11.6369
R3646 VGND.n2026 VGND.n2025 11.6369
R3647 VGND.n2029 VGND.n2026 11.6369
R3648 VGND.n2031 VGND.n2029 11.6369
R3649 VGND.n2032 VGND.n2031 11.6369
R3650 VGND.n2109 VGND.n2032 11.6369
R3651 VGND.n1991 VGND.n1990 11.6369
R3652 VGND.n1990 VGND.n1989 11.6369
R3653 VGND.n1989 VGND.n1987 11.6369
R3654 VGND.n1987 VGND.n1984 11.6369
R3655 VGND.n1984 VGND.n1983 11.6369
R3656 VGND.n1983 VGND.n1980 11.6369
R3657 VGND.n1980 VGND.n1979 11.6369
R3658 VGND.n1979 VGND.n1976 11.6369
R3659 VGND.n1976 VGND.n1975 11.6369
R3660 VGND.n1975 VGND.n1973 11.6369
R3661 VGND.n1121 VGND.n1120 11.6369
R3662 VGND.n1120 VGND.n1021 11.6369
R3663 VGND.n1114 VGND.n1021 11.6369
R3664 VGND.n1114 VGND.n1113 11.6369
R3665 VGND.n1113 VGND.n1112 11.6369
R3666 VGND.n1112 VGND.n1026 11.6369
R3667 VGND.n1106 VGND.n1026 11.6369
R3668 VGND.n1106 VGND.n1105 11.6369
R3669 VGND.n1105 VGND.n1104 11.6369
R3670 VGND.n1104 VGND.n1031 11.6369
R3671 VGND.n1098 VGND.n1031 11.6369
R3672 VGND.n1276 VGND.n1275 11.6369
R3673 VGND.n1275 VGND.n1274 11.6369
R3674 VGND.n1274 VGND.n1122 11.6369
R3675 VGND.n1268 VGND.n1122 11.6369
R3676 VGND.n1268 VGND.n1267 11.6369
R3677 VGND.n1267 VGND.n1266 11.6369
R3678 VGND.n1266 VGND.n1126 11.6369
R3679 VGND.n1260 VGND.n1126 11.6369
R3680 VGND.n1260 VGND.n1259 11.6369
R3681 VGND.n1259 VGND.n1258 11.6369
R3682 VGND.n2144 VGND.n2143 11.6369
R3683 VGND.n2145 VGND.n2144 11.6369
R3684 VGND.n2145 VGND.n1998 11.6369
R3685 VGND.n2151 VGND.n1998 11.6369
R3686 VGND.n2152 VGND.n2151 11.6369
R3687 VGND.n2153 VGND.n2152 11.6369
R3688 VGND.n2153 VGND.n1996 11.6369
R3689 VGND.n2159 VGND.n1996 11.6369
R3690 VGND.n2160 VGND.n2159 11.6369
R3691 VGND.n2161 VGND.n2160 11.6369
R3692 VGND.n2137 VGND.n2000 11.6369
R3693 VGND.n2137 VGND.n2136 11.6369
R3694 VGND.n2136 VGND.n2135 11.6369
R3695 VGND.n2135 VGND.n2114 11.6369
R3696 VGND.n2130 VGND.n2114 11.6369
R3697 VGND.n2130 VGND.n2129 11.6369
R3698 VGND.n2129 VGND.n2128 11.6369
R3699 VGND.n2128 VGND.n2117 11.6369
R3700 VGND.n2123 VGND.n2117 11.6369
R3701 VGND.n2123 VGND.n2122 11.6369
R3702 VGND.n2122 VGND.n350 11.6369
R3703 VGND.n1834 VGND.n1833 11.6369
R3704 VGND.n1833 VGND.n739 11.6369
R3705 VGND.n1828 VGND.n739 11.6369
R3706 VGND.n1828 VGND.n1827 11.6369
R3707 VGND.n1827 VGND.n1826 11.6369
R3708 VGND.n1826 VGND.n741 11.6369
R3709 VGND.n1820 VGND.n741 11.6369
R3710 VGND.n1820 VGND.n1819 11.6369
R3711 VGND.n1819 VGND.n1818 11.6369
R3712 VGND.n1818 VGND.n743 11.6369
R3713 VGND.n1812 VGND.n743 11.6369
R3714 VGND.n714 VGND.n660 11.6369
R3715 VGND.n719 VGND.n714 11.6369
R3716 VGND.n720 VGND.n719 11.6369
R3717 VGND.n721 VGND.n720 11.6369
R3718 VGND.n721 VGND.n712 11.6369
R3719 VGND.n727 VGND.n712 11.6369
R3720 VGND.n728 VGND.n727 11.6369
R3721 VGND.n729 VGND.n728 11.6369
R3722 VGND.n729 VGND.n710 11.6369
R3723 VGND.n735 VGND.n710 11.6369
R3724 VGND.n736 VGND.n735 11.6369
R3725 VGND.n2411 VGND.n2410 11.6369
R3726 VGND.n2410 VGND.n2409 11.6369
R3727 VGND.n2409 VGND.n86 11.6369
R3728 VGND.n2403 VGND.n86 11.6369
R3729 VGND.n2403 VGND.n2402 11.6369
R3730 VGND.n2402 VGND.n2401 11.6369
R3731 VGND.n2401 VGND.n91 11.6369
R3732 VGND.n2395 VGND.n91 11.6369
R3733 VGND.n2395 VGND.n2394 11.6369
R3734 VGND.n2394 VGND.n2393 11.6369
R3735 VGND.n2436 VGND.n2435 11.6369
R3736 VGND.n2435 VGND.n2434 11.6369
R3737 VGND.n2434 VGND.n73 11.6369
R3738 VGND.n2428 VGND.n73 11.6369
R3739 VGND.n2428 VGND.n2427 11.6369
R3740 VGND.n2427 VGND.n2426 11.6369
R3741 VGND.n2426 VGND.n77 11.6369
R3742 VGND.n2420 VGND.n77 11.6369
R3743 VGND.n2420 VGND.n2419 11.6369
R3744 VGND.n2419 VGND.n2418 11.6369
R3745 VGND.n2418 VGND.n81 11.6369
R3746 VGND.n1096 VGND.n1035 11.6369
R3747 VGND.n1090 VGND.n1035 11.6369
R3748 VGND.n1090 VGND.n1089 11.6369
R3749 VGND.n1089 VGND.n1088 11.6369
R3750 VGND.n1088 VGND.n60 11.6369
R3751 VGND.n2451 VGND.n61 11.6369
R3752 VGND.n66 VGND.n61 11.6369
R3753 VGND.n2444 VGND.n66 11.6369
R3754 VGND.n2444 VGND.n2443 11.6369
R3755 VGND.n2443 VGND.n2442 11.6369
R3756 VGND.n37 VGND.n36 11.563
R3757 VGND.n33 VGND.n31 11.563
R3758 VGND.n1004 VGND.n1002 11.563
R3759 VGND.n1005 VGND.n1003 11.563
R3760 VGND.n2510 VGND.t330 11.4829
R3761 VGND.n2496 VGND.n2495 11.3369
R3762 VGND.n2512 VGND.n2511 11.1724
R3763 VGND.n1287 VGND.n1286 10.8829
R3764 VGND.n1291 VGND.n1290 10.8829
R3765 VGND.n1966 VGND.t81 10.1221
R3766 VGND.t124 VGND.n1894 10.1221
R3767 VGND.n1896 VGND.t16 10.1221
R3768 VGND.n1876 VGND.t208 10.1221
R3769 VGND.n906 VGND.n902 10.0862
R3770 VGND.n895 VGND.n891 10.0862
R3771 VGND.n919 VGND.n915 10.0862
R3772 VGND.n1334 VGND.n1333 10.0317
R3773 VGND.n1413 VGND.n977 9.97782
R3774 VGND.t261 VGND.t166 9.97782
R3775 VGND.t312 VGND.t41 9.97782
R3776 VGND.n1305 VGND.t281 9.6005
R3777 VGND.n1298 VGND.t179 9.6005
R3778 VGND.n1317 VGND.t284 9.6005
R3779 VGND.n1320 VGND.t176 9.6005
R3780 VGND.n1636 VGND.n796 9.36264
R3781 VGND.n2453 VGND.n54 9.36264
R3782 VGND.n1619 VGND.n802 9.36264
R3783 VGND.n902 VGND.n901 9.3005
R3784 VGND.n904 VGND.n903 9.3005
R3785 VGND.n891 VGND.n890 9.3005
R3786 VGND.n893 VGND.n892 9.3005
R3787 VGND.n1392 VGND.n1389 9.3005
R3788 VGND.n1397 VGND.n1388 9.3005
R3789 VGND.n1635 VGND.n797 9.3005
R3790 VGND.n1634 VGND.n1633 9.3005
R3791 VGND.n2483 VGND.n2482 9.3005
R3792 VGND.n2470 VGND.n2469 9.3005
R3793 VGND.n52 VGND.n51 9.3005
R3794 VGND.n39 VGND.n38 9.3005
R3795 VGND.n56 VGND.n55 9.3005
R3796 VGND.n2457 VGND.n2456 9.3005
R3797 VGND.n804 VGND.n803 9.3005
R3798 VGND.n1624 VGND.n1623 9.3005
R3799 VGND.n958 VGND.n957 9.3005
R3800 VGND.n965 VGND.n956 9.3005
R3801 VGND.n915 VGND.n914 9.3005
R3802 VGND.n917 VGND.n916 9.3005
R3803 VGND.n922 VGND.n889 9.3005
R3804 VGND.n912 VGND.n911 9.3005
R3805 VGND.n910 VGND.n909 9.3005
R3806 VGND.n925 VGND.n924 9.3005
R3807 VGND.n2492 VGND.n2486 9.2505
R3808 VGND.n2488 VGND.n2485 9.2505
R3809 VGND.n24 VGND.n18 9.2505
R3810 VGND.n20 VGND.n17 9.2505
R3811 VGND.t218 VGND.t45 8.67615
R3812 VGND.n457 VGND.n364 8.60107
R3813 VGND.n2511 VGND.n2510 7.60845
R3814 VGND.n842 VGND.n841 7.52932
R3815 VGND.n2537 VGND.n1 7.41931
R3816 VGND.n2481 VGND.n2480 7.4005
R3817 VGND.n2477 VGND.n2476 7.4005
R3818 VGND.n1397 VGND.n1389 7.11161
R3819 VGND.n965 VGND.n957 7.11161
R3820 VGND.n2109 VGND.n2108 6.72373
R3821 VGND.n1098 VGND.n1097 6.72373
R3822 VGND.n2336 VGND.n350 6.72373
R3823 VGND.n1812 VGND.n1811 6.72373
R3824 VGND.n737 VGND.n736 6.72373
R3825 VGND.n2442 VGND.n67 6.72373
R3826 VGND.n2478 VGND.n2477 6.30719
R3827 VGND.n2480 VGND.n2479 6.30719
R3828 VGND.n1811 VGND.n745 6.20656
R3829 VGND.n2108 VGND.n2070 6.20656
R3830 VGND.n2336 VGND.n349 6.20656
R3831 VGND.n1834 VGND.n737 6.20656
R3832 VGND.n2436 VGND.n67 6.20656
R3833 VGND.n1097 VGND.n1096 6.20656
R3834 VGND.n2452 VGND.n60 6.07727
R3835 VGND.n2413 VGND.n84 5.89178
R3836 VGND.n924 VGND.n923 5.84425
R3837 VGND.n1331 VGND.n1318 5.81868
R3838 VGND.n1327 VGND.n1318 5.81868
R3839 VGND.n862 VGND.n861 5.68939
R3840 VGND.n861 VGND.n860 5.68939
R3841 VGND.n1353 VGND.n1346 5.68939
R3842 VGND.n1338 VGND.n1337 5.66539
R3843 VGND.n2465 VGND.n2460 5.60656
R3844 VGND.n2461 VGND.n2459 5.60656
R3845 VGND.n50 VGND.n49 5.60656
R3846 VGND.n46 VGND.n45 5.60656
R3847 VGND.n2452 VGND.n2451 5.5601
R3848 VGND.n1548 VGND.n837 5.51161
R3849 VGND.n2258 VGND.n2257 5.51161
R3850 VGND.n1727 VGND.n1644 5.51161
R3851 VGND.n285 VGND.n249 5.51161
R3852 VGND.n2313 VGND.n2312 5.51161
R3853 VGND.n1904 VGND.n684 5.51161
R3854 VGND.n1183 VGND.n1156 5.51161
R3855 VGND.n2207 VGND.n2206 5.51161
R3856 VGND.n2382 VGND.n2381 5.51161
R3857 VGND.n1710 VGND.n1709 5.1717
R3858 VGND.n2320 VGND.n379 5.1717
R3859 VGND.n98 VGND.n95 5.1717
R3860 VGND.n2505 VGND.n2502 5.13939
R3861 VGND.n2509 VGND.n2501 5.13939
R3862 VGND.n909 VGND.n1 5.07862
R3863 VGND.n913 VGND.n912 5.07862
R3864 VGND.n923 VGND.n922 5.07862
R3865 VGND.t160 VGND.t66 4.98916
R3866 VGND.t264 VGND.t170 4.98916
R3867 VGND.t267 VGND.t312 4.98916
R3868 VGND.n1401 VGND.n989 4.98916
R3869 VGND.n968 VGND.n953 4.98488
R3870 VGND.n1353 VGND.n1352 4.97828
R3871 VGND.n1972 VGND.n662 4.9157
R3872 VGND.n1252 VGND.n1251 4.9157
R3873 VGND.n2168 VGND.n651 4.9157
R3874 VGND.n2466 VGND.n2465 4.90189
R3875 VGND.n2463 VGND.n2461 4.90189
R3876 VGND.n47 VGND.n46 4.90189
R3877 VGND.n49 VGND.n48 4.90189
R3878 VGND.n1417 VGND.n1416 4.78398
R3879 VGND.n971 VGND.n942 4.78398
R3880 VGND.n1387 VGND.n1386 4.64112
R3881 VGND.n2458 VGND.n2457 4.5005
R3882 VGND.n1625 VGND.n1624 4.5005
R3883 VGND.n1633 VGND.n1632 4.5005
R3884 VGND.n801 VGND.n799 4.5005
R3885 VGND.n1316 VGND.n1294 4.5005
R3886 VGND.n1313 VGND.n800 4.5005
R3887 VGND.n1316 VGND.n800 4.5005
R3888 VGND.n2531 VGND.n8 4.48804
R3889 VGND.n2527 VGND.n11 4.48804
R3890 VGND.n2483 VGND.t32 4.34657
R3891 VGND.n1782 VGND.t324 4.33832
R3892 VGND.n1795 VGND.t190 4.33832
R3893 VGND.t195 VGND.n1793 4.33832
R3894 VGND.n1718 VGND.t142 4.33832
R3895 VGND.n2535 VGND.n5 4.32167
R3896 VGND.n1838 VGND.n708 4.26717
R3897 VGND.n1844 VGND.n708 4.26717
R3898 VGND.n1844 VGND.n706 4.26717
R3899 VGND.n1850 VGND.n706 4.26717
R3900 VGND.n1850 VGND.n704 4.26717
R3901 VGND.n1856 VGND.n704 4.26717
R3902 VGND.n1856 VGND.n702 4.26717
R3903 VGND.n1862 VGND.n702 4.26717
R3904 VGND.n1862 VGND.n700 4.26717
R3905 VGND.n1868 VGND.n700 4.26717
R3906 VGND.n1868 VGND.n697 4.26717
R3907 VGND.n2335 VGND.n352 4.26717
R3908 VGND.n549 VGND.n352 4.26717
R3909 VGND.n549 VGND.n545 4.26717
R3910 VGND.n557 VGND.n545 4.26717
R3911 VGND.n558 VGND.n557 4.26717
R3912 VGND.n561 VGND.n558 4.26717
R3913 VGND.n561 VGND.n543 4.26717
R3914 VGND.n568 VGND.n543 4.26717
R3915 VGND.n571 VGND.n568 4.26717
R3916 VGND.n571 VGND.n541 4.26717
R3917 VGND.n2214 VGND.n541 4.26717
R3918 VGND.n1042 VGND.n1034 4.26717
R3919 VGND.n1077 VGND.n1042 4.26717
R3920 VGND.n1077 VGND.n1076 4.26717
R3921 VGND.n1076 VGND.n1075 4.26717
R3922 VGND.n1075 VGND.n1073 4.26717
R3923 VGND.n1073 VGND.n1070 4.26717
R3924 VGND.n1070 VGND.n1069 4.26717
R3925 VGND.n1069 VGND.n1066 4.26717
R3926 VGND.n1066 VGND.n1065 4.26717
R3927 VGND.n1065 VGND.n1062 4.26717
R3928 VGND.n1062 VGND.n1061 4.26717
R3929 VGND.n195 VGND.n193 4.26717
R3930 VGND.n195 VGND.n190 4.26717
R3931 VGND.n201 VGND.n190 4.26717
R3932 VGND.n202 VGND.n201 4.26717
R3933 VGND.n202 VGND.n186 4.26717
R3934 VGND.n209 VGND.n186 4.26717
R3935 VGND.n210 VGND.n209 4.26717
R3936 VGND.n210 VGND.n182 4.26717
R3937 VGND.n216 VGND.n182 4.26717
R3938 VGND.n217 VGND.n216 4.26717
R3939 VGND.n217 VGND.n179 4.26717
R3940 VGND.n2107 VGND.n2071 4.26717
R3941 VGND.n2102 VGND.n2071 4.26717
R3942 VGND.n2102 VGND.n2101 4.26717
R3943 VGND.n2101 VGND.n2079 4.26717
R3944 VGND.n2096 VGND.n2079 4.26717
R3945 VGND.n2096 VGND.n2095 4.26717
R3946 VGND.n2095 VGND.n2094 4.26717
R3947 VGND.n2094 VGND.n2089 4.26717
R3948 VGND.n2089 VGND.n461 4.26717
R3949 VGND.n2267 VGND.n461 4.26717
R3950 VGND.n2267 VGND.n459 4.26717
R3951 VGND.n1810 VGND.n746 4.26717
R3952 VGND.n1504 VGND.n746 4.26717
R3953 VGND.n1505 VGND.n1504 4.26717
R3954 VGND.n1510 VGND.n1505 4.26717
R3955 VGND.n1511 VGND.n1510 4.26717
R3956 VGND.n1516 VGND.n1511 4.26717
R3957 VGND.n1517 VGND.n1516 4.26717
R3958 VGND.n1522 VGND.n1517 4.26717
R3959 VGND.n1523 VGND.n1522 4.26717
R3960 VGND.n1526 VGND.n1523 4.26717
R3961 VGND.n1526 VGND.n790 4.26717
R3962 VGND.n2470 VGND.t38 4.22295
R3963 VGND.n52 VGND.t101 4.22295
R3964 VGND.n1838 VGND.n737 3.93531
R3965 VGND.n2336 VGND.n2335 3.93531
R3966 VGND.n1097 VGND.n1034 3.93531
R3967 VGND.n193 VGND.n67 3.93531
R3968 VGND.n2108 VGND.n2107 3.93531
R3969 VGND.n1811 VGND.n1810 3.93531
R3970 VGND.n1616 VGND.n1615 3.7893
R3971 VGND.n1612 VGND.n811 3.7893
R3972 VGND.n1611 VGND.n814 3.7893
R3973 VGND.n818 VGND.n817 3.7893
R3974 VGND.n1605 VGND.n1604 3.7893
R3975 VGND.n1531 VGND.n819 3.7893
R3976 VGND.n1537 VGND.n1536 3.7893
R3977 VGND.n1533 VGND.n1532 3.7893
R3978 VGND.n1545 VGND.n838 3.7893
R3979 VGND.n2220 VGND.n477 3.7893
R3980 VGND.n2229 VGND.n2228 3.7893
R3981 VGND.n475 VGND.n474 3.7893
R3982 VGND.n2237 VGND.n2235 3.7893
R3983 VGND.n2236 VGND.n472 3.7893
R3984 VGND.n2244 VGND.n2243 3.7893
R3985 VGND.n470 VGND.n469 3.7893
R3986 VGND.n2252 VGND.n2250 3.7893
R3987 VGND.n2251 VGND.n465 3.7893
R3988 VGND.n1798 VGND.n780 3.7893
R3989 VGND.n1797 VGND.n781 3.7893
R3990 VGND.n1786 VGND.n1785 3.7893
R3991 VGND.n1791 VGND.n1790 3.7893
R3992 VGND.n1787 VGND.n758 3.7893
R3993 VGND.n1804 VGND.n1803 3.7893
R3994 VGND.n1713 VGND.n759 3.7893
R3995 VGND.n1716 VGND.n1715 3.7893
R3996 VGND.n1724 VGND.n1645 3.7893
R3997 VGND.n345 VGND.n228 3.7893
R3998 VGND.n341 VGND.n340 3.7893
R3999 VGND.n258 VGND.n230 3.7893
R4000 VGND.n259 VGND.n254 3.7893
R4001 VGND.n264 VGND.n263 3.7893
R4002 VGND.n267 VGND.n252 3.7893
R4003 VGND.n269 VGND.n268 3.7893
R4004 VGND.n273 VGND.n272 3.7893
R4005 VGND.n282 VGND.n250 3.7893
R4006 VGND.n2275 VGND.n394 3.7893
R4007 VGND.n2284 VGND.n2283 3.7893
R4008 VGND.n392 VGND.n391 3.7893
R4009 VGND.n2292 VGND.n2290 3.7893
R4010 VGND.n2291 VGND.n389 3.7893
R4011 VGND.n2299 VGND.n2298 3.7893
R4012 VGND.n387 VGND.n386 3.7893
R4013 VGND.n2307 VGND.n2305 3.7893
R4014 VGND.n2306 VGND.n382 3.7893
R4015 VGND.n1958 VGND.n664 3.7893
R4016 VGND.n1957 VGND.n667 3.7893
R4017 VGND.n1964 VGND.n1963 3.7893
R4018 VGND.n1882 VGND.n668 3.7893
R4019 VGND.n1885 VGND.n1884 3.7893
R4020 VGND.n1890 VGND.n1881 3.7893
R4021 VGND.n1892 VGND.n1891 3.7893
R4022 VGND.n1899 VGND.n688 3.7893
R4023 VGND.n1898 VGND.n686 3.7893
R4024 VGND.n1247 VGND.n1246 3.7893
R4025 VGND.n1243 VGND.n1132 3.7893
R4026 VGND.n1242 VGND.n1135 3.7893
R4027 VGND.n1238 VGND.n1237 3.7893
R4028 VGND.n1159 VGND.n1137 3.7893
R4029 VGND.n1165 VGND.n1163 3.7893
R4030 VGND.n1167 VGND.n1166 3.7893
R4031 VGND.n1171 VGND.n1170 3.7893
R4032 VGND.n1180 VGND.n1157 3.7893
R4033 VGND.n2169 VGND.n589 3.7893
R4034 VGND.n2178 VGND.n2177 3.7893
R4035 VGND.n587 VGND.n586 3.7893
R4036 VGND.n2186 VGND.n2184 3.7893
R4037 VGND.n2185 VGND.n584 3.7893
R4038 VGND.n2193 VGND.n2192 3.7893
R4039 VGND.n582 VGND.n581 3.7893
R4040 VGND.n2201 VGND.n2199 3.7893
R4041 VGND.n2200 VGND.n577 3.7893
R4042 VGND.n2344 VGND.n113 3.7893
R4043 VGND.n2353 VGND.n2352 3.7893
R4044 VGND.n111 VGND.n110 3.7893
R4045 VGND.n2361 VGND.n2359 3.7893
R4046 VGND.n2360 VGND.n108 3.7893
R4047 VGND.n2368 VGND.n2367 3.7893
R4048 VGND.n106 VGND.n105 3.7893
R4049 VGND.n2376 VGND.n2374 3.7893
R4050 VGND.n2375 VGND.n101 3.7893
R4051 VGND.t283 VGND.n0 1.95574
R4052 VGND.n1393 VGND.n1392 3.55702
R4053 VGND.n959 VGND.n958 3.55702
R4054 VGND.n2503 VGND.n2501 3.52815
R4055 VGND.n2506 VGND.n2505 3.52815
R4056 VGND.n1390 VGND.n1389 3.48951
R4057 VGND.n1391 VGND.n1390 3.48951
R4058 VGND.n957 VGND.n954 3.48951
R4059 VGND.n960 VGND.n954 3.48951
R4060 VGND.n2535 VGND.n2533 3.4105
R4061 VGND.n2536 VGND.n2535 3.4105
R4062 VGND.n2531 VGND.n2529 3.4105
R4063 VGND.n2532 VGND.n2531 3.4105
R4064 VGND.n2527 VGND.n2525 3.4105
R4065 VGND.n2528 VGND.n2527 3.4105
R4066 VGND.n2523 VGND.n2521 3.4105
R4067 VGND.n2524 VGND.n2523 3.4105
R4068 VGND.n2519 VGND.n2517 3.4105
R4069 VGND.n2520 VGND.n2519 3.4105
R4070 VGND.n2514 VGND.n2512 3.4105
R4071 VGND.n2516 VGND.n2515 3.4105
R4072 VGND.n2514 VGND.n2513 3.4105
R4073 VGND.n2515 VGND.n2514 3.4105
R4074 VGND.n2523 VGND.n14 3.39037
R4075 VGND.n1404 VGND.n1014 3.16744
R4076 VGND.n1386 VGND.n14 3.16281
R4077 VGND.n985 VGND.n979 3.14514
R4078 VGND.n950 VGND.n946 3.14514
R4079 VGND.n986 VGND.n985 3.1005
R4080 VGND.n983 VGND.n973 3.1005
R4081 VGND.n1416 VGND.n1415 3.1005
R4082 VGND.n951 VGND.n950 3.1005
R4083 VGND.n949 VGND.n944 3.1005
R4084 VGND.n1424 VGND.n942 3.1005
R4085 VGND.n1309 VGND.n1297 2.86505
R4086 VGND.n1309 VGND.n1308 2.86505
R4087 VGND.n1306 VGND.n1300 2.86505
R4088 VGND.n1301 VGND.n1300 2.86505
R4089 VGND.n1308 VGND.n1307 2.86505
R4090 VGND.n1304 VGND.n1301 2.86505
R4091 VGND.n1312 VGND.n1297 2.86505
R4092 VGND.n1307 VGND.n1306 2.86505
R4093 VGND.n1326 VGND.n1325 2.86505
R4094 VGND.n1325 VGND.n1324 2.86505
R4095 VGND.n1324 VGND.n1323 2.86505
R4096 VGND.n1327 VGND.n1326 2.86505
R4097 VGND.n1333 VGND.n1332 2.8366
R4098 VGND.n810 VGND.n809 2.6629
R4099 VGND.n1643 VGND.n788 2.6629
R4100 VGND.n2221 VGND.n2219 2.6629
R4101 VGND.n463 VGND.n456 2.6629
R4102 VGND.n1780 VGND.n1779 2.6629
R4103 VGND.n347 VGND.n346 2.6629
R4104 VGND.n277 VGND.n175 2.6629
R4105 VGND.n2276 VGND.n2274 2.6629
R4106 VGND.n1953 VGND.n662 2.6629
R4107 VGND.n694 VGND.n693 2.6629
R4108 VGND.n1251 VGND.n1130 2.6629
R4109 VGND.n1175 VGND.n348 2.6629
R4110 VGND.n2170 VGND.n2168 2.6629
R4111 VGND.n575 VGND.n539 2.6629
R4112 VGND.n2345 VGND.n2343 2.6629
R4113 VGND.n1395 VGND.n1393 2.60059
R4114 VGND.n959 VGND.n955 2.60059
R4115 VGND.n1393 VGND.n1391 2.55763
R4116 VGND.n960 VGND.n959 2.55763
R4117 VGND.n809 VGND.n694 2.4581
R4118 VGND.n837 VGND.n788 2.4581
R4119 VGND.n2219 VGND.n539 2.4581
R4120 VGND.n2258 VGND.n463 2.4581
R4121 VGND.n1780 VGND.n1643 2.4581
R4122 VGND.n1710 VGND.n1644 2.4581
R4123 VGND.n348 VGND.n347 2.4581
R4124 VGND.n277 VGND.n249 2.4581
R4125 VGND.n2274 VGND.n456 2.4581
R4126 VGND.n2313 VGND.n379 2.4581
R4127 VGND.n693 VGND.n684 2.4581
R4128 VGND.n1175 VGND.n1156 2.4581
R4129 VGND.n2207 VGND.n575 2.4581
R4130 VGND.n2343 VGND.n175 2.4581
R4131 VGND.n2382 VGND.n98 2.4581
R4132 VGND.n1335 VGND.n1334 2.44675
R4133 VGND.n1334 VGND.n1281 2.44675
R4134 VGND.n1009 VGND.t19 2.37317
R4135 VGND.t19 VGND.n1008 2.37317
R4136 VGND.n35 VGND.t287 2.2941
R4137 VGND.n32 VGND.t287 2.2941
R4138 VGND.n2519 VGND.n2496 2.27233
R4139 VGND.n1626 VGND.n798 2.26187
R4140 VGND.n1315 VGND.n1314 2.26187
R4141 VGND.n983 VGND.n975 2.25882
R4142 VGND.n984 VGND.n983 2.25882
R4143 VGND.n982 VGND.n979 2.25882
R4144 VGND.n986 VGND.n984 2.25882
R4145 VGND.n1415 VGND.n975 2.25882
R4146 VGND.n986 VGND.n982 2.25882
R4147 VGND.n1423 VGND.n944 2.25882
R4148 VGND.n948 VGND.n944 2.25882
R4149 VGND.n952 VGND.n946 2.25882
R4150 VGND.n951 VGND.n948 2.25882
R4151 VGND.n1424 VGND.n1423 2.25882
R4152 VGND.n952 VGND.n951 2.25882
R4153 VGND.n1627 VGND.n1626 2.24063
R4154 VGND.n1314 VGND.n1313 2.24063
R4155 VGND.n1296 VGND.n1295 2.24063
R4156 VGND.n1629 VGND.n1628 2.24063
R4157 VGND.n1631 VGND.n1630 2.24063
R4158 VGND.n2458 VGND.n54 2.22018
R4159 VGND.n1625 VGND.n802 2.22018
R4160 VGND.n1632 VGND.n796 2.22018
R4161 VGND.n1288 VGND.t185 2.20954
R4162 VGND.t185 VGND.n1284 2.20954
R4163 VGND.n697 VGND.n694 2.18124
R4164 VGND.n2214 VGND.n539 2.18124
R4165 VGND.n1061 VGND.n348 2.18124
R4166 VGND.n179 VGND.n175 2.18124
R4167 VGND.n459 VGND.n456 2.18124
R4168 VGND.n1643 VGND.n790 2.18124
R4169 VGND.n1544 VGND.n837 2.1509
R4170 VGND.n2259 VGND.n2258 2.1509
R4171 VGND.n1723 VGND.n1644 2.1509
R4172 VGND.n281 VGND.n249 2.1509
R4173 VGND.n2314 VGND.n2313 2.1509
R4174 VGND.n691 VGND.n684 2.1509
R4175 VGND.n1179 VGND.n1156 2.1509
R4176 VGND.n2208 VGND.n2207 2.1509
R4177 VGND.n2383 VGND.n2382 2.1509
R4178 VGND.n1584 VGND.n810 2.13383
R4179 VGND.n2222 VGND.n2221 2.13383
R4180 VGND.n1779 VGND.n1778 2.13383
R4181 VGND.n346 VGND.n227 2.13383
R4182 VGND.n2277 VGND.n2276 2.13383
R4183 VGND.n1954 VGND.n1953 2.13383
R4184 VGND.n1219 VGND.n1130 2.13383
R4185 VGND.n2171 VGND.n2170 2.13383
R4186 VGND.n2346 VGND.n2345 2.13383
R4187 VGND.n1873 VGND.n694 2.08643
R4188 VGND.n540 VGND.n539 2.08643
R4189 VGND.n2337 VGND.n348 2.08643
R4190 VGND.n177 VGND.n175 2.08643
R4191 VGND.n458 VGND.n456 2.08643
R4192 VGND.n1643 VGND.n1642 2.08643
R4193 VGND.n2484 VGND.n2483 2.03694
R4194 VGND.n2471 VGND.n2470 2.03694
R4195 VGND.n53 VGND.n52 2.03694
R4196 VGND.n40 VGND.n39 2.03694
R4197 VGND.n1616 VGND.n810 1.9461
R4198 VGND.n2221 VGND.n2220 1.9461
R4199 VGND.n1779 VGND.n780 1.9461
R4200 VGND.n346 VGND.n345 1.9461
R4201 VGND.n2276 VGND.n2275 1.9461
R4202 VGND.n1953 VGND.n664 1.9461
R4203 VGND.n1247 VGND.n1130 1.9461
R4204 VGND.n2170 VGND.n2169 1.9461
R4205 VGND.n2345 VGND.n2344 1.9461
R4206 VGND.n1994 VGND.n0 3.39918
R4207 VGND.n2491 VGND.t155 1.78135
R4208 VGND.t155 VGND.n2487 1.78135
R4209 VGND.n23 VGND.t18 1.78135
R4210 VGND.t18 VGND.n19 1.78135
R4211 VGND.n2533 VGND.n3 1.70675
R4212 VGND.n2529 VGND.n7 1.70675
R4213 VGND.n2517 VGND.n16 1.70675
R4214 VGND.n2525 VGND.n10 1.70675
R4215 VGND.n2521 VGND.n13 1.70675
R4216 VGND.n2536 VGND.n3 1.706
R4217 VGND.n2532 VGND.n7 1.706
R4218 VGND.n2528 VGND.n10 1.706
R4219 VGND.n2524 VGND.n13 1.706
R4220 VGND.n2520 VGND.n16 1.706
R4221 VGND.n2534 VGND.n2 1.70307
R4222 VGND.n2530 VGND.n6 1.70307
R4223 VGND.n2526 VGND.n9 1.70307
R4224 VGND.n2522 VGND.n12 1.70307
R4225 VGND.n2518 VGND.n15 1.70307
R4226 VGND.n2499 VGND.n2497 1.70248
R4227 VGND.n2516 VGND.n2498 1.70149
R4228 VGND.n2506 VGND.t46 1.60927
R4229 VGND.n2503 VGND.t46 1.60927
R4230 VGND.n1709 VGND.n1708 1.47392
R4231 VGND.n2321 VGND.n2320 1.47392
R4232 VGND.n1973 VGND.n1972 1.47392
R4233 VGND.n1258 VGND.n1252 1.47392
R4234 VGND.n2161 VGND.n651 1.47392
R4235 VGND.n2393 VGND.n95 1.47392
R4236 VGND.n2471 VGND.n2458 1.33383
R4237 VGND.t323 VGND.t10 1.31787
R4238 VGND.t180 VGND.t6 1.31787
R4239 VGND.t47 VGND.t94 1.31787
R4240 VGND.n2458 VGND.n53 1.26612
R4241 VGND.n2521 VGND.n2520 1.20488
R4242 VGND.n2479 VGND.t31 1.08466
R4243 VGND.t31 VGND.n2478 1.08466
R4244 VGND.n1485 VGND.n1483 1.063
R4245 VGND.n841 VGND.n84 1.03743
R4246 VGND.n1468 VGND.n848 1.03175
R4247 VGND.n1463 VGND.n1461 0.891125
R4248 VGND.n1449 VGND.n1447 0.859875
R4249 VGND.n1457 VGND.n1455 0.859875
R4250 VGND.n1615 VGND.n811 0.8197
R4251 VGND.n1612 VGND.n1611 0.8197
R4252 VGND.n817 VGND.n814 0.8197
R4253 VGND.n1605 VGND.n818 0.8197
R4254 VGND.n1604 VGND.n819 0.8197
R4255 VGND.n1537 VGND.n1531 0.8197
R4256 VGND.n1536 VGND.n1532 0.8197
R4257 VGND.n1533 VGND.n838 0.8197
R4258 VGND.n1545 VGND.n1544 0.8197
R4259 VGND.n2229 VGND.n477 0.8197
R4260 VGND.n2228 VGND.n475 0.8197
R4261 VGND.n2235 VGND.n474 0.8197
R4262 VGND.n2237 VGND.n2236 0.8197
R4263 VGND.n2244 VGND.n472 0.8197
R4264 VGND.n2243 VGND.n470 0.8197
R4265 VGND.n2250 VGND.n469 0.8197
R4266 VGND.n2252 VGND.n2251 0.8197
R4267 VGND.n2259 VGND.n465 0.8197
R4268 VGND.n1798 VGND.n1797 0.8197
R4269 VGND.n1785 VGND.n781 0.8197
R4270 VGND.n1791 VGND.n1786 0.8197
R4271 VGND.n1790 VGND.n1787 0.8197
R4272 VGND.n1804 VGND.n758 0.8197
R4273 VGND.n1803 VGND.n759 0.8197
R4274 VGND.n1716 VGND.n1713 0.8197
R4275 VGND.n1715 VGND.n1645 0.8197
R4276 VGND.n1724 VGND.n1723 0.8197
R4277 VGND.n341 VGND.n228 0.8197
R4278 VGND.n340 VGND.n230 0.8197
R4279 VGND.n259 VGND.n258 0.8197
R4280 VGND.n263 VGND.n254 0.8197
R4281 VGND.n264 VGND.n252 0.8197
R4282 VGND.n268 VGND.n267 0.8197
R4283 VGND.n273 VGND.n269 0.8197
R4284 VGND.n272 VGND.n250 0.8197
R4285 VGND.n282 VGND.n281 0.8197
R4286 VGND.n2284 VGND.n394 0.8197
R4287 VGND.n2283 VGND.n392 0.8197
R4288 VGND.n2290 VGND.n391 0.8197
R4289 VGND.n2292 VGND.n2291 0.8197
R4290 VGND.n2299 VGND.n389 0.8197
R4291 VGND.n2298 VGND.n387 0.8197
R4292 VGND.n2305 VGND.n386 0.8197
R4293 VGND.n2307 VGND.n2306 0.8197
R4294 VGND.n2314 VGND.n382 0.8197
R4295 VGND.n1958 VGND.n1957 0.8197
R4296 VGND.n1964 VGND.n667 0.8197
R4297 VGND.n1963 VGND.n668 0.8197
R4298 VGND.n1884 VGND.n1882 0.8197
R4299 VGND.n1885 VGND.n1881 0.8197
R4300 VGND.n1892 VGND.n1890 0.8197
R4301 VGND.n1891 VGND.n688 0.8197
R4302 VGND.n1899 VGND.n1898 0.8197
R4303 VGND.n691 VGND.n686 0.8197
R4304 VGND.n1246 VGND.n1132 0.8197
R4305 VGND.n1243 VGND.n1242 0.8197
R4306 VGND.n1238 VGND.n1135 0.8197
R4307 VGND.n1237 VGND.n1137 0.8197
R4308 VGND.n1163 VGND.n1159 0.8197
R4309 VGND.n1166 VGND.n1165 0.8197
R4310 VGND.n1171 VGND.n1167 0.8197
R4311 VGND.n1170 VGND.n1157 0.8197
R4312 VGND.n1180 VGND.n1179 0.8197
R4313 VGND.n2178 VGND.n589 0.8197
R4314 VGND.n2177 VGND.n587 0.8197
R4315 VGND.n2184 VGND.n586 0.8197
R4316 VGND.n2186 VGND.n2185 0.8197
R4317 VGND.n2193 VGND.n584 0.8197
R4318 VGND.n2192 VGND.n582 0.8197
R4319 VGND.n2199 VGND.n581 0.8197
R4320 VGND.n2201 VGND.n2200 0.8197
R4321 VGND.n2208 VGND.n577 0.8197
R4322 VGND.n2353 VGND.n113 0.8197
R4323 VGND.n2352 VGND.n111 0.8197
R4324 VGND.n2359 VGND.n110 0.8197
R4325 VGND.n2361 VGND.n2360 0.8197
R4326 VGND.n2368 VGND.n108 0.8197
R4327 VGND.n2367 VGND.n106 0.8197
R4328 VGND.n2374 VGND.n105 0.8197
R4329 VGND.n2376 VGND.n2375 0.8197
R4330 VGND.n2383 VGND.n101 0.8197
R4331 VGND.n1372 VGND.n1017 0.813
R4332 VGND.n923 VGND.n913 0.813
R4333 VGND.n913 VGND.n1 0.813
R4334 VGND.n908 VGND.n907 0.788301
R4335 VGND.n897 VGND.n896 0.788301
R4336 VGND.n921 VGND.n920 0.788301
R4337 VGND.n2484 VGND.n2471 0.7505
R4338 VGND.n1488 VGND.n1487 0.734875
R4339 VGND.n1477 VGND.n1476 0.734875
R4340 VGND.n1488 VGND.n1474 0.71925
R4341 VGND.n2466 VGND.t37 0.701195
R4342 VGND.n2463 VGND.t37 0.701195
R4343 VGND.n48 VGND.t100 0.701195
R4344 VGND.t100 VGND.n47 0.701195
R4345 VGND.n1483 VGND.n1481 0.688
R4346 VGND.n873 VGND.n853 0.688
R4347 VGND.n1366 VGND.n1365 0.688
R4348 VGND.n970 VGND.n968 0.688
R4349 VGND.n1420 VGND.n1419 0.688
R4350 VGND.n1385 VGND.n972 0.688
R4351 VGND.n874 VGND.n852 0.672375
R4352 VGND.n1332 VGND.n1316 0.65675
R4353 VGND.n1358 VGND.n1357 0.6255
R4354 VGND.n997 VGND.n936 0.6255
R4355 VGND.n999 VGND.n997 0.6255
R4356 VGND.n1001 VGND.n999 0.6255
R4357 VGND.n881 VGND.n852 0.609875
R4358 VGND.n53 VGND.n40 0.578625
R4359 VGND.n1474 VGND.n1473 0.547375
R4360 VGND.n1629 VGND.n800 0.542167
R4361 VGND.n1479 VGND.n1477 0.53175
R4362 VGND.n1470 VGND.n1468 0.516125
R4363 VGND.n874 VGND.n873 0.516125
R4364 VGND.n1365 VGND.n1339 0.516125
R4365 VGND.n1358 VGND.n1339 0.516125
R4366 VGND.n971 VGND.n970 0.5005
R4367 VGND.n1420 VGND.n971 0.5005
R4368 VGND.n1419 VGND.n1417 0.5005
R4369 VGND.n1417 VGND.n972 0.5005
R4370 VGND.n1293 VGND.n1014 0.472458
R4371 VGND.n866 VGND.n853 0.46925
R4372 VGND.n865 VGND.n864 0.46925
R4373 VGND.n855 VGND.n854 0.46925
R4374 VGND.n1347 VGND.n1340 0.46925
R4375 VGND.n1350 VGND.n1349 0.46925
R4376 VGND.n1450 VGND.n1449 0.438
R4377 VGND.n1455 VGND.n1453 0.438
R4378 VGND.n2496 VGND.n2484 0.411958
R4379 VGND.n1464 VGND.n1463 0.40675
R4380 VGND.n1366 VGND.n1017 0.40675
R4381 VGND.n1450 VGND.n1445 0.391125
R4382 VGND.n1453 VGND.n850 0.391125
R4383 VGND.n1464 VGND.n1459 0.391125
R4384 VGND.n1473 VGND.n1472 0.391125
R4385 VGND.n1407 VGND.n1406 0.3755
R4386 VGND.n1351 VGND.n1350 0.359875
R4387 VGND.n1445 VGND.n1443 0.34425
R4388 VGND.n1447 VGND.n850 0.34425
R4389 VGND.n1459 VGND.n1457 0.34425
R4390 VGND.n1461 VGND.n848 0.34425
R4391 VGND.n1472 VGND.n1470 0.34425
R4392 VGND.n1487 VGND.n1485 0.34425
R4393 VGND.n1481 VGND.n1479 0.34425
R4394 VGND.n1476 VGND.n5 0.34425
R4395 VGND.n866 VGND.n865 0.34425
R4396 VGND.n864 VGND.n863 0.34425
R4397 VGND.n856 VGND.n855 0.34425
R4398 VGND.n854 VGND.n8 0.34425
R4399 VGND.n1357 VGND.n1340 0.34425
R4400 VGND.n1348 VGND.n1347 0.34425
R4401 VGND.n1349 VGND.n11 0.34425
R4402 VGND.n1386 VGND.n1385 0.34425
R4403 VGND.n2533 VGND.n2532 0.3389
R4404 VGND.n38 VGND.n28 0.3205
R4405 VGND.n1431 VGND.n936 0.313
R4406 VGND.n1406 VGND.n1404 0.313
R4407 VGND.n909 VGND.n908 0.279967
R4408 VGND.n912 VGND.n897 0.279967
R4409 VGND.n922 VGND.n921 0.279967
R4410 VGND.n2529 VGND.n2528 0.26605
R4411 VGND.n863 VGND.n856 0.2505
R4412 VGND.n1407 VGND.n1001 0.2505
R4413 VGND.n1351 VGND.n1348 0.234875
R4414 VGND.n1014 VGND.n1013 0.219833
R4415 VGND.n1388 VGND.n1387 0.188
R4416 VGND.n1627 VGND.n1625 0.188
R4417 VGND.n1632 VGND.n1631 0.188
R4418 VGND.n956 VGND.n953 0.188
R4419 VGND.n1013 VGND.n14 0.172833
R4420 VGND.n2537 VGND.n2536 0.16108
R4421 VGND.n2495 VGND.n2494 0.1605
R4422 VGND.n27 VGND.n26 0.1605
R4423 VGND.n1392 VGND.n1388 0.15675
R4424 VGND.n958 VGND.n956 0.15675
R4425 VGND.n1333 VGND.n1293 0.132155
R4426 VGND.n903 VGND.n901 0.1255
R4427 VGND.n907 VGND.n901 0.1255
R4428 VGND.n892 VGND.n890 0.1255
R4429 VGND.n896 VGND.n890 0.1255
R4430 VGND.n1633 VGND.n797 0.1255
R4431 VGND.n2457 VGND.n55 0.1255
R4432 VGND.n1624 VGND.n803 0.1255
R4433 VGND.n916 VGND.n914 0.1255
R4434 VGND.n920 VGND.n914 0.1255
R4435 VGND.n2517 VGND.n2516 0.0804
R4436 VGND VGND.n2537 0.0647243
R4437 VGND.n797 VGND.n796 0.0626438
R4438 VGND.n55 VGND.n54 0.0626438
R4439 VGND.n803 VGND.n802 0.0626438
R4440 VGND.n1416 VGND.n973 0.0451429
R4441 VGND.n985 VGND.n973 0.0451429
R4442 VGND.n949 VGND.n942 0.0451429
R4443 VGND.n950 VGND.n949 0.0451429
R4444 VGND.n1313 VGND.n1296 0.0421667
R4445 VGND.n2525 VGND.n2524 0.029875
R4446 VGND.n2534 VGND.n3 0.0256998
R4447 VGND.n2530 VGND.n7 0.0256998
R4448 VGND.n2518 VGND.n16 0.0256998
R4449 VGND.n2526 VGND.n10 0.0256998
R4450 VGND.n2522 VGND.n13 0.0256998
R4451 VGND.n1631 VGND.n798 0.0217373
R4452 VGND.n1295 VGND.n800 0.0217373
R4453 VGND.n1626 VGND.n799 0.0217373
R4454 VGND.n801 VGND.n798 0.0217373
R4455 VGND.n1314 VGND.n1294 0.0217373
R4456 VGND.n1295 VGND.n1294 0.0217373
R4457 VGND.n1628 VGND.n801 0.0217373
R4458 VGND.n1630 VGND.n799 0.0217373
R4459 VGND.n1630 VGND.n1629 0.0217373
R4460 VGND.n1628 VGND.n1627 0.0217373
R4461 VGND.n1316 VGND.n1315 0.0217373
R4462 VGND.n1315 VGND.n1296 0.0217373
R4463 VGND.n2535 VGND.n2534 0.0200833
R4464 VGND.n2531 VGND.n2530 0.0200833
R4465 VGND.n2519 VGND.n2518 0.0200833
R4466 VGND.n2527 VGND.n2526 0.0200833
R4467 VGND.n2523 VGND.n2522 0.0200833
R4468 VGND.n2513 VGND.n2499 0.0185769
R4469 VGND.n2515 VGND.n2499 0.0185769
R4470 VGND.n2513 VGND.n2498 0.0100146
R4471 VGND.n2512 VGND.n2498 0.0100146
R4472 VGND.n2516 VGND.n2497 0.00803545
R4473 VGND.n2514 VGND.n2497 0.00803545
R4474 VGND.n2520 VGND.n15 0.0068649
R4475 VGND.n2524 VGND.n12 0.0068649
R4476 VGND.n2528 VGND.n9 0.0068649
R4477 VGND.n2532 VGND.n6 0.0068649
R4478 VGND.n2536 VGND.n2 0.0068649
R4479 VGND.n2533 VGND.n2 0.0068649
R4480 VGND.n2529 VGND.n6 0.0068649
R4481 VGND.n2525 VGND.n9 0.0068649
R4482 VGND.n2521 VGND.n12 0.0068649
R4483 VGND.n2517 VGND.n15 0.0068649
R4484 I_IN.n13 I_IN.n12 1269.42
R4485 I_IN.n2 I_IN.n0 299.368
R4486 I_IN.n2 I_IN.n1 299.252
R4487 I_IN.n4 I_IN.n3 299.252
R4488 I_IN.n6 I_IN.n5 299.252
R4489 I_IN.n8 I_IN.n7 299.252
R4490 I_IN.n10 I_IN.n9 299.252
R4491 I_IN.t13 I_IN.n13 275.325
R4492 I_IN.n16 I_IN.t7 238.891
R4493 I_IN.n14 I_IN.t13 178.34
R4494 I_IN.n14 I_IN.t15 178.34
R4495 I_IN.n16 I_IN.t10 161.371
R4496 I_IN.n15 I_IN.n14 152
R4497 I_IN.n12 I_IN.t18 151.792
R4498 I_IN.n13 I_IN.t15 80.3338
R4499 I_IN.n17 I_IN.n16 73.5727
R4500 I_IN.n15 I_IN.n11 68.0438
R4501 I_IN.n12 I_IN.t19 44.2902
R4502 I_IN.n0 I_IN.t5 39.4005
R4503 I_IN.n0 I_IN.t1 39.4005
R4504 I_IN.n1 I_IN.t6 39.4005
R4505 I_IN.n1 I_IN.t11 39.4005
R4506 I_IN.n3 I_IN.t8 39.4005
R4507 I_IN.n3 I_IN.t17 39.4005
R4508 I_IN.n5 I_IN.t9 39.4005
R4509 I_IN.n5 I_IN.t0 39.4005
R4510 I_IN.n7 I_IN.t12 39.4005
R4511 I_IN.n7 I_IN.t3 39.4005
R4512 I_IN.n9 I_IN.t2 39.4005
R4513 I_IN.n9 I_IN.t4 39.4005
R4514 I_IN.n17 I_IN.n15 15.7983
R4515 I_IN.n11 I_IN.t16 15.0005
R4516 I_IN.n11 I_IN.t14 15.0005
R4517 I_IN I_IN.n17 1.66073
R4518 I_IN.n10 I_IN.n8 0.115083
R4519 I_IN.n8 I_IN.n6 0.115083
R4520 I_IN.n6 I_IN.n4 0.115083
R4521 I_IN.n4 I_IN.n2 0.115083
R4522 I_IN I_IN.n10 3.29118
R4523 a_10710_11860.n13 a_10710_11860.t20 362.341
R4524 a_10710_11860.n3 a_10710_11860.t19 355.094
R4525 a_10710_11860.n3 a_10710_11860.n8 302.183
R4526 a_10710_11860.n3 a_10710_11860.n6 302.183
R4527 a_10710_11860.n14 a_10710_11860.n5 302.183
R4528 a_10710_11860.n4 a_10710_11860.t3 242.968
R4529 a_10710_11860.n11 a_10710_11860.n9 200.477
R4530 a_10710_11860.n11 a_10710_11860.n10 199.727
R4531 a_10710_11860.n12 a_10710_11860.t27 194.809
R4532 a_10710_11860.n12 a_10710_11860.t14 194.809
R4533 a_10710_11860.n7 a_10710_11860.t23 194.809
R4534 a_10710_11860.n7 a_10710_11860.t33 194.809
R4535 a_10710_11860.n3 a_10710_11860.n7 166.03
R4536 a_10710_11860.n4 a_10710_11860.n12 161.53
R4537 a_10710_11860.n10 a_10710_11860.t8 48.0005
R4538 a_10710_11860.n10 a_10710_11860.t5 48.0005
R4539 a_10710_11860.n9 a_10710_11860.t10 48.0005
R4540 a_10710_11860.n9 a_10710_11860.t6 48.0005
R4541 a_10710_11860.n13 a_10710_11860.n2 42.714
R4542 a_10710_11860.n8 a_10710_11860.t2 39.4005
R4543 a_10710_11860.n8 a_10710_11860.t1 39.4005
R4544 a_10710_11860.n6 a_10710_11860.t7 39.4005
R4545 a_10710_11860.n6 a_10710_11860.t9 39.4005
R4546 a_10710_11860.n14 a_10710_11860.t4 39.4005
R4547 a_10710_11860.t0 a_10710_11860.n14 39.4005
R4548 a_10710_11860.n4 a_10710_11860.n11 5.2505
R4549 a_10710_11860.n5 a_10710_11860.n4 4.92238
R4550 a_10710_11860.n0 a_10710_11860.t22 4.8248
R4551 a_10710_11860.n1 a_10710_11860.t15 4.5005
R4552 a_10710_11860.n1 a_10710_11860.t32 4.5005
R4553 a_10710_11860.n1 a_10710_11860.t36 4.5005
R4554 a_10710_11860.n0 a_10710_11860.t29 4.5005
R4555 a_10710_11860.n0 a_10710_11860.t25 4.5005
R4556 a_10710_11860.n0 a_10710_11860.t17 4.5005
R4557 a_10710_11860.n0 a_10710_11860.t21 4.5005
R4558 a_10710_11860.n0 a_10710_11860.t12 4.5005
R4559 a_10710_11860.n0 a_10710_11860.t18 4.5005
R4560 a_10710_11860.n1 a_10710_11860.t31 4.5005
R4561 a_10710_11860.n1 a_10710_11860.t26 4.5005
R4562 a_10710_11860.n2 a_10710_11860.t28 4.5005
R4563 a_10710_11860.n2 a_10710_11860.t24 4.5005
R4564 a_10710_11860.n2 a_10710_11860.t16 4.5005
R4565 a_10710_11860.n2 a_10710_11860.t34 4.5005
R4566 a_10710_11860.n2 a_10710_11860.t11 4.5005
R4567 a_10710_11860.n2 a_10710_11860.t30 4.5005
R4568 a_10710_11860.n2 a_10710_11860.t35 4.5005
R4569 a_10710_11860.n2 a_10710_11860.t13 4.5005
R4570 a_10710_11860.n2 a_10710_11860.n1 3.2388
R4571 a_10710_11860.n5 a_10710_11860.n13 2.90725
R4572 a_10710_11860.n1 a_10710_11860.n0 2.6325
R4573 a_10710_11860.n5 a_10710_11860.n3 2.2505
R4574 a_8454_18026.t0 a_8454_18026.t12 78.0006
R4575 a_8454_18026.t2 a_8454_18026.t18 0.1603
R4576 a_8454_18026.t6 a_8454_18026.t2 0.1603
R4577 a_8454_18026.t20 a_8454_18026.t6 0.1603
R4578 a_8454_18026.t3 a_8454_18026.t20 0.1603
R4579 a_8454_18026.t16 a_8454_18026.t3 0.1603
R4580 a_8454_18026.t11 a_8454_18026.t16 0.1603
R4581 a_8454_18026.t8 a_8454_18026.t11 0.1603
R4582 a_8454_18026.t9 a_8454_18026.t8 0.1603
R4583 a_8454_18026.t1 a_8454_18026.t4 0.1603
R4584 a_8454_18026.t7 a_8454_18026.t1 0.1603
R4585 a_8454_18026.t10 a_8454_18026.t7 0.1603
R4586 a_8454_18026.t15 a_8454_18026.t10 0.1603
R4587 a_8454_18026.t13 a_8454_18026.t15 0.1603
R4588 a_8454_18026.t19 a_8454_18026.t13 0.1603
R4589 a_8454_18026.t14 a_8454_18026.t19 0.1603
R4590 a_8454_18026.t12 a_8454_18026.t14 0.1603
R4591 a_8454_18026.t17 a_8454_18026.n0 0.159278
R4592 a_8454_18026.t4 a_8454_18026.t17 0.137822
R4593 a_8454_18026.n0 a_8454_18026.t9 0.1368
R4594 a_8454_18026.n0 a_8454_18026.t5 0.00152174
R4595 VDPWR.n162 VDPWR.n161 7755
R4596 VDPWR.n196 VDPWR.n161 7665
R4597 VDPWR.n196 VDPWR.n160 5025
R4598 VDPWR.n193 VDPWR.n160 2985
R4599 VDPWR.t34 VDPWR.t100 2804.76
R4600 VDPWR.t244 VDPWR.t81 2533.33
R4601 VDPWR.t188 VDPWR.t206 2307.14
R4602 VDPWR.t73 VDPWR.t61 2216.67
R4603 VDPWR.t283 VDPWR.t133 2216.67
R4604 VDPWR.t208 VDPWR.t395 2216.67
R4605 VDPWR.t227 VDPWR.t104 2126.19
R4606 VDPWR.t14 VDPWR.t40 1538.1
R4607 VDPWR.t424 VDPWR.t397 1492.86
R4608 VDPWR.t404 VDPWR.t250 1492.86
R4609 VDPWR.n45 VDPWR.t44 1289.29
R4610 VDPWR.n46 VDPWR.t402 1289.29
R4611 VDPWR.t75 VDPWR.t22 1130.95
R4612 VDPWR.t410 VDPWR.t220 1130.95
R4613 VDPWR.t118 VDPWR.t246 1130.95
R4614 VDPWR.t167 VDPWR.t102 1130.95
R4615 VDPWR.t48 VDPWR.t58 1130.95
R4616 VDPWR.n13 VDPWR.t371 927.381
R4617 VDPWR.n14 VDPWR.t4 927.381
R4618 VDPWR.n25 VDPWR.t194 927.381
R4619 VDPWR.n26 VDPWR.t30 927.381
R4620 VDPWR.n222 VDPWR.n213 831.25
R4621 VDPWR.n216 VDPWR.n215 831.25
R4622 VDPWR.n396 VDPWR.n210 831.25
R4623 VDPWR.n391 VDPWR.n390 831.25
R4624 VDPWR.n163 VDPWR.n159 827.201
R4625 VDPWR.n197 VDPWR.n159 817.601
R4626 VDPWR.n34 VDPWR.t49 740.534
R4627 VDPWR.n33 VDPWR.t105 740.534
R4628 VDPWR.t325 VDPWR.n521 708.125
R4629 VDPWR.n544 VDPWR.t325 708.125
R4630 VDPWR.n541 VDPWR.t301 708.125
R4631 VDPWR.t301 VDPWR.n522 708.125
R4632 VDPWR.t295 VDPWR.n501 708.125
R4633 VDPWR.n554 VDPWR.t295 708.125
R4634 VDPWR.n551 VDPWR.t311 708.125
R4635 VDPWR.t311 VDPWR.n502 708.125
R4636 VDPWR.t334 VDPWR.n624 708.125
R4637 VDPWR.n631 VDPWR.t334 708.125
R4638 VDPWR.t328 VDPWR.n651 708.125
R4639 VDPWR.n667 VDPWR.t328 708.125
R4640 VDPWR.t322 VDPWR.n638 708.125
R4641 VDPWR.n677 VDPWR.t322 708.125
R4642 VDPWR.n628 VDPWR.t355 694.444
R4643 VDPWR.t355 VDPWR.n625 694.444
R4644 VDPWR.n12 VDPWR.t62 663.801
R4645 VDPWR.n47 VDPWR.t84 663.801
R4646 VDPWR.n44 VDPWR.t101 663.801
R4647 VDPWR.n27 VDPWR.t189 663.801
R4648 VDPWR.n24 VDPWR.t396 663.801
R4649 VDPWR.n15 VDPWR.t284 663.801
R4650 VDPWR.n8 VDPWR.n6 662.297
R4651 VDPWR.n1 VDPWR.n0 661.734
R4652 VDPWR.n40 VDPWR.n39 661.734
R4653 VDPWR.n38 VDPWR.n37 661.734
R4654 VDPWR.n36 VDPWR.n35 661.734
R4655 VDPWR.n32 VDPWR.n31 661.734
R4656 VDPWR.n30 VDPWR.n29 661.734
R4657 VDPWR.n3 VDPWR.n2 661.734
R4658 VDPWR.n22 VDPWR.n21 661.734
R4659 VDPWR.n20 VDPWR.n19 661.734
R4660 VDPWR.n18 VDPWR.n17 661.734
R4661 VDPWR.n5 VDPWR.n4 661.734
R4662 VDPWR.n10 VDPWR.n9 661.734
R4663 VDPWR.n8 VDPWR.n7 661.734
R4664 VDPWR.n42 VDPWR.n41 660.514
R4665 VDPWR.n543 VDPWR.t324 657.76
R4666 VDPWR.n553 VDPWR.t294 657.76
R4667 VDPWR.n630 VDPWR.t333 640.794
R4668 VDPWR.n666 VDPWR.t327 640.794
R4669 VDPWR.n676 VDPWR.t321 640.794
R4670 VDPWR.t61 VDPWR.n13 610.715
R4671 VDPWR.n14 VDPWR.t283 610.715
R4672 VDPWR.t395 VDPWR.n25 610.715
R4673 VDPWR.n26 VDPWR.t188 610.715
R4674 VDPWR.t100 VDPWR.n45 610.715
R4675 VDPWR.n46 VDPWR.t83 610.715
R4676 VDPWR.n577 VDPWR.n575 587.407
R4677 VDPWR.n581 VDPWR.n578 587.407
R4678 VDPWR.n607 VDPWR.n606 587.407
R4679 VDPWR.n602 VDPWR.n568 587.407
R4680 VDPWR.n491 VDPWR.n490 585
R4681 VDPWR.n470 VDPWR.n435 585
R4682 VDPWR.n606 VDPWR.n605 585
R4683 VDPWR.n604 VDPWR.n602 585
R4684 VDPWR.n588 VDPWR.n577 585
R4685 VDPWR.n585 VDPWR.n578 585
R4686 VDPWR.n211 VDPWR.n210 585
R4687 VDPWR.n393 VDPWR.n391 585
R4688 VDPWR.n214 VDPWR.n213 585
R4689 VDPWR.n219 VDPWR.n216 585
R4690 VDPWR.n309 VDPWR.n245 585
R4691 VDPWR.n304 VDPWR.n245 585
R4692 VDPWR.n253 VDPWR.n246 585
R4693 VDPWR.n248 VDPWR.n246 585
R4694 VDPWR.n300 VDPWR.n255 585
R4695 VDPWR.n293 VDPWR.n255 585
R4696 VDPWR.n290 VDPWR.n262 585
R4697 VDPWR.n285 VDPWR.n262 585
R4698 VDPWR.n270 VDPWR.n263 585
R4699 VDPWR.n265 VDPWR.n263 585
R4700 VDPWR.n282 VDPWR.n271 585
R4701 VDPWR.n278 VDPWR.n271 585
R4702 VDPWR.n126 VDPWR.n125 585
R4703 VDPWR.n119 VDPWR.n117 585
R4704 VDPWR.n148 VDPWR.n147 585
R4705 VDPWR.n141 VDPWR.n139 585
R4706 VDPWR.n179 VDPWR.n178 585
R4707 VDPWR.n172 VDPWR.n170 585
R4708 VDPWR.n104 VDPWR.n53 585
R4709 VDPWR.n108 VDPWR.n53 585
R4710 VDPWR.n97 VDPWR.n59 585
R4711 VDPWR.n88 VDPWR.n59 585
R4712 VDPWR.n77 VDPWR.n76 585
R4713 VDPWR.n77 VDPWR.n64 585
R4714 VDPWR.n127 VDPWR.n126 584.514
R4715 VDPWR.n120 VDPWR.n119 584.514
R4716 VDPWR.n149 VDPWR.n148 584.514
R4717 VDPWR.n142 VDPWR.n141 584.514
R4718 VDPWR.n180 VDPWR.n179 584.514
R4719 VDPWR.n173 VDPWR.n172 584.514
R4720 VDPWR.t354 VDPWR.n629 557.783
R4721 VDPWR.t300 VDPWR.n542 540.818
R4722 VDPWR.t310 VDPWR.n552 540.818
R4723 VDPWR.t336 VDPWR.n665 523.855
R4724 VDPWR.t330 VDPWR.n675 523.855
R4725 VDPWR.n118 VDPWR.t430 500.986
R4726 VDPWR.n140 VDPWR.t428 500.986
R4727 VDPWR.n171 VDPWR.t432 500.986
R4728 VDPWR.t22 VDPWR.t380 497.62
R4729 VDPWR.t371 VDPWR.t75 497.62
R4730 VDPWR.t220 VDPWR.t73 497.62
R4731 VDPWR.t4 VDPWR.t410 497.62
R4732 VDPWR.t133 VDPWR.t118 497.62
R4733 VDPWR.t246 VDPWR.t194 497.62
R4734 VDPWR.t102 VDPWR.t208 497.62
R4735 VDPWR.t30 VDPWR.t167 497.62
R4736 VDPWR.t206 VDPWR.t424 497.62
R4737 VDPWR.t397 VDPWR.t227 497.62
R4738 VDPWR.t104 VDPWR.t48 497.62
R4739 VDPWR.t58 VDPWR.t14 497.62
R4740 VDPWR.t40 VDPWR.t44 497.62
R4741 VDPWR.t32 VDPWR.t34 497.62
R4742 VDPWR.t250 VDPWR.t32 497.62
R4743 VDPWR.t81 VDPWR.t404 497.62
R4744 VDPWR.t402 VDPWR.t244 497.62
R4745 VDPWR.n221 VDPWR.t159 465.079
R4746 VDPWR.t159 VDPWR.n220 465.079
R4747 VDPWR.n395 VDPWR.t172 465.079
R4748 VDPWR.t172 VDPWR.n394 465.079
R4749 VDPWR.n356 VDPWR.t39 464.281
R4750 VDPWR.t39 VDPWR.n355 464.281
R4751 VDPWR.t72 VDPWR.n204 464.281
R4752 VDPWR.n400 VDPWR.t72 464.281
R4753 VDPWR.n410 VDPWR.t178 464.281
R4754 VDPWR.t178 VDPWR.n409 464.281
R4755 VDPWR.t107 VDPWR.n226 464.281
R4756 VDPWR.n370 VDPWR.t107 464.281
R4757 VDPWR.n380 VDPWR.t233 464.281
R4758 VDPWR.t233 VDPWR.n379 464.281
R4759 VDPWR.n365 VDPWR.t3 464.281
R4760 VDPWR.t3 VDPWR.n364 464.281
R4761 VDPWR.t415 VDPWR.n337 464.281
R4762 VDPWR.n340 VDPWR.t415 464.281
R4763 VDPWR.n332 VDPWR.t161 464.281
R4764 VDPWR.t161 VDPWR.n235 464.281
R4765 VDPWR.n325 VDPWR.t109 464.281
R4766 VDPWR.t109 VDPWR.n324 464.281
R4767 VDPWR.n315 VDPWR.t421 464.281
R4768 VDPWR.t421 VDPWR.n239 464.281
R4769 VDPWR.n133 VDPWR.t383 461.389
R4770 VDPWR.t383 VDPWR.n132 461.389
R4771 VDPWR.n155 VDPWR.t55 461.389
R4772 VDPWR.t55 VDPWR.n154 461.389
R4773 VDPWR.n186 VDPWR.t413 461.389
R4774 VDPWR.t413 VDPWR.n185 461.389
R4775 VDPWR.n633 VDPWR.t332 422.384
R4776 VDPWR.n626 VDPWR.t353 422.384
R4777 VDPWR.n669 VDPWR.t326 418.368
R4778 VDPWR.n662 VDPWR.t335 418.368
R4779 VDPWR.n679 VDPWR.t320 418.368
R4780 VDPWR.n672 VDPWR.t329 418.368
R4781 VDPWR.n254 VDPWR.t429 411.101
R4782 VDPWR.t324 VDPWR.t279 407.144
R4783 VDPWR.t279 VDPWR.t248 407.144
R4784 VDPWR.t248 VDPWR.t285 407.144
R4785 VDPWR.t285 VDPWR.t151 407.144
R4786 VDPWR.t151 VDPWR.t216 407.144
R4787 VDPWR.t216 VDPWR.t271 407.144
R4788 VDPWR.t271 VDPWR.t275 407.144
R4789 VDPWR.t275 VDPWR.t96 407.144
R4790 VDPWR.t96 VDPWR.t52 407.144
R4791 VDPWR.t52 VDPWR.t240 407.144
R4792 VDPWR.t240 VDPWR.t94 407.144
R4793 VDPWR.t94 VDPWR.t281 407.144
R4794 VDPWR.t281 VDPWR.t273 407.144
R4795 VDPWR.t273 VDPWR.t182 407.144
R4796 VDPWR.t182 VDPWR.t0 407.144
R4797 VDPWR.t0 VDPWR.t179 407.144
R4798 VDPWR.t179 VDPWR.t149 407.144
R4799 VDPWR.t149 VDPWR.t277 407.144
R4800 VDPWR.t277 VDPWR.t300 407.144
R4801 VDPWR.t294 VDPWR.t257 407.144
R4802 VDPWR.t257 VDPWR.t50 407.144
R4803 VDPWR.t50 VDPWR.t126 407.144
R4804 VDPWR.t126 VDPWR.t289 407.144
R4805 VDPWR.t289 VDPWR.t184 407.144
R4806 VDPWR.t184 VDPWR.t263 407.144
R4807 VDPWR.t263 VDPWR.t259 407.144
R4808 VDPWR.t259 VDPWR.t65 407.144
R4809 VDPWR.t65 VDPWR.t140 407.144
R4810 VDPWR.t140 VDPWR.t69 407.144
R4811 VDPWR.t69 VDPWR.t364 407.144
R4812 VDPWR.t364 VDPWR.t253 407.144
R4813 VDPWR.t253 VDPWR.t255 407.144
R4814 VDPWR.t255 VDPWR.t251 407.144
R4815 VDPWR.t251 VDPWR.t287 407.144
R4816 VDPWR.t287 VDPWR.t291 407.144
R4817 VDPWR.t291 VDPWR.t20 407.144
R4818 VDPWR.t20 VDPWR.t261 407.144
R4819 VDPWR.t261 VDPWR.t310 407.144
R4820 VDPWR.n475 VDPWR.t347 384.967
R4821 VDPWR.n479 VDPWR.t312 384.967
R4822 VDPWR.n442 VDPWR.t350 384.967
R4823 VDPWR.n446 VDPWR.t360 384.967
R4824 VDPWR.n47 VDPWR.n46 382.8
R4825 VDPWR.n45 VDPWR.n44 382.8
R4826 VDPWR.n27 VDPWR.n26 382.8
R4827 VDPWR.n25 VDPWR.n24 382.8
R4828 VDPWR.n15 VDPWR.n14 382.8
R4829 VDPWR.n13 VDPWR.n12 382.8
R4830 VDPWR.t333 VDPWR.t219 373.214
R4831 VDPWR.t219 VDPWR.t218 373.214
R4832 VDPWR.t218 VDPWR.t354 373.214
R4833 VDPWR.t327 VDPWR.t390 373.214
R4834 VDPWR.t390 VDPWR.t406 373.214
R4835 VDPWR.t406 VDPWR.t24 373.214
R4836 VDPWR.t24 VDPWR.t124 373.214
R4837 VDPWR.t124 VDPWR.t155 373.214
R4838 VDPWR.t155 VDPWR.t128 373.214
R4839 VDPWR.t128 VDPWR.t26 373.214
R4840 VDPWR.t26 VDPWR.t374 373.214
R4841 VDPWR.t374 VDPWR.t222 373.214
R4842 VDPWR.t222 VDPWR.t200 373.214
R4843 VDPWR.t200 VDPWR.t336 373.214
R4844 VDPWR.t321 VDPWR.t77 373.214
R4845 VDPWR.t77 VDPWR.t214 373.214
R4846 VDPWR.t214 VDPWR.t63 373.214
R4847 VDPWR.t63 VDPWR.t164 373.214
R4848 VDPWR.t164 VDPWR.t9 373.214
R4849 VDPWR.t9 VDPWR.t162 373.214
R4850 VDPWR.t162 VDPWR.t392 373.214
R4851 VDPWR.t392 VDPWR.t115 373.214
R4852 VDPWR.t115 VDPWR.t204 373.214
R4853 VDPWR.t204 VDPWR.t79 373.214
R4854 VDPWR.t79 VDPWR.t330 373.214
R4855 VDPWR.n546 VDPWR.t323 370.168
R4856 VDPWR.n539 VDPWR.t299 370.168
R4857 VDPWR.n556 VDPWR.t293 370.168
R4858 VDPWR.n549 VDPWR.t309 370.168
R4859 VDPWR.n460 VDPWR.t344 362.134
R4860 VDPWR.n559 VDPWR.t296 360.868
R4861 VDPWR.n613 VDPWR.t338 360.868
R4862 VDPWR.t307 VDPWR.t225 360.346
R4863 VDPWR.t225 VDPWR.t238 360.346
R4864 VDPWR.t238 VDPWR.t190 360.346
R4865 VDPWR.t190 VDPWR.t231 360.346
R4866 VDPWR.t231 VDPWR.t357 360.346
R4867 VDPWR.t18 VDPWR.t342 360.346
R4868 VDPWR.t234 VDPWR.t18 360.346
R4869 VDPWR.t236 VDPWR.t234 360.346
R4870 VDPWR.t153 VDPWR.t236 360.346
R4871 VDPWR.t303 VDPWR.t153 360.346
R4872 VDPWR.n496 VDPWR.t316 352.834
R4873 VDPWR.n653 VDPWR.t337 351.793
R4874 VDPWR.n640 VDPWR.t331 351.793
R4875 VDPWR.n198 VDPWR.n197 347.2
R4876 VDPWR.n74 VDPWR.t307 343.966
R4877 VDPWR.n99 VDPWR.t357 343.966
R4878 VDPWR.t342 VDPWR.n99 343.966
R4879 VDPWR.n106 VDPWR.t303 343.966
R4880 VDPWR.n480 VDPWR.t315 341.752
R4881 VDPWR.n474 VDPWR.t349 341.752
R4882 VDPWR.n445 VDPWR.t363 341.752
R4883 VDPWR.n441 VDPWR.t352 341.752
R4884 VDPWR.n57 VDPWR.t341 336.329
R4885 VDPWR.n57 VDPWR.t356 336.329
R4886 VDPWR.n62 VDPWR.t306 330
R4887 VDPWR.n110 VDPWR.t302 330
R4888 VDPWR.n448 VDPWR.n439 315.647
R4889 VDPWR.n447 VDPWR.n444 315.647
R4890 VDPWR.n443 VDPWR.n440 315.647
R4891 VDPWR.t132 VDPWR.t117 314.113
R4892 VDPWR.t11 VDPWR.t171 314.113
R4893 VDPWR.n477 VDPWR.n429 313.846
R4894 VDPWR.n478 VDPWR.n427 313.846
R4895 VDPWR.n476 VDPWR.n430 313.846
R4896 VDPWR.n232 VDPWR.t177 308.849
R4897 VDPWR.n441 VDPWR.t351 304.659
R4898 VDPWR.n661 VDPWR.n660 301.933
R4899 VDPWR.n659 VDPWR.n658 301.933
R4900 VDPWR.n657 VDPWR.n656 301.933
R4901 VDPWR.n655 VDPWR.n654 301.933
R4902 VDPWR.n650 VDPWR.n649 301.933
R4903 VDPWR.n648 VDPWR.n647 301.933
R4904 VDPWR.n646 VDPWR.n645 301.933
R4905 VDPWR.n644 VDPWR.n643 301.933
R4906 VDPWR.n642 VDPWR.n641 301.933
R4907 VDPWR.n637 VDPWR.n636 301.933
R4908 VDPWR.n538 VDPWR.n537 299.231
R4909 VDPWR.n536 VDPWR.n535 299.231
R4910 VDPWR.n534 VDPWR.n533 299.231
R4911 VDPWR.n532 VDPWR.n531 299.231
R4912 VDPWR.n530 VDPWR.n529 299.231
R4913 VDPWR.n528 VDPWR.n527 299.231
R4914 VDPWR.n526 VDPWR.n525 299.231
R4915 VDPWR.n524 VDPWR.n523 299.231
R4916 VDPWR.n520 VDPWR.n519 299.231
R4917 VDPWR.n518 VDPWR.n517 299.231
R4918 VDPWR.n516 VDPWR.n515 299.231
R4919 VDPWR.n514 VDPWR.n513 299.231
R4920 VDPWR.n512 VDPWR.n511 299.231
R4921 VDPWR.n510 VDPWR.n509 299.231
R4922 VDPWR.n508 VDPWR.n507 299.231
R4923 VDPWR.n506 VDPWR.n505 299.231
R4924 VDPWR.n504 VDPWR.n503 299.231
R4925 VDPWR.n500 VDPWR.n499 299.231
R4926 VDPWR.n84 VDPWR.n59 291.363
R4927 VDPWR.n96 VDPWR.n95 291.363
R4928 VDPWR.n95 VDPWR.n61 291.363
R4929 VDPWR.n490 VDPWR.n489 290.733
R4930 VDPWR.n490 VDPWR.n425 290.733
R4931 VDPWR.n438 VDPWR.n435 290.733
R4932 VDPWR.n463 VDPWR.n435 290.733
R4933 VDPWR.n307 VDPWR.n245 290.733
R4934 VDPWR.n247 VDPWR.n246 290.733
R4935 VDPWR.n294 VDPWR.n255 290.733
R4936 VDPWR.n288 VDPWR.n262 290.733
R4937 VDPWR.n264 VDPWR.n263 290.733
R4938 VDPWR.n276 VDPWR.n271 290.733
R4939 VDPWR.n101 VDPWR.n53 290.733
R4940 VDPWR.n77 VDPWR.n63 290.733
R4941 VDPWR.t90 VDPWR.t297 251.471
R4942 VDPWR.t92 VDPWR.t90 251.471
R4943 VDPWR.t366 VDPWR.t92 251.471
R4944 VDPWR.t400 VDPWR.t366 251.471
R4945 VDPWR.t110 VDPWR.t400 251.471
R4946 VDPWR.t197 VDPWR.t110 251.471
R4947 VDPWR.t145 VDPWR.t197 251.471
R4948 VDPWR.t212 VDPWR.t145 251.471
R4949 VDPWR.t143 VDPWR.t212 251.471
R4950 VDPWR.t138 VDPWR.t143 251.471
R4951 VDPWR.t416 VDPWR.t138 251.471
R4952 VDPWR.t418 VDPWR.t416 251.471
R4953 VDPWR.t210 VDPWR.t418 251.471
R4954 VDPWR.t174 VDPWR.t210 251.471
R4955 VDPWR.t147 VDPWR.t174 251.471
R4956 VDPWR.t386 VDPWR.t147 251.471
R4957 VDPWR.t339 VDPWR.t386 251.471
R4958 VDPWR.n411 VDPWR.n410 243.698
R4959 VDPWR.n381 VDPWR.n380 243.698
R4960 VDPWR.n357 VDPWR.n356 243.698
R4961 VDPWR.n333 VDPWR.n332 243.698
R4962 VDPWR.n316 VDPWR.n315 243.698
R4963 VDPWR.n404 VDPWR.n400 243.698
R4964 VDPWR.n374 VDPWR.n370 243.698
R4965 VDPWR.n364 VDPWR.n359 243.698
R4966 VDPWR.n340 VDPWR.n339 243.698
R4967 VDPWR.n324 VDPWR.n237 243.698
R4968 VDPWR.n542 VDPWR.n541 238.367
R4969 VDPWR.n542 VDPWR.n522 238.367
R4970 VDPWR.n552 VDPWR.n551 238.367
R4971 VDPWR.n552 VDPWR.n502 238.367
R4972 VDPWR.n609 VDPWR.n608 238.367
R4973 VDPWR.n629 VDPWR.n628 238.367
R4974 VDPWR.n629 VDPWR.n625 238.367
R4975 VDPWR.n665 VDPWR.n664 238.367
R4976 VDPWR.n665 VDPWR.n652 238.367
R4977 VDPWR.n675 VDPWR.n674 238.367
R4978 VDPWR.n675 VDPWR.n639 238.367
R4979 VDPWR.n399 VDPWR.n203 238.367
R4980 VDPWR.n397 VDPWR.n396 238.367
R4981 VDPWR.n390 VDPWR.n206 238.367
R4982 VDPWR.n369 VDPWR.n225 238.367
R4983 VDPWR.n352 VDPWR.n229 238.367
R4984 VDPWR.n336 VDPWR.n335 238.367
R4985 VDPWR.n319 VDPWR.n318 238.367
R4986 VDPWR.n414 VDPWR.n413 238.367
R4987 VDPWR.n222 VDPWR.n208 238.367
R4988 VDPWR.n384 VDPWR.n383 238.367
R4989 VDPWR.n367 VDPWR.n366 238.367
R4990 VDPWR.n345 VDPWR.n344 238.367
R4991 VDPWR.n327 VDPWR.n326 238.367
R4992 VDPWR.n215 VDPWR.n207 238.367
R4993 VDPWR.t297 VDPWR.n593 237.5
R4994 VDPWR.n610 VDPWR.t339 237.5
R4995 VDPWR.n190 VDPWR.t121 236.043
R4996 VDPWR.n492 VDPWR.n491 230.308
R4997 VDPWR.n495 VDPWR.n494 230.308
R4998 VDPWR.n462 VDPWR.n433 230.308
R4999 VDPWR.n310 VDPWR.n309 230.308
R5000 VDPWR.n304 VDPWR.n241 230.308
R5001 VDPWR.n291 VDPWR.n290 230.308
R5002 VDPWR.n285 VDPWR.n258 230.308
R5003 VDPWR.n253 VDPWR.n243 230.308
R5004 VDPWR.n300 VDPWR.n299 230.308
R5005 VDPWR.n297 VDPWR.n293 230.308
R5006 VDPWR.n270 VDPWR.n260 230.308
R5007 VDPWR.n265 VDPWR.n259 230.308
R5008 VDPWR.n248 VDPWR.n242 230.308
R5009 VDPWR.n105 VDPWR.n104 230.308
R5010 VDPWR.n108 VDPWR.n107 230.308
R5011 VDPWR.n98 VDPWR.n97 230.308
R5012 VDPWR.n88 VDPWR.n55 230.308
R5013 VDPWR.t6 VDPWR.t186 222.178
R5014 VDPWR.n192 VDPWR.n163 221.601
R5015 VDPWR.t412 VDPWR.t120 221.525
R5016 VDPWR.n317 VDPWR.n311 199.195
R5017 VDPWR.n445 VDPWR.n431 185.001
R5018 VDPWR.n474 VDPWR.n473 185.001
R5019 VDPWR.n481 VDPWR.n480 185.001
R5020 VDPWR.n485 VDPWR.n483 185
R5021 VDPWR.n488 VDPWR.n482 185
R5022 VDPWR.n493 VDPWR.n482 185
R5023 VDPWR.n487 VDPWR.n426 185
R5024 VDPWR.n471 VDPWR.n470 185
R5025 VDPWR.n472 VDPWR.n471 185
R5026 VDPWR.n436 VDPWR.n434 185
R5027 VDPWR.n467 VDPWR.n466 185
R5028 VDPWR.n465 VDPWR.n464 185
R5029 VDPWR.n598 VDPWR.n596 185
R5030 VDPWR.n605 VDPWR.n595 185
R5031 VDPWR.n610 VDPWR.n595 185
R5032 VDPWR.n604 VDPWR.n603 185
R5033 VDPWR.n601 VDPWR.n570 185
R5034 VDPWR.n612 VDPWR.n611 185
R5035 VDPWR.n611 VDPWR.n610 185
R5036 VDPWR.n592 VDPWR.n591 185
R5037 VDPWR.n593 VDPWR.n592 185
R5038 VDPWR.n589 VDPWR.n574 185
R5039 VDPWR.n588 VDPWR.n587 185
R5040 VDPWR.n586 VDPWR.n585 185
R5041 VDPWR.n580 VDPWR.n579 185
R5042 VDPWR.n582 VDPWR.n573 185
R5043 VDPWR.n593 VDPWR.n573 185
R5044 VDPWR.n269 VDPWR.n268 185
R5045 VDPWR.n267 VDPWR.n266 185
R5046 VDPWR.n257 VDPWR.n256 185
R5047 VDPWR.n296 VDPWR.n295 185
R5048 VDPWR.n252 VDPWR.n251 185
R5049 VDPWR.n250 VDPWR.n249 185
R5050 VDPWR.n321 VDPWR.n238 185
R5051 VDPWR.n323 VDPWR.n322 185
R5052 VDPWR.n343 VDPWR.n342 185
R5053 VDPWR.n341 VDPWR.n338 185
R5054 VDPWR.n361 VDPWR.n360 185
R5055 VDPWR.n363 VDPWR.n362 185
R5056 VDPWR.n371 VDPWR.n227 185
R5057 VDPWR.n373 VDPWR.n372 185
R5058 VDPWR.n217 VDPWR.n214 185
R5059 VDPWR.n219 VDPWR.n218 185
R5060 VDPWR.n401 VDPWR.n205 185
R5061 VDPWR.n403 VDPWR.n402 185
R5062 VDPWR.n289 VDPWR.n261 185
R5063 VDPWR.n287 VDPWR.n286 185
R5064 VDPWR.n308 VDPWR.n244 185
R5065 VDPWR.n306 VDPWR.n305 185
R5066 VDPWR.n314 VDPWR.n312 185
R5067 VDPWR.n313 VDPWR.n240 185
R5068 VDPWR.n331 VDPWR.n329 185
R5069 VDPWR.n330 VDPWR.n236 185
R5070 VDPWR.n231 VDPWR.n230 185
R5071 VDPWR.n354 VDPWR.n353 185
R5072 VDPWR.n376 VDPWR.n375 185
R5073 VDPWR.n378 VDPWR.n377 185
R5074 VDPWR.n211 VDPWR.n209 185
R5075 VDPWR.n393 VDPWR.n392 185
R5076 VDPWR.n406 VDPWR.n405 185
R5077 VDPWR.n408 VDPWR.n407 185
R5078 VDPWR.n282 VDPWR.n281 185
R5079 VDPWR.n281 VDPWR.n280 185
R5080 VDPWR.n273 VDPWR.n272 185
R5081 VDPWR.n277 VDPWR.n275 185
R5082 VDPWR.n279 VDPWR.n278 185
R5083 VDPWR.n280 VDPWR.n279 185
R5084 VDPWR.n193 VDPWR.n192 185
R5085 VDPWR.n60 VDPWR.n56 185
R5086 VDPWR.n86 VDPWR.n85 185
R5087 VDPWR.n102 VDPWR.n100 185
R5088 VDPWR.n54 VDPWR.n52 185
R5089 VDPWR.n76 VDPWR.n75 185
R5090 VDPWR.n75 VDPWR.n74 185
R5091 VDPWR.n67 VDPWR.n66 185
R5092 VDPWR.n72 VDPWR.n71 185
R5093 VDPWR.n73 VDPWR.n64 185
R5094 VDPWR.n74 VDPWR.n73 185
R5095 VDPWR.n280 VDPWR.t6 172.38
R5096 VDPWR.t229 VDPWR.n292 172.38
R5097 VDPWR.n298 VDPWR.t98 172.38
R5098 VDPWR.n97 VDPWR.n57 166.63
R5099 VDPWR.n194 VDPWR.n193 164.12
R5100 VDPWR.t382 VDPWR.t224 163.588
R5101 VDPWR.n191 VDPWR.n165 153.601
R5102 VDPWR.n198 VDPWR.n158 153.601
R5103 VDPWR.n50 VDPWR.n49 153.573
R5104 VDPWR.n92 VDPWR.n91 153.573
R5105 VDPWR.n94 VDPWR.n93 153.573
R5106 VDPWR.n83 VDPWR.n82 153.573
R5107 VDPWR.n81 VDPWR.n80 153.573
R5108 VDPWR.n79 VDPWR.n78 153.573
R5109 VDPWR.n596 VDPWR.n595 150
R5110 VDPWR.n603 VDPWR.n595 150
R5111 VDPWR.n611 VDPWR.n570 150
R5112 VDPWR.n592 VDPWR.n574 150
R5113 VDPWR.n587 VDPWR.n586 150
R5114 VDPWR.n579 VDPWR.n573 150
R5115 VDPWR.n407 VDPWR.n405 150
R5116 VDPWR.n392 VDPWR.n209 150
R5117 VDPWR.n377 VDPWR.n375 150
R5118 VDPWR.n353 VDPWR.n230 150
R5119 VDPWR.n329 VDPWR.n236 150
R5120 VDPWR.n312 VDPWR.n240 150
R5121 VDPWR.n403 VDPWR.n205 150
R5122 VDPWR.n218 VDPWR.n217 150
R5123 VDPWR.n373 VDPWR.n227 150
R5124 VDPWR.n362 VDPWR.n360 150
R5125 VDPWR.n343 VDPWR.n338 150
R5126 VDPWR.n322 VDPWR.n238 150
R5127 VDPWR.t67 VDPWR.t88 145.038
R5128 VDPWR.n165 VDPWR.n164 144
R5129 VDPWR.n614 VDPWR.n567 141.712
R5130 VDPWR.n615 VDPWR.n566 141.712
R5131 VDPWR.n616 VDPWR.n565 141.712
R5132 VDPWR.n617 VDPWR.n564 141.712
R5133 VDPWR.n618 VDPWR.n563 141.712
R5134 VDPWR.n619 VDPWR.n562 141.712
R5135 VDPWR.n620 VDPWR.n561 141.712
R5136 VDPWR.n621 VDPWR.n560 141.712
R5137 VDPWR.n334 VDPWR.n328 137.904
R5138 VDPWR.n358 VDPWR.n228 137.904
R5139 VDPWR.n280 VDPWR.t408 126.412
R5140 VDPWR.n292 VDPWR.t186 126.412
R5141 VDPWR.n298 VDPWR.t229 126.412
R5142 VDPWR.n311 VDPWR.t98 126.412
R5143 VDPWR.n423 VDPWR.n422 123.987
R5144 VDPWR.n450 VDPWR.n449 123.987
R5145 VDPWR.n452 VDPWR.n451 123.987
R5146 VDPWR.n458 VDPWR.n457 123.987
R5147 VDPWR.t298 VDPWR.n577 123.126
R5148 VDPWR.n578 VDPWR.t298 123.126
R5149 VDPWR.n606 VDPWR.t340 123.126
R5150 VDPWR.n602 VDPWR.t340 123.126
R5151 VDPWR.t43 VDPWR.n213 123.126
R5152 VDPWR.n216 VDPWR.t43 123.126
R5153 VDPWR.t199 VDPWR.n210 123.126
R5154 VDPWR.n391 VDPWR.t199 123.126
R5155 VDPWR.n126 VDPWR.t268 123.126
R5156 VDPWR.n119 VDPWR.t268 123.126
R5157 VDPWR.n148 VDPWR.t270 123.126
R5158 VDPWR.n141 VDPWR.t270 123.126
R5159 VDPWR.n179 VDPWR.t266 123.126
R5160 VDPWR.n172 VDPWR.t266 123.126
R5161 VDPWR.n483 VDPWR.n482 120.001
R5162 VDPWR.n482 VDPWR.n426 120.001
R5163 VDPWR.n471 VDPWR.n434 120.001
R5164 VDPWR.n466 VDPWR.n465 120.001
R5165 VDPWR.n305 VDPWR.n244 120.001
R5166 VDPWR.n286 VDPWR.n261 120.001
R5167 VDPWR.n251 VDPWR.n250 120.001
R5168 VDPWR.n296 VDPWR.n257 120.001
R5169 VDPWR.n268 VDPWR.n267 120.001
R5170 VDPWR.n281 VDPWR.n273 120.001
R5171 VDPWR.n279 VDPWR.n275 120.001
R5172 VDPWR.n100 VDPWR.n54 120.001
R5173 VDPWR.n85 VDPWR.n56 120.001
R5174 VDPWR.n75 VDPWR.n67 120.001
R5175 VDPWR.n73 VDPWR.n72 120.001
R5176 VDPWR.t361 VDPWR.n431 119.656
R5177 VDPWR.n454 VDPWR.n453 119.424
R5178 VDPWR.n196 VDPWR.t166 115.386
R5179 VDPWR.n473 VDPWR.n472 108.779
R5180 VDPWR.n382 VDPWR.n368 107.258
R5181 VDPWR.n382 VDPWR.t106 103.427
R5182 VDPWR.n398 VDPWR.t158 103.427
R5183 VDPWR.t42 VDPWR.n398 103.427
R5184 VDPWR.n412 VDPWR.t71 103.427
R5185 VDPWR.t54 VDPWR.n195 102.243
R5186 VDPWR.n368 VDPWR.t38 95.7666
R5187 VDPWR.t351 VDPWR.t113 94.2753
R5188 VDPWR.t113 VDPWR.t12 94.2753
R5189 VDPWR.t12 VDPWR.t7 94.2753
R5190 VDPWR.t7 VDPWR.t16 94.2753
R5191 VDPWR.t16 VDPWR.t361 94.2753
R5192 VDPWR.t369 VDPWR.t28 94.2753
R5193 VDPWR.t242 VDPWR.t313 94.2753
R5194 VDPWR.n481 VDPWR.t130 94.2753
R5195 VDPWR.t85 VDPWR.t373 94.2753
R5196 VDPWR.t157 VDPWR.t394 94.2753
R5197 VDPWR.n164 VDPWR.n160 92.5005
R5198 VDPWR.n195 VDPWR.n160 92.5005
R5199 VDPWR.n161 VDPWR.n159 92.5005
R5200 VDPWR.n195 VDPWR.n161 92.5005
R5201 VDPWR.t108 VDPWR.t420 91.936
R5202 VDPWR.t414 VDPWR.t160 91.936
R5203 VDPWR.t120 VDPWR.n194 89.6985
R5204 VDPWR.t2 VDPWR.t176 84.2747
R5205 VDPWR.t106 VDPWR.t132 84.2747
R5206 VDPWR.t117 VDPWR.t158 84.2747
R5207 VDPWR.t171 VDPWR.t42 84.2747
R5208 VDPWR.t71 VDPWR.t11 84.2747
R5209 VDPWR.t345 VDPWR.t348 83.3974
R5210 VDPWR.t60 VDPWR.t86 83.3974
R5211 VDPWR.n477 VDPWR.n476 83.2005
R5212 VDPWR.n478 VDPWR.n477 83.2005
R5213 VDPWR.n448 VDPWR.n443 83.2005
R5214 VDPWR.n448 VDPWR.n447 83.2005
R5215 VDPWR.n0 VDPWR.t245 78.8005
R5216 VDPWR.n0 VDPWR.t403 78.8005
R5217 VDPWR.n39 VDPWR.t405 78.8005
R5218 VDPWR.n39 VDPWR.t82 78.8005
R5219 VDPWR.n41 VDPWR.t35 78.8005
R5220 VDPWR.n41 VDPWR.t33 78.8005
R5221 VDPWR.n37 VDPWR.t41 78.8005
R5222 VDPWR.n37 VDPWR.t45 78.8005
R5223 VDPWR.n35 VDPWR.t59 78.8005
R5224 VDPWR.n35 VDPWR.t15 78.8005
R5225 VDPWR.n31 VDPWR.t398 78.8005
R5226 VDPWR.n31 VDPWR.t228 78.8005
R5227 VDPWR.n29 VDPWR.t207 78.8005
R5228 VDPWR.n29 VDPWR.t425 78.8005
R5229 VDPWR.n2 VDPWR.t168 78.8005
R5230 VDPWR.n2 VDPWR.t31 78.8005
R5231 VDPWR.n21 VDPWR.t209 78.8005
R5232 VDPWR.n21 VDPWR.t103 78.8005
R5233 VDPWR.n19 VDPWR.t247 78.8005
R5234 VDPWR.n19 VDPWR.t195 78.8005
R5235 VDPWR.n17 VDPWR.t134 78.8005
R5236 VDPWR.n17 VDPWR.t119 78.8005
R5237 VDPWR.n4 VDPWR.t411 78.8005
R5238 VDPWR.n4 VDPWR.t5 78.8005
R5239 VDPWR.n9 VDPWR.t74 78.8005
R5240 VDPWR.n9 VDPWR.t221 78.8005
R5241 VDPWR.n7 VDPWR.t76 78.8005
R5242 VDPWR.n7 VDPWR.t372 78.8005
R5243 VDPWR.n6 VDPWR.t381 78.8005
R5244 VDPWR.n6 VDPWR.t23 78.8005
R5245 VDPWR.n194 VDPWR.n162 76.2865
R5246 VDPWR.t378 VDPWR.t192 76.1455
R5247 VDPWR.t389 VDPWR.t317 76.1455
R5248 VDPWR.n283 VDPWR.n282 72.1074
R5249 VDPWR.n366 VDPWR.n224 71.8576
R5250 VDPWR.n301 VDPWR.n300 71.0449
R5251 VDPWR.n493 VDPWR.n492 69.8479
R5252 VDPWR.n494 VDPWR.n493 69.8479
R5253 VDPWR.n472 VDPWR.n432 69.8479
R5254 VDPWR.n472 VDPWR.n433 69.8479
R5255 VDPWR.n292 VDPWR.n260 69.8479
R5256 VDPWR.n292 VDPWR.n259 69.8479
R5257 VDPWR.n299 VDPWR.n298 69.8479
R5258 VDPWR.n298 VDPWR.n297 69.8479
R5259 VDPWR.n311 VDPWR.n243 69.8479
R5260 VDPWR.n311 VDPWR.n242 69.8479
R5261 VDPWR.n292 VDPWR.n291 69.8479
R5262 VDPWR.n292 VDPWR.n258 69.8479
R5263 VDPWR.n311 VDPWR.n310 69.8479
R5264 VDPWR.n311 VDPWR.n241 69.8479
R5265 VDPWR.n280 VDPWR.n274 69.8479
R5266 VDPWR.n99 VDPWR.n98 69.8479
R5267 VDPWR.n99 VDPWR.n55 69.8479
R5268 VDPWR.n106 VDPWR.n105 69.8479
R5269 VDPWR.n107 VDPWR.n106 69.8479
R5270 VDPWR.n74 VDPWR.n68 69.8479
R5271 VDPWR.t192 VDPWR.t36 68.8936
R5272 VDPWR.n493 VDPWR.t389 68.8936
R5273 VDPWR.n48 VDPWR.n47 68.2005
R5274 VDPWR.n44 VDPWR.n43 68.2005
R5275 VDPWR.n28 VDPWR.n27 68.2005
R5276 VDPWR.n24 VDPWR.n23 68.2005
R5277 VDPWR.n16 VDPWR.n15 68.2005
R5278 VDPWR.n12 VDPWR.n11 68.2005
R5279 VDPWR.n610 VDPWR.n609 65.8183
R5280 VDPWR.n610 VDPWR.n594 65.8183
R5281 VDPWR.n593 VDPWR.n571 65.8183
R5282 VDPWR.n593 VDPWR.n572 65.8183
R5283 VDPWR.n328 VDPWR.n327 65.8183
R5284 VDPWR.n328 VDPWR.n237 65.8183
R5285 VDPWR.n344 VDPWR.n228 65.8183
R5286 VDPWR.n339 VDPWR.n228 65.8183
R5287 VDPWR.n368 VDPWR.n367 65.8183
R5288 VDPWR.n368 VDPWR.n359 65.8183
R5289 VDPWR.n383 VDPWR.n382 65.8183
R5290 VDPWR.n382 VDPWR.n374 65.8183
R5291 VDPWR.n398 VDPWR.n208 65.8183
R5292 VDPWR.n398 VDPWR.n207 65.8183
R5293 VDPWR.n413 VDPWR.n412 65.8183
R5294 VDPWR.n412 VDPWR.n404 65.8183
R5295 VDPWR.n317 VDPWR.n316 65.8183
R5296 VDPWR.n318 VDPWR.n317 65.8183
R5297 VDPWR.n334 VDPWR.n333 65.8183
R5298 VDPWR.n335 VDPWR.n334 65.8183
R5299 VDPWR.n358 VDPWR.n357 65.8183
R5300 VDPWR.n358 VDPWR.n229 65.8183
R5301 VDPWR.n382 VDPWR.n381 65.8183
R5302 VDPWR.n382 VDPWR.n369 65.8183
R5303 VDPWR.n398 VDPWR.n397 65.8183
R5304 VDPWR.n398 VDPWR.n206 65.8183
R5305 VDPWR.n412 VDPWR.n411 65.8183
R5306 VDPWR.n412 VDPWR.n399 65.8183
R5307 VDPWR.t348 VDPWR.t135 61.6417
R5308 VDPWR.t169 VDPWR.t60 61.6417
R5309 VDPWR.n195 VDPWR.t181 61.3458
R5310 VDPWR.n419 VDPWR.t426 58.8005
R5311 VDPWR.n418 VDPWR.t427 58.8005
R5312 VDPWR.n415 VDPWR.n203 58.0576
R5313 VDPWR.n415 VDPWR.n414 58.0576
R5314 VDPWR.n385 VDPWR.n225 58.0576
R5315 VDPWR.n385 VDPWR.n384 58.0576
R5316 VDPWR.n346 VDPWR.n336 58.0576
R5317 VDPWR.n346 VDPWR.n345 58.0576
R5318 VDPWR.n320 VDPWR.n319 58.0576
R5319 VDPWR.n326 VDPWR.n320 58.0576
R5320 VDPWR.t265 VDPWR.t412 57.5117
R5321 VDPWR.t269 VDPWR.t54 57.5117
R5322 VDPWR.t267 VDPWR.t382 57.5117
R5323 VDPWR.n304 VDPWR.n303 57.2449
R5324 VDPWR.n303 VDPWR.n253 57.2449
R5325 VDPWR.n285 VDPWR.n284 57.2449
R5326 VDPWR.n284 VDPWR.n270 57.2449
R5327 VDPWR.n459 VDPWR.n448 56.338
R5328 VDPWR.n352 VDPWR.n351 54.8576
R5329 VDPWR.n389 VDPWR.n212 54.4005
R5330 VDPWR.n223 VDPWR.n212 54.4005
R5331 VDPWR.n389 VDPWR.n388 54.4005
R5332 VDPWR.n388 VDPWR.n223 54.4005
R5333 VDPWR.n603 VDPWR.n594 53.3664
R5334 VDPWR.n609 VDPWR.n596 53.3664
R5335 VDPWR.n594 VDPWR.n570 53.3664
R5336 VDPWR.n574 VDPWR.n571 53.3664
R5337 VDPWR.n586 VDPWR.n572 53.3664
R5338 VDPWR.n587 VDPWR.n571 53.3664
R5339 VDPWR.n579 VDPWR.n572 53.3664
R5340 VDPWR.n404 VDPWR.n403 53.3664
R5341 VDPWR.n218 VDPWR.n207 53.3664
R5342 VDPWR.n374 VDPWR.n373 53.3664
R5343 VDPWR.n327 VDPWR.n238 53.3664
R5344 VDPWR.n322 VDPWR.n237 53.3664
R5345 VDPWR.n344 VDPWR.n343 53.3664
R5346 VDPWR.n339 VDPWR.n338 53.3664
R5347 VDPWR.n367 VDPWR.n360 53.3664
R5348 VDPWR.n362 VDPWR.n359 53.3664
R5349 VDPWR.n383 VDPWR.n227 53.3664
R5350 VDPWR.n217 VDPWR.n208 53.3664
R5351 VDPWR.n413 VDPWR.n205 53.3664
R5352 VDPWR.n316 VDPWR.n312 53.3664
R5353 VDPWR.n318 VDPWR.n240 53.3664
R5354 VDPWR.n333 VDPWR.n329 53.3664
R5355 VDPWR.n335 VDPWR.n236 53.3664
R5356 VDPWR.n357 VDPWR.n230 53.3664
R5357 VDPWR.n353 VDPWR.n229 53.3664
R5358 VDPWR.n381 VDPWR.n375 53.3664
R5359 VDPWR.n377 VDPWR.n369 53.3664
R5360 VDPWR.n397 VDPWR.n209 53.3664
R5361 VDPWR.n392 VDPWR.n206 53.3664
R5362 VDPWR.n411 VDPWR.n405 53.3664
R5363 VDPWR.n407 VDPWR.n399 53.3664
R5364 VDPWR.n477 VDPWR.n428 50.9005
R5365 VDPWR.t88 VDPWR.n481 50.7639
R5366 VDPWR.n429 VDPWR.t29 49.2505
R5367 VDPWR.n429 VDPWR.t193 49.2505
R5368 VDPWR.n427 VDPWR.t243 49.2505
R5369 VDPWR.n427 VDPWR.t314 49.2505
R5370 VDPWR.t349 VDPWR.n430 49.2505
R5371 VDPWR.n430 VDPWR.t370 49.2505
R5372 VDPWR.n439 VDPWR.t13 49.2505
R5373 VDPWR.n439 VDPWR.t8 49.2505
R5374 VDPWR.n444 VDPWR.t17 49.2505
R5375 VDPWR.n444 VDPWR.t362 49.2505
R5376 VDPWR.t352 VDPWR.n440 49.2505
R5377 VDPWR.n440 VDPWR.t114 49.2505
R5378 VDPWR.n418 VDPWR.t431 49.1638
R5379 VDPWR.n420 VDPWR.t433 48.5162
R5380 VDPWR.n494 VDPWR.n426 45.3071
R5381 VDPWR.n492 VDPWR.n483 45.3071
R5382 VDPWR.n434 VDPWR.n432 45.3071
R5383 VDPWR.n465 VDPWR.n433 45.3071
R5384 VDPWR.n466 VDPWR.n432 45.3071
R5385 VDPWR.n250 VDPWR.n242 45.3071
R5386 VDPWR.n267 VDPWR.n259 45.3071
R5387 VDPWR.n268 VDPWR.n260 45.3071
R5388 VDPWR.n299 VDPWR.n257 45.3071
R5389 VDPWR.n297 VDPWR.n296 45.3071
R5390 VDPWR.n251 VDPWR.n243 45.3071
R5391 VDPWR.n291 VDPWR.n261 45.3071
R5392 VDPWR.n286 VDPWR.n258 45.3071
R5393 VDPWR.n310 VDPWR.n244 45.3071
R5394 VDPWR.n305 VDPWR.n241 45.3071
R5395 VDPWR.n274 VDPWR.n273 45.3071
R5396 VDPWR.n275 VDPWR.n274 45.3071
R5397 VDPWR.n98 VDPWR.n56 45.3071
R5398 VDPWR.n85 VDPWR.n55 45.3071
R5399 VDPWR.n105 VDPWR.n100 45.3071
R5400 VDPWR.n107 VDPWR.n54 45.3071
R5401 VDPWR.n68 VDPWR.n67 45.3071
R5402 VDPWR.n72 VDPWR.n68 45.3071
R5403 VDPWR.t373 VDPWR.t67 39.886
R5404 VDPWR.n537 VDPWR.t150 39.4005
R5405 VDPWR.n537 VDPWR.t278 39.4005
R5406 VDPWR.n535 VDPWR.t1 39.4005
R5407 VDPWR.n535 VDPWR.t180 39.4005
R5408 VDPWR.n533 VDPWR.t274 39.4005
R5409 VDPWR.n533 VDPWR.t183 39.4005
R5410 VDPWR.n531 VDPWR.t95 39.4005
R5411 VDPWR.n531 VDPWR.t282 39.4005
R5412 VDPWR.n529 VDPWR.t53 39.4005
R5413 VDPWR.n529 VDPWR.t241 39.4005
R5414 VDPWR.n527 VDPWR.t276 39.4005
R5415 VDPWR.n527 VDPWR.t97 39.4005
R5416 VDPWR.n525 VDPWR.t217 39.4005
R5417 VDPWR.n525 VDPWR.t272 39.4005
R5418 VDPWR.n523 VDPWR.t286 39.4005
R5419 VDPWR.n523 VDPWR.t152 39.4005
R5420 VDPWR.n519 VDPWR.t280 39.4005
R5421 VDPWR.n519 VDPWR.t249 39.4005
R5422 VDPWR.n517 VDPWR.t21 39.4005
R5423 VDPWR.n517 VDPWR.t262 39.4005
R5424 VDPWR.n515 VDPWR.t288 39.4005
R5425 VDPWR.n515 VDPWR.t292 39.4005
R5426 VDPWR.n513 VDPWR.t256 39.4005
R5427 VDPWR.n513 VDPWR.t252 39.4005
R5428 VDPWR.n511 VDPWR.t365 39.4005
R5429 VDPWR.n511 VDPWR.t254 39.4005
R5430 VDPWR.n509 VDPWR.t141 39.4005
R5431 VDPWR.n509 VDPWR.t70 39.4005
R5432 VDPWR.n507 VDPWR.t260 39.4005
R5433 VDPWR.n507 VDPWR.t66 39.4005
R5434 VDPWR.n505 VDPWR.t185 39.4005
R5435 VDPWR.n505 VDPWR.t264 39.4005
R5436 VDPWR.n503 VDPWR.t127 39.4005
R5437 VDPWR.n503 VDPWR.t290 39.4005
R5438 VDPWR.n499 VDPWR.t258 39.4005
R5439 VDPWR.n499 VDPWR.t51 39.4005
R5440 VDPWR.n660 VDPWR.t223 39.4005
R5441 VDPWR.n660 VDPWR.t201 39.4005
R5442 VDPWR.n658 VDPWR.t27 39.4005
R5443 VDPWR.n658 VDPWR.t375 39.4005
R5444 VDPWR.n656 VDPWR.t156 39.4005
R5445 VDPWR.n656 VDPWR.t129 39.4005
R5446 VDPWR.n654 VDPWR.t25 39.4005
R5447 VDPWR.n654 VDPWR.t125 39.4005
R5448 VDPWR.n649 VDPWR.t391 39.4005
R5449 VDPWR.n649 VDPWR.t407 39.4005
R5450 VDPWR.n647 VDPWR.t205 39.4005
R5451 VDPWR.n647 VDPWR.t80 39.4005
R5452 VDPWR.n645 VDPWR.t393 39.4005
R5453 VDPWR.n645 VDPWR.t116 39.4005
R5454 VDPWR.n643 VDPWR.t10 39.4005
R5455 VDPWR.n643 VDPWR.t163 39.4005
R5456 VDPWR.n641 VDPWR.t64 39.4005
R5457 VDPWR.n641 VDPWR.t165 39.4005
R5458 VDPWR.n636 VDPWR.t78 39.4005
R5459 VDPWR.n636 VDPWR.t215 39.4005
R5460 VDPWR.n197 VDPWR.n196 37.0005
R5461 VDPWR.n163 VDPWR.n162 37.0005
R5462 VDPWR.n473 VDPWR.t345 36.26
R5463 VDPWR.t135 VDPWR.t369 32.6341
R5464 VDPWR.t394 VDPWR.t169 32.6341
R5465 VDPWR.n446 VDPWR.n445 30.754
R5466 VDPWR.n442 VDPWR.n441 30.186
R5467 VDPWR.n480 VDPWR.n479 30.18
R5468 VDPWR.n475 VDPWR.n474 29.7151
R5469 VDPWR.t36 VDPWR.t242 25.3822
R5470 VDPWR.t313 VDPWR.t130 25.3822
R5471 VDPWR.n246 VDPWR.t99 24.6255
R5472 VDPWR.n245 VDPWR.t203 24.6255
R5473 VDPWR.n255 VDPWR.t230 24.6255
R5474 VDPWR.n263 VDPWR.t202 24.6255
R5475 VDPWR.n262 VDPWR.t187 24.6255
R5476 VDPWR.n271 VDPWR.t409 24.6255
R5477 VDPWR.n49 VDPWR.t154 24.6255
R5478 VDPWR.n49 VDPWR.t304 24.6255
R5479 VDPWR.n91 VDPWR.t235 24.6255
R5480 VDPWR.n91 VDPWR.t237 24.6255
R5481 VDPWR.t343 VDPWR.n94 24.6255
R5482 VDPWR.n94 VDPWR.t19 24.6255
R5483 VDPWR.n82 VDPWR.t232 24.6255
R5484 VDPWR.n82 VDPWR.t358 24.6255
R5485 VDPWR.n80 VDPWR.t239 24.6255
R5486 VDPWR.n80 VDPWR.t191 24.6255
R5487 VDPWR.n78 VDPWR.t308 24.6255
R5488 VDPWR.n78 VDPWR.t226 24.6255
R5489 VDPWR.t308 VDPWR.n77 24.6255
R5490 VDPWR.n53 VDPWR.t305 24.6255
R5491 VDPWR.n95 VDPWR.t343 24.6255
R5492 VDPWR.n59 VDPWR.t359 24.6255
R5493 VDPWR.n613 VDPWR.n612 22.8576
R5494 VDPWR.n582 VDPWR.n559 22.8576
R5495 VDPWR.n134 VDPWR.n133 21.6365
R5496 VDPWR.n132 VDPWR.n129 21.6365
R5497 VDPWR.n128 VDPWR.n127 21.6365
R5498 VDPWR.n120 VDPWR.n118 21.6365
R5499 VDPWR.n156 VDPWR.n155 21.6365
R5500 VDPWR.n154 VDPWR.n151 21.6365
R5501 VDPWR.n150 VDPWR.n149 21.6365
R5502 VDPWR.n142 VDPWR.n140 21.6365
R5503 VDPWR.n187 VDPWR.n186 21.6365
R5504 VDPWR.n185 VDPWR.n182 21.6365
R5505 VDPWR.n181 VDPWR.n180 21.6365
R5506 VDPWR.n173 VDPWR.n171 21.6365
R5507 VDPWR.n131 VDPWR.n114 21.3338
R5508 VDPWR.n125 VDPWR.n116 21.3338
R5509 VDPWR.n125 VDPWR.n117 21.3338
R5510 VDPWR.n121 VDPWR.n117 21.3338
R5511 VDPWR.n153 VDPWR.n136 21.3338
R5512 VDPWR.n147 VDPWR.n138 21.3338
R5513 VDPWR.n147 VDPWR.n139 21.3338
R5514 VDPWR.n143 VDPWR.n139 21.3338
R5515 VDPWR.n184 VDPWR.n167 21.3338
R5516 VDPWR.n178 VDPWR.n169 21.3338
R5517 VDPWR.n178 VDPWR.n170 21.3338
R5518 VDPWR.n174 VDPWR.n170 21.3338
R5519 VDPWR.n453 VDPWR.t379 19.7005
R5520 VDPWR.n453 VDPWR.t37 19.7005
R5521 VDPWR.n422 VDPWR.t170 19.7005
R5522 VDPWR.n422 VDPWR.t318 19.7005
R5523 VDPWR.n449 VDPWR.t68 19.7005
R5524 VDPWR.n449 VDPWR.t87 19.7005
R5525 VDPWR.n451 VDPWR.t131 19.7005
R5526 VDPWR.n451 VDPWR.t89 19.7005
R5527 VDPWR.n457 VDPWR.t346 19.7005
R5528 VDPWR.n457 VDPWR.t136 19.7005
R5529 VDPWR.t346 VDPWR.n435 19.7005
R5530 VDPWR.n490 VDPWR.t319 19.7005
R5531 VDPWR.n421 VDPWR.t423 18.7777
R5532 VDPWR.t28 VDPWR.t378 18.1303
R5533 VDPWR.t317 VDPWR.t157 18.1303
R5534 VDPWR.n479 VDPWR.n478 16.0005
R5535 VDPWR.n476 VDPWR.n475 16.0005
R5536 VDPWR.n447 VDPWR.n446 16.0005
R5537 VDPWR.n443 VDPWR.n442 16.0005
R5538 VDPWR.n496 VDPWR.n495 15.6449
R5539 VDPWR.n497 VDPWR.n496 14.0505
R5540 VDPWR.n284 VDPWR.n283 13.8005
R5541 VDPWR.n303 VDPWR.n302 13.8005
R5542 VDPWR.n320 VDPWR.n234 13.8005
R5543 VDPWR.n347 VDPWR.n346 13.8005
R5544 VDPWR.n386 VDPWR.n385 13.8005
R5545 VDPWR.n388 VDPWR.n387 13.8005
R5546 VDPWR.n212 VDPWR.n202 13.8005
R5547 VDPWR.n416 VDPWR.n415 13.8005
R5548 VDPWR.n567 VDPWR.t148 13.1338
R5549 VDPWR.n567 VDPWR.t387 13.1338
R5550 VDPWR.n566 VDPWR.t211 13.1338
R5551 VDPWR.n566 VDPWR.t175 13.1338
R5552 VDPWR.n565 VDPWR.t417 13.1338
R5553 VDPWR.n565 VDPWR.t419 13.1338
R5554 VDPWR.n564 VDPWR.t144 13.1338
R5555 VDPWR.n564 VDPWR.t139 13.1338
R5556 VDPWR.n563 VDPWR.t146 13.1338
R5557 VDPWR.n563 VDPWR.t213 13.1338
R5558 VDPWR.n562 VDPWR.t111 13.1338
R5559 VDPWR.n562 VDPWR.t198 13.1338
R5560 VDPWR.n561 VDPWR.t367 13.1338
R5561 VDPWR.n561 VDPWR.t401 13.1338
R5562 VDPWR.n560 VDPWR.t91 13.1338
R5563 VDPWR.n560 VDPWR.t93 13.1338
R5564 VDPWR.n351 VDPWR.n232 12.8005
R5565 VDPWR.n317 VDPWR.t108 11.4924
R5566 VDPWR.n328 VDPWR.t420 11.4924
R5567 VDPWR.n334 VDPWR.t414 11.4924
R5568 VDPWR.t160 VDPWR.n228 11.4924
R5569 VDPWR.t176 VDPWR.n358 11.4924
R5570 VDPWR.n614 VDPWR.n613 11.0575
R5571 VDPWR.t86 VDPWR.t85 10.8784
R5572 VDPWR.n622 VDPWR.n559 10.87
R5573 VDPWR.n129 VDPWR.n128 10.1932
R5574 VDPWR.n151 VDPWR.n150 10.1932
R5575 VDPWR.n182 VDPWR.n181 10.1932
R5576 VDPWR.n164 VDPWR.n158 9.6005
R5577 VDPWR.n545 VDPWR.n521 9.50883
R5578 VDPWR.n555 VDPWR.n501 9.50883
R5579 VDPWR.n591 VDPWR.n590 9.50883
R5580 VDPWR.n583 VDPWR.n582 9.50883
R5581 VDPWR.n608 VDPWR.n597 9.50883
R5582 VDPWR.n612 VDPWR.n569 9.50883
R5583 VDPWR.n632 VDPWR.n624 9.50883
R5584 VDPWR.n495 VDPWR.n424 9.45675
R5585 VDPWR.n487 VDPWR.n424 9.3005
R5586 VDPWR.n488 VDPWR.n486 9.3005
R5587 VDPWR.n464 VDPWR.n437 9.3005
R5588 VDPWR.n468 VDPWR.n467 9.3005
R5589 VDPWR.n462 VDPWR.n461 9.3005
R5590 VDPWR.n545 VDPWR.n544 9.3005
R5591 VDPWR.n555 VDPWR.n554 9.3005
R5592 VDPWR.n601 VDPWR.n569 9.3005
R5593 VDPWR.n604 VDPWR.n600 9.3005
R5594 VDPWR.n605 VDPWR.n599 9.3005
R5595 VDPWR.n598 VDPWR.n597 9.3005
R5596 VDPWR.n583 VDPWR.n580 9.3005
R5597 VDPWR.n585 VDPWR.n584 9.3005
R5598 VDPWR.n588 VDPWR.n576 9.3005
R5599 VDPWR.n590 VDPWR.n589 9.3005
R5600 VDPWR.n632 VDPWR.n631 9.3005
R5601 VDPWR.n351 VDPWR.n350 9.3005
R5602 VDPWR.n233 VDPWR.n232 9.3005
R5603 VDPWR.n122 VDPWR.n121 9.3005
R5604 VDPWR.n123 VDPWR.n117 9.3005
R5605 VDPWR.n125 VDPWR.n124 9.3005
R5606 VDPWR.n116 VDPWR.n115 9.3005
R5607 VDPWR.n131 VDPWR.n130 9.3005
R5608 VDPWR.n114 VDPWR.n113 9.3005
R5609 VDPWR.n144 VDPWR.n143 9.3005
R5610 VDPWR.n145 VDPWR.n139 9.3005
R5611 VDPWR.n147 VDPWR.n146 9.3005
R5612 VDPWR.n138 VDPWR.n137 9.3005
R5613 VDPWR.n153 VDPWR.n152 9.3005
R5614 VDPWR.n136 VDPWR.n135 9.3005
R5615 VDPWR.n175 VDPWR.n174 9.3005
R5616 VDPWR.n176 VDPWR.n170 9.3005
R5617 VDPWR.n178 VDPWR.n177 9.3005
R5618 VDPWR.n169 VDPWR.n168 9.3005
R5619 VDPWR.n184 VDPWR.n183 9.3005
R5620 VDPWR.n167 VDPWR.n166 9.3005
R5621 VDPWR.n188 VDPWR.n165 9.3005
R5622 VDPWR.n158 VDPWR.n157 9.3005
R5623 VDPWR.n199 VDPWR.n198 9.3005
R5624 VDPWR.n191 VDPWR.n190 9.3005
R5625 VDPWR.n52 VDPWR.n51 9.3005
R5626 VDPWR.n109 VDPWR.n108 9.3005
R5627 VDPWR.n71 VDPWR.n70 9.3005
R5628 VDPWR.n69 VDPWR.n64 9.3005
R5629 VDPWR.n605 VDPWR.n598 9.14336
R5630 VDPWR.n605 VDPWR.n604 9.14336
R5631 VDPWR.n604 VDPWR.n601 9.14336
R5632 VDPWR.n589 VDPWR.n588 9.14336
R5633 VDPWR.n588 VDPWR.n585 9.14336
R5634 VDPWR.n585 VDPWR.n580 9.14336
R5635 VDPWR.n354 VDPWR.n231 9.14336
R5636 VDPWR.n408 VDPWR.n406 9.14336
R5637 VDPWR.n402 VDPWR.n401 9.14336
R5638 VDPWR.n378 VDPWR.n376 9.14336
R5639 VDPWR.n372 VDPWR.n371 9.14336
R5640 VDPWR.n363 VDPWR.n361 9.14336
R5641 VDPWR.n331 VDPWR.n330 9.14336
R5642 VDPWR.n342 VDPWR.n341 9.14336
R5643 VDPWR.n314 VDPWR.n313 9.14336
R5644 VDPWR.n323 VDPWR.n321 9.14336
R5645 VDPWR.n133 VDPWR.n114 8.68224
R5646 VDPWR.n132 VDPWR.n131 8.68224
R5647 VDPWR.n127 VDPWR.n116 8.68224
R5648 VDPWR.n121 VDPWR.n120 8.68224
R5649 VDPWR.n155 VDPWR.n136 8.68224
R5650 VDPWR.n154 VDPWR.n153 8.68224
R5651 VDPWR.n149 VDPWR.n138 8.68224
R5652 VDPWR.n143 VDPWR.n142 8.68224
R5653 VDPWR.n186 VDPWR.n167 8.68224
R5654 VDPWR.n185 VDPWR.n184 8.68224
R5655 VDPWR.n180 VDPWR.n169 8.68224
R5656 VDPWR.n174 VDPWR.n173 8.68224
R5657 VDPWR.t38 VDPWR.t2 7.66179
R5658 VDPWR.n472 VDPWR.n431 7.25241
R5659 VDPWR.n488 VDPWR.n487 7.11161
R5660 VDPWR.n467 VDPWR.n464 7.11161
R5661 VDPWR.n309 VDPWR.n308 7.11161
R5662 VDPWR.n306 VDPWR.n304 7.11161
R5663 VDPWR.n253 VDPWR.n252 7.11161
R5664 VDPWR.n249 VDPWR.n248 7.11161
R5665 VDPWR.n300 VDPWR.n256 7.11161
R5666 VDPWR.n295 VDPWR.n293 7.11161
R5667 VDPWR.n290 VDPWR.n289 7.11161
R5668 VDPWR.n287 VDPWR.n285 7.11161
R5669 VDPWR.n270 VDPWR.n269 7.11161
R5670 VDPWR.n266 VDPWR.n265 7.11161
R5671 VDPWR.n282 VDPWR.n272 7.11161
R5672 VDPWR.n278 VDPWR.n277 7.11161
R5673 VDPWR.n108 VDPWR.n52 7.11161
R5674 VDPWR.n71 VDPWR.n64 7.11161
R5675 VDPWR.n681 VDPWR.n680 6.74656
R5676 VDPWR.n393 VDPWR.n211 5.81868
R5677 VDPWR.n219 VDPWR.n214 5.81868
R5678 VDPWR.n190 VDPWR.n189 5.46925
R5679 VDPWR.n608 VDPWR.n607 5.33286
R5680 VDPWR.n612 VDPWR.n568 5.33286
R5681 VDPWR.n591 VDPWR.n575 5.33286
R5682 VDPWR.n582 VDPWR.n581 5.33286
R5683 VDPWR.n355 VDPWR.n352 5.33286
R5684 VDPWR.n409 VDPWR.n203 5.33286
R5685 VDPWR.n414 VDPWR.n204 5.33286
R5686 VDPWR.n379 VDPWR.n225 5.33286
R5687 VDPWR.n384 VDPWR.n226 5.33286
R5688 VDPWR.n366 VDPWR.n365 5.33286
R5689 VDPWR.n336 VDPWR.n235 5.33286
R5690 VDPWR.n345 VDPWR.n337 5.33286
R5691 VDPWR.n319 VDPWR.n239 5.33286
R5692 VDPWR.n326 VDPWR.n325 5.33286
R5693 VDPWR.n684 VDPWR.n48 5.13102
R5694 VDPWR.n682 VDPWR.n416 5.04739
R5695 VDPWR.n79 VDPWR.n62 5.01612
R5696 VDPWR.n662 VDPWR.n661 4.84425
R5697 VDPWR.n90 VDPWR.n89 4.81523
R5698 VDPWR.n460 VDPWR.n459 4.7505
R5699 VDPWR.n664 VDPWR.n663 4.73979
R5700 VDPWR.n668 VDPWR.n651 4.73979
R5701 VDPWR.n674 VDPWR.n673 4.73979
R5702 VDPWR.n678 VDPWR.n638 4.73979
R5703 VDPWR.n111 VDPWR.n110 4.67238
R5704 VDPWR.n200 VDPWR.n199 4.65675
R5705 VDPWR.n157 VDPWR.n112 4.65675
R5706 VDPWR.n189 VDPWR.n188 4.65675
R5707 VDPWR.n663 VDPWR.n652 4.6505
R5708 VDPWR.n668 VDPWR.n667 4.6505
R5709 VDPWR.n673 VDPWR.n639 4.6505
R5710 VDPWR.n678 VDPWR.n677 4.6505
R5711 VDPWR.n653 VDPWR.n652 4.54311
R5712 VDPWR.n664 VDPWR.n653 4.54311
R5713 VDPWR.n640 VDPWR.n639 4.54311
R5714 VDPWR.n674 VDPWR.n640 4.54311
R5715 VDPWR.n455 VDPWR.n454 4.5005
R5716 VDPWR.n456 VDPWR.n428 4.5005
R5717 VDPWR.n680 VDPWR.n679 4.5005
R5718 VDPWR.n672 VDPWR.n671 4.5005
R5719 VDPWR.n670 VDPWR.n669 4.5005
R5720 VDPWR.n350 VDPWR.n349 4.5005
R5721 VDPWR.n348 VDPWR.n233 4.5005
R5722 VDPWR.n544 VDPWR.n543 4.48641
R5723 VDPWR.n543 VDPWR.n521 4.48641
R5724 VDPWR.n554 VDPWR.n553 4.48641
R5725 VDPWR.n553 VDPWR.n501 4.48641
R5726 VDPWR.n631 VDPWR.n630 4.48641
R5727 VDPWR.n630 VDPWR.n624 4.48641
R5728 VDPWR.n667 VDPWR.n666 4.48641
R5729 VDPWR.n666 VDPWR.n651 4.48641
R5730 VDPWR.n677 VDPWR.n676 4.48641
R5731 VDPWR.n676 VDPWR.n638 4.48641
R5732 VDPWR.n682 VDPWR.n681 4.17751
R5733 VDPWR.n683 VDPWR.n201 4.12598
R5734 VDPWR.n201 VDPWR.n200 3.83321
R5735 VDPWR.n498 VDPWR.n497 3.82369
R5736 VDPWR.n607 VDPWR.n598 3.75335
R5737 VDPWR.n601 VDPWR.n568 3.75335
R5738 VDPWR.n589 VDPWR.n575 3.75335
R5739 VDPWR.n581 VDPWR.n580 3.75335
R5740 VDPWR.n356 VDPWR.n231 3.75335
R5741 VDPWR.n355 VDPWR.n354 3.75335
R5742 VDPWR.n410 VDPWR.n406 3.75335
R5743 VDPWR.n409 VDPWR.n408 3.75335
R5744 VDPWR.n401 VDPWR.n204 3.75335
R5745 VDPWR.n402 VDPWR.n400 3.75335
R5746 VDPWR.n380 VDPWR.n376 3.75335
R5747 VDPWR.n379 VDPWR.n378 3.75335
R5748 VDPWR.n371 VDPWR.n226 3.75335
R5749 VDPWR.n372 VDPWR.n370 3.75335
R5750 VDPWR.n365 VDPWR.n361 3.75335
R5751 VDPWR.n364 VDPWR.n363 3.75335
R5752 VDPWR.n332 VDPWR.n331 3.75335
R5753 VDPWR.n330 VDPWR.n235 3.75335
R5754 VDPWR.n342 VDPWR.n337 3.75335
R5755 VDPWR.n341 VDPWR.n340 3.75335
R5756 VDPWR.n315 VDPWR.n314 3.75335
R5757 VDPWR.n313 VDPWR.n239 3.75335
R5758 VDPWR.n325 VDPWR.n321 3.75335
R5759 VDPWR.n324 VDPWR.n323 3.75335
R5760 VDPWR.n486 VDPWR.n484 3.55702
R5761 VDPWR.n469 VDPWR.n468 3.55702
R5762 VDPWR.n103 VDPWR.n51 3.55702
R5763 VDPWR.n70 VDPWR.n65 3.55702
R5764 VDPWR.n489 VDPWR.n485 3.53508
R5765 VDPWR.n487 VDPWR.n425 3.53508
R5766 VDPWR.n489 VDPWR.n488 3.53508
R5767 VDPWR.n495 VDPWR.n425 3.53508
R5768 VDPWR.n438 VDPWR.n436 3.53508
R5769 VDPWR.n464 VDPWR.n463 3.53508
R5770 VDPWR.n467 VDPWR.n438 3.53508
R5771 VDPWR.n463 VDPWR.n462 3.53508
R5772 VDPWR.n308 VDPWR.n307 3.53508
R5773 VDPWR.n307 VDPWR.n306 3.53508
R5774 VDPWR.n252 VDPWR.n247 3.53508
R5775 VDPWR.n249 VDPWR.n247 3.53508
R5776 VDPWR.n294 VDPWR.n256 3.53508
R5777 VDPWR.n295 VDPWR.n294 3.53508
R5778 VDPWR.n289 VDPWR.n288 3.53508
R5779 VDPWR.n288 VDPWR.n287 3.53508
R5780 VDPWR.n269 VDPWR.n264 3.53508
R5781 VDPWR.n266 VDPWR.n264 3.53508
R5782 VDPWR.n276 VDPWR.n272 3.53508
R5783 VDPWR.n277 VDPWR.n276 3.53508
R5784 VDPWR.n102 VDPWR.n101 3.53508
R5785 VDPWR.n101 VDPWR.n52 3.53508
R5786 VDPWR.n66 VDPWR.n63 3.53508
R5787 VDPWR.n71 VDPWR.n63 3.53508
R5788 VDPWR.n627 VDPWR.n626 3.46433
R5789 VDPWR.n540 VDPWR.n539 3.41464
R5790 VDPWR.n550 VDPWR.n549 3.41464
R5791 VDPWR.n396 VDPWR.n395 3.40194
R5792 VDPWR.n394 VDPWR.n390 3.40194
R5793 VDPWR.n222 VDPWR.n221 3.40194
R5794 VDPWR.n220 VDPWR.n215 3.40194
R5795 VDPWR.n97 VDPWR.n58 3.14514
R5796 VDPWR.n541 VDPWR.n540 3.11118
R5797 VDPWR.n551 VDPWR.n550 3.11118
R5798 VDPWR.n87 VDPWR.n86 3.1005
R5799 VDPWR.n60 VDPWR.n58 3.1005
R5800 VDPWR.n89 VDPWR.n88 3.1005
R5801 VDPWR.n540 VDPWR.n522 3.04304
R5802 VDPWR.n550 VDPWR.n502 3.04304
R5803 VDPWR.n628 VDPWR.n627 2.96855
R5804 VDPWR.n627 VDPWR.n625 2.90353
R5805 VDPWR.n491 VDPWR.n484 2.60059
R5806 VDPWR.n470 VDPWR.n469 2.60059
R5807 VDPWR.n104 VDPWR.n103 2.60059
R5808 VDPWR.n76 VDPWR.n65 2.60059
R5809 VDPWR.n485 VDPWR.n484 2.55763
R5810 VDPWR.n469 VDPWR.n436 2.55763
R5811 VDPWR.n103 VDPWR.n102 2.55763
R5812 VDPWR.n66 VDPWR.n65 2.55763
R5813 VDPWR.n395 VDPWR.n211 2.39444
R5814 VDPWR.n394 VDPWR.n393 2.39444
R5815 VDPWR.n221 VDPWR.n214 2.39444
R5816 VDPWR.n220 VDPWR.n219 2.39444
R5817 VDPWR.n421 VDPWR.n420 2.35874
R5818 VDPWR.n390 VDPWR.n389 2.32777
R5819 VDPWR.n223 VDPWR.n222 2.32777
R5820 VDPWR.n96 VDPWR.n60 2.27782
R5821 VDPWR.n84 VDPWR.n60 2.27782
R5822 VDPWR.n88 VDPWR.n61 2.27782
R5823 VDPWR.n86 VDPWR.n84 2.27782
R5824 VDPWR.n97 VDPWR.n96 2.27782
R5825 VDPWR.n86 VDPWR.n61 2.27782
R5826 VDPWR.n201 VDPWR.n111 2.13269
R5827 VDPWR.n635 VDPWR.n634 1.97722
R5828 VDPWR.n558 VDPWR.n557 1.9616
R5829 VDPWR.n626 VDPWR.n623 1.94497
R5830 VDPWR.n634 VDPWR.n633 1.94497
R5831 VDPWR.n539 VDPWR.n538 1.90331
R5832 VDPWR.n547 VDPWR.n546 1.77831
R5833 VDPWR.n549 VDPWR.n548 1.77831
R5834 VDPWR.n557 VDPWR.n556 1.77831
R5835 VDPWR.n387 VDPWR.n386 1.15675
R5836 VDPWR.n416 VDPWR.n202 1.15675
R5837 VDPWR.n43 VDPWR.n42 1.10988
R5838 VDPWR.n40 VDPWR.n1 1.04738
R5839 VDPWR.n30 VDPWR.n28 0.96925
R5840 VDPWR.n11 VDPWR.n10 0.938
R5841 VDPWR.n18 VDPWR.n16 0.938
R5842 VDPWR.n23 VDPWR.n22 0.938
R5843 VDPWR.n671 VDPWR.n670 0.90675
R5844 VDPWR.n42 VDPWR.n40 0.891125
R5845 VDPWR.n189 VDPWR.n112 0.813
R5846 VDPWR.n200 VDPWR.n112 0.813
R5847 VDPWR.n192 VDPWR.n191 0.8005
R5848 VDPWR.n419 VDPWR.n418 0.75233
R5849 VDPWR.n33 VDPWR.n32 0.734875
R5850 VDPWR.n302 VDPWR.n234 0.688
R5851 VDPWR.n81 VDPWR.n79 0.688
R5852 VDPWR.n83 VDPWR.n81 0.688
R5853 VDPWR.n93 VDPWR.n92 0.688
R5854 VDPWR.n92 VDPWR.n50 0.688
R5855 VDPWR.n32 VDPWR.n30 0.688
R5856 VDPWR.n38 VDPWR.n36 0.688
R5857 VDPWR.n43 VDPWR.n38 0.672375
R5858 VDPWR.n48 VDPWR.n1 0.65675
R5859 VDPWR.n420 VDPWR.n419 0.648711
R5860 VDPWR.n455 VDPWR.n452 0.6255
R5861 VDPWR.n452 VDPWR.n450 0.6255
R5862 VDPWR.n450 VDPWR.n423 0.6255
R5863 VDPWR.n302 VDPWR.n301 0.609875
R5864 VDPWR.n10 VDPWR.n5 0.563
R5865 VDPWR.n20 VDPWR.n18 0.563
R5866 VDPWR.n22 VDPWR.n3 0.563
R5867 VDPWR.n11 VDPWR.n8 0.53175
R5868 VDPWR.n16 VDPWR.n5 0.53175
R5869 VDPWR.n23 VDPWR.n20 0.53175
R5870 VDPWR.n28 VDPWR.n3 0.53175
R5871 VDPWR.n347 VDPWR.n234 0.516125
R5872 VDPWR.n458 VDPWR.n456 0.5005
R5873 VDPWR.n90 VDPWR.n83 0.5005
R5874 VDPWR.n93 VDPWR.n90 0.5005
R5875 VDPWR.t181 VDPWR.t265 0.426509
R5876 VDPWR.t224 VDPWR.t269 0.426509
R5877 VDPWR.t166 VDPWR.t267 0.426509
R5878 VDPWR.n386 VDPWR.n224 0.391125
R5879 VDPWR.n36 VDPWR.n34 0.391125
R5880 VDPWR.n680 VDPWR.n637 0.34425
R5881 VDPWR.n642 VDPWR.n637 0.34425
R5882 VDPWR.n644 VDPWR.n642 0.34425
R5883 VDPWR.n646 VDPWR.n644 0.34425
R5884 VDPWR.n648 VDPWR.n646 0.34425
R5885 VDPWR.n671 VDPWR.n648 0.34425
R5886 VDPWR.n670 VDPWR.n650 0.34425
R5887 VDPWR.n655 VDPWR.n650 0.34425
R5888 VDPWR.n657 VDPWR.n655 0.34425
R5889 VDPWR.n659 VDPWR.n657 0.34425
R5890 VDPWR.n661 VDPWR.n659 0.34425
R5891 VDPWR.n111 VDPWR.n50 0.34425
R5892 VDPWR.n34 VDPWR.n33 0.34425
R5893 VDPWR.n548 VDPWR.n547 0.333833
R5894 VDPWR.n623 VDPWR.n622 0.328625
R5895 VDPWR.n301 VDPWR.n254 0.328625
R5896 VDPWR.n348 VDPWR.n347 0.328625
R5897 VDPWR VDPWR.n684 0.320874
R5898 VDPWR.n459 VDPWR.n458 0.313
R5899 VDPWR.n497 VDPWR.n423 0.313
R5900 VDPWR.n349 VDPWR.n224 0.297375
R5901 VDPWR.n635 VDPWR.n558 0.285347
R5902 VDPWR.n283 VDPWR.n254 0.28175
R5903 VDPWR.n546 VDPWR.n545 0.2505
R5904 VDPWR.n556 VDPWR.n555 0.2505
R5905 VDPWR.n387 VDPWR.n202 0.2505
R5906 VDPWR.n199 VDPWR.n134 0.2505
R5907 VDPWR.n157 VDPWR.n156 0.2505
R5908 VDPWR.n188 VDPWR.n187 0.2505
R5909 VDPWR.n633 VDPWR.n632 0.229667
R5910 VDPWR.n634 VDPWR.n623 0.229667
R5911 VDPWR.n684 VDPWR.n683 0.227655
R5912 VDPWR.n590 VDPWR.n576 0.208833
R5913 VDPWR.n584 VDPWR.n576 0.208833
R5914 VDPWR.n584 VDPWR.n583 0.208833
R5915 VDPWR.n599 VDPWR.n597 0.208833
R5916 VDPWR.n600 VDPWR.n599 0.208833
R5917 VDPWR.n600 VDPWR.n569 0.208833
R5918 VDPWR.n128 VDPWR.n115 0.208833
R5919 VDPWR.n124 VDPWR.n115 0.208833
R5920 VDPWR.n124 VDPWR.n123 0.208833
R5921 VDPWR.n123 VDPWR.n122 0.208833
R5922 VDPWR.n122 VDPWR.n118 0.208833
R5923 VDPWR.n134 VDPWR.n113 0.208833
R5924 VDPWR.n130 VDPWR.n113 0.208833
R5925 VDPWR.n130 VDPWR.n129 0.208833
R5926 VDPWR.n150 VDPWR.n137 0.208833
R5927 VDPWR.n146 VDPWR.n137 0.208833
R5928 VDPWR.n146 VDPWR.n145 0.208833
R5929 VDPWR.n145 VDPWR.n144 0.208833
R5930 VDPWR.n144 VDPWR.n140 0.208833
R5931 VDPWR.n156 VDPWR.n135 0.208833
R5932 VDPWR.n152 VDPWR.n135 0.208833
R5933 VDPWR.n152 VDPWR.n151 0.208833
R5934 VDPWR.n181 VDPWR.n168 0.208833
R5935 VDPWR.n177 VDPWR.n168 0.208833
R5936 VDPWR.n177 VDPWR.n176 0.208833
R5937 VDPWR.n176 VDPWR.n175 0.208833
R5938 VDPWR.n175 VDPWR.n171 0.208833
R5939 VDPWR.n187 VDPWR.n166 0.208833
R5940 VDPWR.n183 VDPWR.n166 0.208833
R5941 VDPWR.n183 VDPWR.n182 0.208833
R5942 VDPWR.n498 VDPWR.n421 0.20853
R5943 VDPWR.n461 VDPWR.n460 0.188
R5944 VDPWR.n622 VDPWR.n621 0.188
R5945 VDPWR.n621 VDPWR.n620 0.188
R5946 VDPWR.n620 VDPWR.n619 0.188
R5947 VDPWR.n619 VDPWR.n618 0.188
R5948 VDPWR.n618 VDPWR.n617 0.188
R5949 VDPWR.n617 VDPWR.n616 0.188
R5950 VDPWR.n616 VDPWR.n615 0.188
R5951 VDPWR.n615 VDPWR.n614 0.188
R5952 VDPWR.n110 VDPWR.n109 0.188
R5953 VDPWR.n69 VDPWR.n62 0.188
R5954 VDPWR.n669 VDPWR.n668 0.182048
R5955 VDPWR.n679 VDPWR.n678 0.182048
R5956 VDPWR.n663 VDPWR.n662 0.182048
R5957 VDPWR.n673 VDPWR.n672 0.182048
R5958 VDPWR.n683 VDPWR.n682 0.178305
R5959 VDPWR.t173 VDPWR.t399 0.1603
R5960 VDPWR.t137 VDPWR.t173 0.1603
R5961 VDPWR.t384 VDPWR.t137 0.1603
R5962 VDPWR.t112 VDPWR.t384 0.1603
R5963 VDPWR.t377 VDPWR.t112 0.1603
R5964 VDPWR.t368 VDPWR.t377 0.1603
R5965 VDPWR.t56 VDPWR.t368 0.1603
R5966 VDPWR.t196 VDPWR.t56 0.1603
R5967 VDPWR.t142 VDPWR.t123 0.1603
R5968 VDPWR.t57 VDPWR.t142 0.1603
R5969 VDPWR.t388 VDPWR.t57 0.1603
R5970 VDPWR.t46 VDPWR.t388 0.1603
R5971 VDPWR.t422 VDPWR.t46 0.1603
R5972 VDPWR.t385 VDPWR.t422 0.1603
R5973 VDPWR.t47 VDPWR.t385 0.1603
R5974 VDPWR.t423 VDPWR.t47 0.1603
R5975 VDPWR.t376 VDPWR.n417 0.159278
R5976 VDPWR.n486 VDPWR.n424 0.15675
R5977 VDPWR.n468 VDPWR.n437 0.15675
R5978 VDPWR.n461 VDPWR.n437 0.15675
R5979 VDPWR.n109 VDPWR.n51 0.15675
R5980 VDPWR.n70 VDPWR.n69 0.15675
R5981 VDPWR.t123 VDPWR.t376 0.137822
R5982 VDPWR.n417 VDPWR.t196 0.1368
R5983 VDPWR.n454 VDPWR.n428 0.1255
R5984 VDPWR.n456 VDPWR.n455 0.1255
R5985 VDPWR.n557 VDPWR.n500 0.1255
R5986 VDPWR.n504 VDPWR.n500 0.1255
R5987 VDPWR.n506 VDPWR.n504 0.1255
R5988 VDPWR.n508 VDPWR.n506 0.1255
R5989 VDPWR.n510 VDPWR.n508 0.1255
R5990 VDPWR.n512 VDPWR.n510 0.1255
R5991 VDPWR.n514 VDPWR.n512 0.1255
R5992 VDPWR.n516 VDPWR.n514 0.1255
R5993 VDPWR.n518 VDPWR.n516 0.1255
R5994 VDPWR.n548 VDPWR.n518 0.1255
R5995 VDPWR.n547 VDPWR.n520 0.1255
R5996 VDPWR.n524 VDPWR.n520 0.1255
R5997 VDPWR.n526 VDPWR.n524 0.1255
R5998 VDPWR.n528 VDPWR.n526 0.1255
R5999 VDPWR.n530 VDPWR.n528 0.1255
R6000 VDPWR.n532 VDPWR.n530 0.1255
R6001 VDPWR.n534 VDPWR.n532 0.1255
R6002 VDPWR.n536 VDPWR.n534 0.1255
R6003 VDPWR.n538 VDPWR.n536 0.1255
R6004 VDPWR.n350 VDPWR.n233 0.1255
R6005 VDPWR.n349 VDPWR.n348 0.1255
R6006 VDPWR.n558 VDPWR.n498 0.118442
R6007 VDPWR.n681 VDPWR.n635 0.10278
R6008 VDPWR.n87 VDPWR.n58 0.0451429
R6009 VDPWR.n89 VDPWR.n87 0.0451429
R6010 VDPWR.n417 VDPWR.t122 0.00152174
R6011 a_11880_10030.n1 a_11880_10030.t32 312.798
R6012 a_11880_10030.n8 a_11880_10030.t24 312.781
R6013 a_11880_10030.n14 a_11880_10030.t45 312.5
R6014 a_11880_10030.n8 a_11880_10030.t31 310.401
R6015 a_11880_10030.n9 a_11880_10030.t43 310.401
R6016 a_11880_10030.n10 a_11880_10030.t18 310.401
R6017 a_11880_10030.n11 a_11880_10030.t27 310.401
R6018 a_11880_10030.n12 a_11880_10030.t26 310.401
R6019 a_11880_10030.n13 a_11880_10030.t37 310.401
R6020 a_11880_10030.n5 a_11880_10030.t29 310.401
R6021 a_11880_10030.n4 a_11880_10030.t40 310.401
R6022 a_11880_10030.n3 a_11880_10030.t49 310.401
R6023 a_11880_10030.n2 a_11880_10030.t22 310.401
R6024 a_11880_10030.n1 a_11880_10030.t33 310.401
R6025 a_11880_10030.n16 a_11880_10030.t19 308
R6026 a_11880_10030.n28 a_11880_10030.n26 306.808
R6027 a_11880_10030.n0 a_11880_10030.t30 305.901
R6028 a_11880_10030.n20 a_11880_10030.n19 301.933
R6029 a_11880_10030.n22 a_11880_10030.n21 301.933
R6030 a_11880_10030.n24 a_11880_10030.n23 301.933
R6031 a_11880_10030.n29 a_11880_10030.n25 297.433
R6032 a_11880_10030.n28 a_11880_10030.n27 297.433
R6033 a_11880_10030.n18 a_11880_10030.t9 98.9217
R6034 a_11880_10030.n25 a_11880_10030.t10 39.4005
R6035 a_11880_10030.n25 a_11880_10030.t5 39.4005
R6036 a_11880_10030.n26 a_11880_10030.t1 39.4005
R6037 a_11880_10030.n26 a_11880_10030.t13 39.4005
R6038 a_11880_10030.n27 a_11880_10030.t12 39.4005
R6039 a_11880_10030.n27 a_11880_10030.t2 39.4005
R6040 a_11880_10030.n19 a_11880_10030.t7 39.4005
R6041 a_11880_10030.n19 a_11880_10030.t11 39.4005
R6042 a_11880_10030.n21 a_11880_10030.t3 39.4005
R6043 a_11880_10030.n21 a_11880_10030.t4 39.4005
R6044 a_11880_10030.n23 a_11880_10030.t8 39.4005
R6045 a_11880_10030.n23 a_11880_10030.t6 39.4005
R6046 a_11880_10030.n50 a_11880_10030.n30 15.2817
R6047 a_11880_10030.n50 a_11880_10030.n49 13.0946
R6048 a_11880_10030.n20 a_11880_10030.n18 4.90675
R6049 a_11880_10030.n31 a_11880_10030.t21 4.8248
R6050 a_11880_10030.n6 a_11880_10030.n0 4.5005
R6051 a_11880_10030.n17 a_11880_10030.n7 4.5005
R6052 a_11880_10030.n16 a_11880_10030.n15 4.5005
R6053 a_11880_10030.n30 a_11880_10030.n29 4.5005
R6054 a_11880_10030.n39 a_11880_10030.t14 4.5005
R6055 a_11880_10030.n38 a_11880_10030.t39 4.5005
R6056 a_11880_10030.n37 a_11880_10030.t44 4.5005
R6057 a_11880_10030.n36 a_11880_10030.t35 4.5005
R6058 a_11880_10030.n35 a_11880_10030.t25 4.5005
R6059 a_11880_10030.n34 a_11880_10030.t16 4.5005
R6060 a_11880_10030.n33 a_11880_10030.t20 4.5005
R6061 a_11880_10030.n32 a_11880_10030.t47 4.5005
R6062 a_11880_10030.n31 a_11880_10030.t17 4.5005
R6063 a_11880_10030.n40 a_11880_10030.t38 4.5005
R6064 a_11880_10030.n41 a_11880_10030.t28 4.5005
R6065 a_11880_10030.n42 a_11880_10030.t34 4.5005
R6066 a_11880_10030.n43 a_11880_10030.t23 4.5005
R6067 a_11880_10030.n44 a_11880_10030.t15 4.5005
R6068 a_11880_10030.n45 a_11880_10030.t41 4.5005
R6069 a_11880_10030.n46 a_11880_10030.t46 4.5005
R6070 a_11880_10030.n47 a_11880_10030.t36 4.5005
R6071 a_11880_10030.n48 a_11880_10030.t42 4.5005
R6072 a_11880_10030.n49 a_11880_10030.t48 4.5005
R6073 a_11880_10030.t0 a_11880_10030.n50 4.16699
R6074 a_11880_10030.n29 a_11880_10030.n28 1.59425
R6075 a_11880_10030.n18 a_11880_10030.n17 1.21925
R6076 a_11880_10030.n30 a_11880_10030.n24 1.1255
R6077 a_11880_10030.n24 a_11880_10030.n22 1.1255
R6078 a_11880_10030.n22 a_11880_10030.n20 1.1255
R6079 a_11880_10030.n39 a_11880_10030.n38 0.3295
R6080 a_11880_10030.n38 a_11880_10030.n37 0.3295
R6081 a_11880_10030.n37 a_11880_10030.n36 0.3295
R6082 a_11880_10030.n36 a_11880_10030.n35 0.3295
R6083 a_11880_10030.n35 a_11880_10030.n34 0.3295
R6084 a_11880_10030.n34 a_11880_10030.n33 0.3295
R6085 a_11880_10030.n33 a_11880_10030.n32 0.3295
R6086 a_11880_10030.n32 a_11880_10030.n31 0.3295
R6087 a_11880_10030.n41 a_11880_10030.n40 0.3295
R6088 a_11880_10030.n42 a_11880_10030.n41 0.3295
R6089 a_11880_10030.n43 a_11880_10030.n42 0.3295
R6090 a_11880_10030.n44 a_11880_10030.n43 0.3295
R6091 a_11880_10030.n45 a_11880_10030.n44 0.3295
R6092 a_11880_10030.n46 a_11880_10030.n45 0.3295
R6093 a_11880_10030.n47 a_11880_10030.n46 0.3295
R6094 a_11880_10030.n48 a_11880_10030.n47 0.3295
R6095 a_11880_10030.n49 a_11880_10030.n48 0.3248
R6096 a_11880_10030.n40 a_11880_10030.n39 0.2825
R6097 a_11880_10030.n2 a_11880_10030.n1 0.28175
R6098 a_11880_10030.n3 a_11880_10030.n2 0.28175
R6099 a_11880_10030.n4 a_11880_10030.n3 0.28175
R6100 a_11880_10030.n5 a_11880_10030.n4 0.28175
R6101 a_11880_10030.n6 a_11880_10030.n5 0.28175
R6102 a_11880_10030.n15 a_11880_10030.n14 0.28175
R6103 a_11880_10030.n14 a_11880_10030.n13 0.28175
R6104 a_11880_10030.n13 a_11880_10030.n12 0.28175
R6105 a_11880_10030.n12 a_11880_10030.n11 0.28175
R6106 a_11880_10030.n11 a_11880_10030.n10 0.28175
R6107 a_11880_10030.n10 a_11880_10030.n9 0.28175
R6108 a_11880_10030.n9 a_11880_10030.n8 0.28175
R6109 a_11880_10030.n7 a_11880_10030.n6 0.141125
R6110 a_11880_10030.n15 a_11880_10030.n7 0.141125
R6111 a_11880_10030.n17 a_11880_10030.n0 0.141125
R6112 a_11880_10030.n17 a_11880_10030.n16 0.141125
R6113 a_21100_10960.t3 a_21100_10960.n6 818.074
R6114 a_21100_10960.n2 a_21100_10960.n0 297.503
R6115 a_21100_10960.n6 a_21100_10960.t5 289.2
R6116 a_21100_10960.n5 a_21100_10960.t8 289.2
R6117 a_21100_10960.n4 a_21100_10960.t7 289.2
R6118 a_21100_10960.n3 a_21100_10960.t6 232.968
R6119 a_21100_10960.n6 a_21100_10960.n5 208.868
R6120 a_21100_10960.n5 a_21100_10960.n4 208.868
R6121 a_21100_10960.n4 a_21100_10960.n3 199.829
R6122 a_21100_10960.n2 a_21100_10960.n1 195.55
R6123 a_21100_10960.n3 a_21100_10960.n2 172.582
R6124 a_21100_10960.n1 a_21100_10960.t1 60.0005
R6125 a_21100_10960.n1 a_21100_10960.t2 60.0005
R6126 a_21100_10960.n0 a_21100_10960.t4 49.2505
R6127 a_21100_10960.n0 a_21100_10960.t0 49.2505
R6128 a_17450_6090.n14 a_17450_6090.n13 424.447
R6129 a_17450_6090.n3 a_17450_6090.n2 380.8
R6130 a_17450_6090.n14 a_17450_6090.n12 380.8
R6131 a_17450_6090.n15 a_17450_6090.n14 354.046
R6132 a_17450_6090.n2 a_17450_6090.n1 313
R6133 a_17450_6090.n6 a_17450_6090.t13 297.233
R6134 a_17450_6090.n7 a_17450_6090.t13 297.233
R6135 a_17450_6090.t11 a_17450_6090.n4 297.233
R6136 a_17450_6090.n5 a_17450_6090.t11 297.233
R6137 a_17450_6090.n9 a_17450_6090.t0 281.596
R6138 a_17450_6090.n2 a_17450_6090.n0 242.601
R6139 a_17450_6090.n6 a_17450_6090.n5 216.9
R6140 a_17450_6090.n10 a_17450_6090.n8 167.644
R6141 a_17450_6090.n9 a_17450_6090.t9 118.666
R6142 a_17450_6090.n8 a_17450_6090.n7 81.6727
R6143 a_17450_6090.n8 a_17450_6090.n4 81.6727
R6144 a_17450_6090.n7 a_17450_6090.t15 80.3338
R6145 a_17450_6090.t15 a_17450_6090.n6 80.3338
R6146 a_17450_6090.t14 a_17450_6090.n4 80.3338
R6147 a_17450_6090.n5 a_17450_6090.t14 80.3338
R6148 a_17450_6090.n3 a_17450_6090.t12 70.0829
R6149 a_17450_6090.n11 a_17450_6090.n3 64.0005
R6150 a_17450_6090.n12 a_17450_6090.n11 64.0005
R6151 a_17450_6090.n12 a_17450_6090.t10 63.6829
R6152 a_17450_6090.n10 a_17450_6090.n9 60.4288
R6153 a_17450_6090.n1 a_17450_6090.t1 60.0005
R6154 a_17450_6090.n1 a_17450_6090.t8 60.0005
R6155 a_17450_6090.n0 a_17450_6090.t3 60.0005
R6156 a_17450_6090.n0 a_17450_6090.t2 60.0005
R6157 a_17450_6090.n11 a_17450_6090.n10 52.4255
R6158 a_17450_6090.n13 a_17450_6090.t5 49.2505
R6159 a_17450_6090.n13 a_17450_6090.t6 49.2505
R6160 a_17450_6090.t7 a_17450_6090.n15 49.2505
R6161 a_17450_6090.n15 a_17450_6090.t4 49.2505
R6162 ua[1].n14 ua[1].t6 537.245
R6163 ua[1].t4 ua[1].t2 401.668
R6164 ua[1].n14 ua[1].t5 386.62
R6165 ua[1].n17 ua[1].n16 366.776
R6166 ua[1].n16 ua[1].t3 353.467
R6167 ua[1].n16 ua[1].t4 257.067
R6168 ua[1].n33 ua[1].t0 236.579
R6169 ua[1].n33 ua[1].t1 135.501
R6170 ua[1] ua[1].n37 5.00166
R6171 ua[1].n19 ua[1].n18 4.5005
R6172 ua[1].n15 ua[1].n13 4.5005
R6173 ua[1].n28 ua[1].n8 4.5005
R6174 ua[1].n27 ua[1].n26 4.5005
R6175 ua[1].n28 ua[1].n27 4.5005
R6176 ua[1].n5 ua[1].n4 4.5005
R6177 ua[1].n37 ua[1].n0 4.5005
R6178 ua[1].n36 ua[1].n35 4.5005
R6179 ua[1].n37 ua[1].n36 4.5005
R6180 ua[1].n6 ua[1].n3 2.26187
R6181 ua[1].n7 ua[1].n6 2.26187
R6182 ua[1].n34 ua[1].n1 2.26187
R6183 ua[1].n18 ua[1].n17 2.25615
R6184 ua[1].n20 ua[1].n19 2.24063
R6185 ua[1].n26 ua[1].n25 2.24063
R6186 ua[1].n11 ua[1].n10 2.24063
R6187 ua[1].n35 ua[1].n34 2.24063
R6188 ua[1].n32 ua[1].n2 2.24063
R6189 ua[1].n23 ua[1].n12 2.24063
R6190 ua[1].n22 ua[1].n21 2.24063
R6191 ua[1].n24 ua[1].n9 2.24063
R6192 ua[1].n31 ua[1].n3 2.24063
R6193 ua[1].n30 ua[1].n29 2.24063
R6194 ua[1].n35 ua[1].n33 1.84657
R6195 ua[1].n21 ua[1].n14 1.57053
R6196 ua[1].n29 ua[1].n28 1.14633
R6197 ua[1].n24 ua[1].n23 0.740083
R6198 ua[1].n36 ua[1].n31 0.740083
R6199 ua[1].n19 ua[1].n13 0.0421667
R6200 ua[1].n26 ua[1].n11 0.0421667
R6201 ua[1].n35 ua[1].n32 0.0421667
R6202 ua[1].n17 ua[1].n13 0.0226148
R6203 ua[1].n21 ua[1].n20 0.0217373
R6204 ua[1].n25 ua[1].n24 0.0217373
R6205 ua[1].n27 ua[1].n10 0.0217373
R6206 ua[1].n20 ua[1].n15 0.0217373
R6207 ua[1].n29 ua[1].n7 0.0217373
R6208 ua[1].n25 ua[1].n8 0.0217373
R6209 ua[1].n10 ua[1].n8 0.0217373
R6210 ua[1].n36 ua[1].n2 0.0217373
R6211 ua[1].n6 ua[1].n4 0.0217373
R6212 ua[1].n7 ua[1].n5 0.0217373
R6213 ua[1].n34 ua[1].n0 0.0217373
R6214 ua[1].n2 ua[1].n0 0.0217373
R6215 ua[1].n15 ua[1].n12 0.0217373
R6216 ua[1].n22 ua[1].n13 0.0217373
R6217 ua[1].n18 ua[1].n12 0.0217373
R6218 ua[1].n23 ua[1].n22 0.0217373
R6219 ua[1].n5 ua[1].n3 0.0217373
R6220 ua[1].n28 ua[1].n9 0.0217373
R6221 ua[1].n11 ua[1].n9 0.0217373
R6222 ua[1].n30 ua[1].n4 0.0217373
R6223 ua[1].n31 ua[1].n30 0.0217373
R6224 ua[1].n37 ua[1].n1 0.0217373
R6225 ua[1].n32 ua[1].n1 0.0217373
R6226 a_21810_3370.n0 a_21810_3370.t1 752.333
R6227 a_21810_3370.t2 a_21810_3370.n5 752.333
R6228 a_21810_3370.n1 a_21810_3370.t6 514.134
R6229 a_21810_3370.n4 a_21810_3370.n3 366.856
R6230 a_21810_3370.n0 a_21810_3370.t0 254.333
R6231 a_21810_3370.n4 a_21810_3370.t4 190.123
R6232 a_21810_3370.n5 a_21810_3370.n4 187.201
R6233 a_21810_3370.n3 a_21810_3370.n2 176.733
R6234 a_21810_3370.n2 a_21810_3370.n1 176.733
R6235 a_21810_3370.n1 a_21810_3370.t7 112.468
R6236 a_21810_3370.n2 a_21810_3370.t5 112.468
R6237 a_21810_3370.n3 a_21810_3370.t3 112.468
R6238 a_21810_3370.n5 a_21810_3370.n0 70.4005
R6239 a_16900_6090.n0 a_16900_6090.t5 1205
R6240 a_16900_6090.n2 a_16900_6090.t2 522.168
R6241 a_16900_6090.n1 a_16900_6090.n0 441.834
R6242 a_16900_6090.n3 a_16900_6090.n2 235.201
R6243 a_16900_6090.t1 a_16900_6090.n3 229.127
R6244 a_16900_6090.n1 a_16900_6090.t3 217.905
R6245 a_16900_6090.n0 a_16900_6090.t4 208.868
R6246 a_16900_6090.n3 a_16900_6090.t0 158.335
R6247 a_16900_6090.n2 a_16900_6090.n1 15.063
R6248 a_17290_6090.n1 a_17290_6090.n0 409.067
R6249 a_17290_6090.n0 a_17290_6090.t2 403.38
R6250 a_17290_6090.n0 a_17290_6090.t3 369.534
R6251 a_17290_6090.t1 a_17290_6090.n1 209.928
R6252 a_17290_6090.n1 a_17290_6090.t0 177.536
R6253 a_13440_6060.t7 a_13440_6060.t5 835.467
R6254 a_13440_6060.n2 a_13440_6060.t6 517.347
R6255 a_13440_6060.n0 a_13440_6060.t3 465.933
R6256 a_13440_6060.n1 a_13440_6060.n0 458.469
R6257 a_13440_6060.n1 a_13440_6060.t7 398.767
R6258 a_13440_6060.n0 a_13440_6060.t4 321.334
R6259 a_13440_6060.n5 a_13440_6060.n4 244.716
R6260 a_13440_6060.n2 a_13440_6060.t8 228.148
R6261 a_13440_6060.t1 a_13440_6060.n5 221.411
R6262 a_13440_6060.n3 a_13440_6060.n2 216
R6263 a_13440_6060.n5 a_13440_6060.n3 201.573
R6264 a_13440_6060.n3 a_13440_6060.n1 121.451
R6265 a_13440_6060.n4 a_13440_6060.t2 24.0005
R6266 a_13440_6060.n4 a_13440_6060.t0 24.0005
R6267 a_16510_6090.n0 a_16510_6090.t2 441.834
R6268 a_16510_6090.n0 a_16510_6090.t3 313.3
R6269 a_16510_6090.n1 a_16510_6090.n0 235.201
R6270 a_16510_6090.t1 a_16510_6090.n1 219.528
R6271 a_16510_6090.n1 a_16510_6090.t0 167.935
R6272 a_16740_3080.n3 a_16740_3080.n2 742.51
R6273 a_16740_3080.n9 a_16740_3080.t1 723.534
R6274 a_16740_3080.n8 a_16740_3080.t0 723.534
R6275 a_16740_3080.n2 a_16740_3080.n1 684.806
R6276 a_16740_3080.n7 a_16740_3080.n6 366.856
R6277 a_16740_3080.n0 a_16740_3080.t10 337.401
R6278 a_16740_3080.n0 a_16740_3080.t3 305.267
R6279 a_16740_3080.t2 a_16740_3080.n9 254.333
R6280 a_16740_3080.n4 a_16740_3080.n3 224.934
R6281 a_16740_3080.n7 a_16740_3080.t8 190.123
R6282 a_16740_3080.n8 a_16740_3080.n7 187.201
R6283 a_16740_3080.n1 a_16740_3080.n0 176.733
R6284 a_16740_3080.n6 a_16740_3080.n5 176.733
R6285 a_16740_3080.n5 a_16740_3080.n4 176.733
R6286 a_16740_3080.n3 a_16740_3080.t9 144.601
R6287 a_16740_3080.n2 a_16740_3080.t5 131.976
R6288 a_16740_3080.n0 a_16740_3080.t7 128.534
R6289 a_16740_3080.n1 a_16740_3080.t11 128.534
R6290 a_16740_3080.n4 a_16740_3080.t4 112.468
R6291 a_16740_3080.n5 a_16740_3080.t12 112.468
R6292 a_16740_3080.n6 a_16740_3080.t6 112.468
R6293 a_16740_3080.n9 a_16740_3080.n8 70.4005
R6294 a_16630_3080.n0 a_16630_3080.t3 723.534
R6295 a_16630_3080.n1 a_16630_3080.t4 553.534
R6296 a_16630_3080.n0 a_16630_3080.t0 254.333
R6297 a_16630_3080.n2 a_16630_3080.n1 206.333
R6298 a_16630_3080.n1 a_16630_3080.n0 70.4005
R6299 a_16630_3080.n2 a_16630_3080.t1 48.0005
R6300 a_16630_3080.t2 a_16630_3080.n2 48.0005
R6301 a_19440_11540.n3 a_19440_11540.t4 384.967
R6302 a_19440_11540.n0 a_19440_11540.t7 384.967
R6303 a_19440_11540.n3 a_19440_11540.t6 378.36
R6304 a_19440_11540.t8 a_19440_11540.n0 375.897
R6305 a_19440_11540.n4 a_19440_11540.n2 313.846
R6306 a_19440_11540.n5 a_19440_11540.n1 313.846
R6307 a_19440_11540.n11 a_19440_11540.n10 312.998
R6308 a_19440_11540.n8 a_19440_11540.n7 130.143
R6309 a_19440_11540.n8 a_19440_11540.n6 119.267
R6310 a_19440_11540.n5 a_19440_11540.n4 83.2005
R6311 a_19440_11540.n2 a_19440_11540.t9 49.2505
R6312 a_19440_11540.n2 a_19440_11540.t5 49.2505
R6313 a_19440_11540.n1 a_19440_11540.t0 49.2505
R6314 a_19440_11540.n1 a_19440_11540.t12 49.2505
R6315 a_19440_11540.t8 a_19440_11540.n11 49.2505
R6316 a_19440_11540.n11 a_19440_11540.t1 49.2505
R6317 a_19440_11540.n10 a_19440_11540.n9 49.0672
R6318 a_19440_11540.n6 a_19440_11540.t2 19.7005
R6319 a_19440_11540.n6 a_19440_11540.t10 19.7005
R6320 a_19440_11540.n7 a_19440_11540.t3 19.7005
R6321 a_19440_11540.n7 a_19440_11540.t11 19.7005
R6322 a_19440_11540.n9 a_19440_11540.n5 17.0672
R6323 a_19440_11540.n4 a_19440_11540.n3 16.0005
R6324 a_19440_11540.n10 a_19440_11540.n0 16.0005
R6325 a_19440_11540.n9 a_19440_11540.n8 9.69113
R6326 a_18230_3320.n0 a_18230_3320.t1 713.933
R6327 a_18230_3320.n0 a_18230_3320.t2 314.233
R6328 a_18230_3320.t0 a_18230_3320.n0 308.2
R6329 a_17820_3240.n0 a_17820_3240.t0 721.4
R6330 a_17820_3240.n1 a_17820_3240.t4 350.349
R6331 a_17820_3240.n0 a_17820_3240.t2 276.733
R6332 a_17820_3240.n2 a_17820_3240.n1 206.333
R6333 a_17820_3240.n1 a_17820_3240.n0 48.0005
R6334 a_17820_3240.n2 a_17820_3240.t1 48.0005
R6335 a_17820_3240.t3 a_17820_3240.n2 48.0005
R6336 PFET_GATE.n0 PFET_GATE.t17 403.952
R6337 PFET_GATE.n18 PFET_GATE.t29 403.755
R6338 PFET_GATE.n17 PFET_GATE.t18 403.755
R6339 PFET_GATE.n16 PFET_GATE.t16 403.755
R6340 PFET_GATE.n15 PFET_GATE.t24 403.755
R6341 PFET_GATE.n14 PFET_GATE.t13 403.755
R6342 PFET_GATE.n13 PFET_GATE.t22 403.755
R6343 PFET_GATE.n12 PFET_GATE.t11 403.755
R6344 PFET_GATE.n11 PFET_GATE.t20 403.755
R6345 PFET_GATE.n10 PFET_GATE.t25 403.755
R6346 PFET_GATE.n9 PFET_GATE.t14 403.755
R6347 PFET_GATE.n8 PFET_GATE.t10 403.755
R6348 PFET_GATE.n7 PFET_GATE.t19 403.755
R6349 PFET_GATE.n6 PFET_GATE.t28 403.755
R6350 PFET_GATE.n5 PFET_GATE.t26 403.755
R6351 PFET_GATE.n4 PFET_GATE.t15 403.755
R6352 PFET_GATE.n3 PFET_GATE.t23 403.755
R6353 PFET_GATE.n2 PFET_GATE.t12 403.755
R6354 PFET_GATE.n1 PFET_GATE.t21 403.755
R6355 PFET_GATE.n0 PFET_GATE.t27 403.755
R6356 PFET_GATE.n26 PFET_GATE.n25 301.933
R6357 PFET_GATE.n24 PFET_GATE.n23 301.933
R6358 PFET_GATE.n22 PFET_GATE.n21 301.933
R6359 PFET_GATE.n20 PFET_GATE.n19 301.933
R6360 PFET_GATE.n20 PFET_GATE.t7 103.828
R6361 PFET_GATE.n25 PFET_GATE.t4 39.4005
R6362 PFET_GATE.n25 PFET_GATE.t8 39.4005
R6363 PFET_GATE.n23 PFET_GATE.t6 39.4005
R6364 PFET_GATE.n23 PFET_GATE.t2 39.4005
R6365 PFET_GATE.n21 PFET_GATE.t1 39.4005
R6366 PFET_GATE.n21 PFET_GATE.t3 39.4005
R6367 PFET_GATE.n19 PFET_GATE.t9 39.4005
R6368 PFET_GATE.n19 PFET_GATE.t5 39.4005
R6369 PFET_GATE.n27 PFET_GATE.n18 13.3157
R6370 PFET_GATE.t0 PFET_GATE.n27 12.4345
R6371 PFET_GATE.n27 PFET_GATE.n26 7.92238
R6372 PFET_GATE.n9 PFET_GATE.n8 1.6255
R6373 PFET_GATE.n22 PFET_GATE.n20 1.1255
R6374 PFET_GATE.n24 PFET_GATE.n22 1.1255
R6375 PFET_GATE.n26 PFET_GATE.n24 1.1255
R6376 PFET_GATE.n1 PFET_GATE.n0 0.196929
R6377 PFET_GATE.n2 PFET_GATE.n1 0.196929
R6378 PFET_GATE.n3 PFET_GATE.n2 0.196929
R6379 PFET_GATE.n4 PFET_GATE.n3 0.196929
R6380 PFET_GATE.n5 PFET_GATE.n4 0.196929
R6381 PFET_GATE.n6 PFET_GATE.n5 0.196929
R6382 PFET_GATE.n7 PFET_GATE.n6 0.196929
R6383 PFET_GATE.n8 PFET_GATE.n7 0.196929
R6384 PFET_GATE.n10 PFET_GATE.n9 0.196929
R6385 PFET_GATE.n11 PFET_GATE.n10 0.196929
R6386 PFET_GATE.n12 PFET_GATE.n11 0.196929
R6387 PFET_GATE.n13 PFET_GATE.n12 0.196929
R6388 PFET_GATE.n14 PFET_GATE.n13 0.196929
R6389 PFET_GATE.n15 PFET_GATE.n14 0.196929
R6390 PFET_GATE.n16 PFET_GATE.n15 0.196929
R6391 PFET_GATE.n17 PFET_GATE.n16 0.196929
R6392 PFET_GATE.n18 PFET_GATE.n17 0.196929
R6393 a_21210_3400.t3 a_21210_3400.t5 1012.2
R6394 a_21210_3400.n0 a_21210_3400.t0 663.801
R6395 a_21210_3400.n2 a_21210_3400.n1 431.401
R6396 a_21210_3400.t4 a_21210_3400.t6 401.668
R6397 a_21210_3400.n0 a_21210_3400.t3 361.692
R6398 a_21210_3400.n1 a_21210_3400.t2 353.467
R6399 a_21210_3400.t1 a_21210_3400.n2 298.921
R6400 a_21210_3400.n1 a_21210_3400.t4 257.067
R6401 a_21210_3400.n2 a_21210_3400.n0 67.2005
R6402 a_20510_3370.n4 a_20510_3370.t1 752.333
R6403 a_20510_3370.t2 a_20510_3370.n5 752.333
R6404 a_20510_3370.n0 a_20510_3370.t5 514.134
R6405 a_20510_3370.n3 a_20510_3370.n2 366.856
R6406 a_20510_3370.n5 a_20510_3370.t0 254.333
R6407 a_20510_3370.n3 a_20510_3370.t3 190.123
R6408 a_20510_3370.n4 a_20510_3370.n3 187.201
R6409 a_20510_3370.n2 a_20510_3370.n1 176.733
R6410 a_20510_3370.n1 a_20510_3370.n0 176.733
R6411 a_20510_3370.n0 a_20510_3370.t7 112.468
R6412 a_20510_3370.n1 a_20510_3370.t4 112.468
R6413 a_20510_3370.n2 a_20510_3370.t6 112.468
R6414 a_20510_3370.n5 a_20510_3370.n4 70.4005
R6415 a_19670_10930.n1 a_19670_10930.t6 321.334
R6416 a_19670_10930.n4 a_19670_10930.n0 298.503
R6417 a_19670_10930.n2 a_19670_10930.n1 208.868
R6418 a_19670_10930.n5 a_19670_10930.n4 194.488
R6419 a_19670_10930.n3 a_19670_10930.t3 174.056
R6420 a_19670_10930.n4 a_19670_10930.n3 161.3
R6421 a_19670_10930.n2 a_19670_10930.t1 112.468
R6422 a_19670_10930.n1 a_19670_10930.t7 112.468
R6423 a_19670_10930.n3 a_19670_10930.n2 61.5894
R6424 a_19670_10930.n5 a_19670_10930.t2 60.0005
R6425 a_19670_10930.t4 a_19670_10930.n5 60.0005
R6426 a_19670_10930.n0 a_19670_10930.t5 49.2505
R6427 a_19670_10930.n0 a_19670_10930.t0 49.2505
R6428 ua[0].n0 ua[0].t0 514.134
R6429 ua[0] ua[0].n0 461.62
R6430 ua[0].n0 ua[0].t1 273.134
R6431 a_13360_6510.t0 a_13360_6510.t1 39.4005
R6432 a_13880_11590.n15 a_13880_11590.t21 310.488
R6433 a_13880_11590.n9 a_13880_11590.t20 310.488
R6434 a_13880_11590.n4 a_13880_11590.t19 310.488
R6435 a_13880_11590.n13 a_13880_11590.n12 297.433
R6436 a_13880_11590.n8 a_13880_11590.n7 297.433
R6437 a_13880_11590.n19 a_13880_11590.n18 297.433
R6438 a_13880_11590.n2 a_13880_11590.t0 248.133
R6439 a_13880_11590.n2 a_13880_11590.n1 199.383
R6440 a_13880_11590.n3 a_13880_11590.n0 194.883
R6441 a_13880_11590.n17 a_13880_11590.t14 184.097
R6442 a_13880_11590.n11 a_13880_11590.t12 184.097
R6443 a_13880_11590.n6 a_13880_11590.t4 184.097
R6444 a_13880_11590.n16 a_13880_11590.n15 167.094
R6445 a_13880_11590.n10 a_13880_11590.n9 167.094
R6446 a_13880_11590.n5 a_13880_11590.n4 167.094
R6447 a_13880_11590.n18 a_13880_11590.n17 161.3
R6448 a_13880_11590.n13 a_13880_11590.n11 161.3
R6449 a_13880_11590.n8 a_13880_11590.n6 161.3
R6450 a_13880_11590.n15 a_13880_11590.t17 120.501
R6451 a_13880_11590.n16 a_13880_11590.t8 120.501
R6452 a_13880_11590.n9 a_13880_11590.t18 120.501
R6453 a_13880_11590.n10 a_13880_11590.t6 120.501
R6454 a_13880_11590.n4 a_13880_11590.t22 120.501
R6455 a_13880_11590.n5 a_13880_11590.t10 120.501
R6456 a_13880_11590.n1 a_13880_11590.t3 48.0005
R6457 a_13880_11590.n1 a_13880_11590.t2 48.0005
R6458 a_13880_11590.n0 a_13880_11590.t16 48.0005
R6459 a_13880_11590.n0 a_13880_11590.t1 48.0005
R6460 a_13880_11590.n17 a_13880_11590.n16 40.7027
R6461 a_13880_11590.n11 a_13880_11590.n10 40.7027
R6462 a_13880_11590.n6 a_13880_11590.n5 40.7027
R6463 a_13880_11590.n12 a_13880_11590.t13 39.4005
R6464 a_13880_11590.n12 a_13880_11590.t7 39.4005
R6465 a_13880_11590.n7 a_13880_11590.t5 39.4005
R6466 a_13880_11590.n7 a_13880_11590.t11 39.4005
R6467 a_13880_11590.t15 a_13880_11590.n19 39.4005
R6468 a_13880_11590.n19 a_13880_11590.t9 39.4005
R6469 a_13880_11590.n14 a_13880_11590.n13 6.6255
R6470 a_13880_11590.n14 a_13880_11590.n8 6.6255
R6471 a_13880_11590.n3 a_13880_11590.n2 5.2505
R6472 a_13880_11590.n18 a_13880_11590.n14 4.5005
R6473 a_13880_11590.n18 a_13880_11590.n3 0.78175
R6474 a_23830_2840.n0 a_23830_2840.t2 537.245
R6475 a_23830_2840.n0 a_23830_2840.t3 386.62
R6476 a_23830_2840.t1 a_23830_2840.n1 236.581
R6477 a_23830_2840.n1 a_23830_2840.t0 135.5
R6478 a_23830_2840.n1 a_23830_2840.n0 3.08327
R6479 a_24238_3560.n0 a_24238_3560.t0 236.867
R6480 a_24238_3560.n0 a_24238_3560.t2 237.337
R6481 a_24238_3560.t1 a_24238_3560.n0 209.882
R6482 a_9573_16817.n6 a_9573_16817.t9 287.762
R6483 a_9573_16817.n5 a_9573_16817.t7 287.762
R6484 a_9573_16817.n5 a_9573_16817.t10 287.589
R6485 a_9573_16817.n8 a_9573_16817.t11 287.012
R6486 a_9573_16817.n7 a_9573_16817.t8 287.012
R6487 a_9573_16817.n2 a_9573_16817.n0 107.266
R6488 a_9573_16817.n4 a_9573_16817.n3 105.016
R6489 a_9573_16817.n2 a_9573_16817.n1 105.016
R6490 a_9573_16817.n3 a_9573_16817.t3 13.1338
R6491 a_9573_16817.n3 a_9573_16817.t6 13.1338
R6492 a_9573_16817.n1 a_9573_16817.t4 13.1338
R6493 a_9573_16817.n1 a_9573_16817.t1 13.1338
R6494 a_9573_16817.n0 a_9573_16817.t5 13.1338
R6495 a_9573_16817.n0 a_9573_16817.t2 13.1338
R6496 a_9573_16817.t0 a_9573_16817.n9 10.8051
R6497 a_9573_16817.n9 a_9573_16817.n4 10.0474
R6498 a_9573_16817.n9 a_9573_16817.n8 7.97729
R6499 a_9573_16817.n4 a_9573_16817.n2 2.2505
R6500 a_9573_16817.n7 a_9573_16817.n6 0.579071
R6501 a_9573_16817.n8 a_9573_16817.n7 0.282643
R6502 a_9573_16817.n6 a_9573_16817.n5 0.2755
R6503 a_10840_11590.n15 a_10840_11590.t18 310.488
R6504 a_10840_11590.n9 a_10840_11590.t17 310.488
R6505 a_10840_11590.n0 a_10840_11590.t22 310.488
R6506 a_10840_11590.n13 a_10840_11590.n12 297.433
R6507 a_10840_11590.n4 a_10840_11590.n3 297.433
R6508 a_10840_11590.n19 a_10840_11590.n18 297.433
R6509 a_10840_11590.n7 a_10840_11590.t4 248.133
R6510 a_10840_11590.n7 a_10840_11590.n6 199.383
R6511 a_10840_11590.n8 a_10840_11590.n5 194.883
R6512 a_10840_11590.n17 a_10840_11590.t9 184.097
R6513 a_10840_11590.n11 a_10840_11590.t11 184.097
R6514 a_10840_11590.n2 a_10840_11590.t13 184.097
R6515 a_10840_11590.n16 a_10840_11590.n15 167.094
R6516 a_10840_11590.n10 a_10840_11590.n9 167.094
R6517 a_10840_11590.n1 a_10840_11590.n0 167.094
R6518 a_10840_11590.n18 a_10840_11590.n17 161.3
R6519 a_10840_11590.n13 a_10840_11590.n11 161.3
R6520 a_10840_11590.n4 a_10840_11590.n2 161.3
R6521 a_10840_11590.n15 a_10840_11590.t20 120.501
R6522 a_10840_11590.n16 a_10840_11590.t15 120.501
R6523 a_10840_11590.n9 a_10840_11590.t21 120.501
R6524 a_10840_11590.n10 a_10840_11590.t7 120.501
R6525 a_10840_11590.n0 a_10840_11590.t19 120.501
R6526 a_10840_11590.n1 a_10840_11590.t5 120.501
R6527 a_10840_11590.n6 a_10840_11590.t1 48.0005
R6528 a_10840_11590.n6 a_10840_11590.t0 48.0005
R6529 a_10840_11590.n5 a_10840_11590.t2 48.0005
R6530 a_10840_11590.n5 a_10840_11590.t3 48.0005
R6531 a_10840_11590.n17 a_10840_11590.n16 40.7027
R6532 a_10840_11590.n11 a_10840_11590.n10 40.7027
R6533 a_10840_11590.n2 a_10840_11590.n1 40.7027
R6534 a_10840_11590.n12 a_10840_11590.t8 39.4005
R6535 a_10840_11590.n12 a_10840_11590.t12 39.4005
R6536 a_10840_11590.n3 a_10840_11590.t6 39.4005
R6537 a_10840_11590.n3 a_10840_11590.t14 39.4005
R6538 a_10840_11590.t16 a_10840_11590.n19 39.4005
R6539 a_10840_11590.n19 a_10840_11590.t10 39.4005
R6540 a_10840_11590.n14 a_10840_11590.n4 6.6255
R6541 a_10840_11590.n18 a_10840_11590.n14 6.6255
R6542 a_10840_11590.n8 a_10840_11590.n7 5.2505
R6543 a_10840_11590.n14 a_10840_11590.n13 4.5005
R6544 a_10840_11590.n13 a_10840_11590.n8 0.78175
R6545 a_10740_13170.n1 a_10740_13170.n2 199.935
R6546 a_10740_13170.n0 a_10740_13170.n3 199.53
R6547 a_10740_13170.n0 a_10740_13170.n4 199.53
R6548 a_10740_13170.n1 a_10740_13170.n5 199.53
R6549 a_10740_13170.n6 a_10740_13170.n1 199.53
R6550 a_10740_13170.n0 a_10740_13170.t9 97.5404
R6551 a_10740_13170.n3 a_10740_13170.t0 48.0005
R6552 a_10740_13170.n3 a_10740_13170.t5 48.0005
R6553 a_10740_13170.n4 a_10740_13170.t6 48.0005
R6554 a_10740_13170.n4 a_10740_13170.t3 48.0005
R6555 a_10740_13170.n5 a_10740_13170.t2 48.0005
R6556 a_10740_13170.n5 a_10740_13170.t8 48.0005
R6557 a_10740_13170.n2 a_10740_13170.t1 48.0005
R6558 a_10740_13170.n2 a_10740_13170.t10 48.0005
R6559 a_10740_13170.n6 a_10740_13170.t7 48.0005
R6560 a_10740_13170.t4 a_10740_13170.n6 48.0005
R6561 a_10740_13170.n1 a_10740_13170.n0 1.09425
R6562 a_17574_18026.t0 a_17574_18026.t6 57.1093
R6563 a_17574_18026.t4 a_17574_18026.t1 0.1603
R6564 a_17574_18026.t9 a_17574_18026.t4 0.1603
R6565 a_17574_18026.t2 a_17574_18026.t9 0.1603
R6566 a_17574_18026.t5 a_17574_18026.t2 0.1603
R6567 a_17574_18026.t20 a_17574_18026.t5 0.1603
R6568 a_17574_18026.t17 a_17574_18026.t20 0.1603
R6569 a_17574_18026.t10 a_17574_18026.t17 0.1603
R6570 a_17574_18026.t14 a_17574_18026.t10 0.1603
R6571 a_17574_18026.t16 a_17574_18026.t18 0.1603
R6572 a_17574_18026.t19 a_17574_18026.t16 0.1603
R6573 a_17574_18026.t3 a_17574_18026.t19 0.1603
R6574 a_17574_18026.t12 a_17574_18026.t3 0.1603
R6575 a_17574_18026.t8 a_17574_18026.t12 0.1603
R6576 a_17574_18026.t15 a_17574_18026.t8 0.1603
R6577 a_17574_18026.t11 a_17574_18026.t15 0.1603
R6578 a_17574_18026.t6 a_17574_18026.t11 0.1603
R6579 a_17574_18026.t13 a_17574_18026.n0 0.159278
R6580 a_17574_18026.t18 a_17574_18026.t13 0.137822
R6581 a_17574_18026.n0 a_17574_18026.t14 0.1368
R6582 a_17574_18026.n0 a_17574_18026.t7 0.00152174
R6583 a_11431_12690.n2 a_11431_12690.n0 302.507
R6584 a_11431_12690.n10 a_11431_12690.n9 302.163
R6585 a_11431_12690.n8 a_11431_12690.n7 302.163
R6586 a_11431_12690.n6 a_11431_12690.n5 302.163
R6587 a_11431_12690.n4 a_11431_12690.n3 302.163
R6588 a_11431_12690.n2 a_11431_12690.n1 302.163
R6589 a_11431_12690.n11 a_11431_12690.t13 291.502
R6590 a_11431_12690.n14 a_11431_12690.t14 291.288
R6591 a_11431_12690.n13 a_11431_12690.t17 291.288
R6592 a_11431_12690.n12 a_11431_12690.t15 291.288
R6593 a_11431_12690.n11 a_11431_12690.t16 291.288
R6594 a_11431_12690.n9 a_11431_12690.t0 39.4005
R6595 a_11431_12690.n9 a_11431_12690.t11 39.4005
R6596 a_11431_12690.n7 a_11431_12690.t6 39.4005
R6597 a_11431_12690.n7 a_11431_12690.t5 39.4005
R6598 a_11431_12690.n5 a_11431_12690.t8 39.4005
R6599 a_11431_12690.n5 a_11431_12690.t2 39.4005
R6600 a_11431_12690.n3 a_11431_12690.t9 39.4005
R6601 a_11431_12690.n3 a_11431_12690.t3 39.4005
R6602 a_11431_12690.n1 a_11431_12690.t1 39.4005
R6603 a_11431_12690.n1 a_11431_12690.t4 39.4005
R6604 a_11431_12690.n0 a_11431_12690.t10 39.4005
R6605 a_11431_12690.n0 a_11431_12690.t7 39.4005
R6606 a_11431_12690.t12 a_11431_12690.n15 30.8342
R6607 a_11431_12690.n15 a_11431_12690.n10 13.0943
R6608 a_11431_12690.n15 a_11431_12690.n14 7.59693
R6609 a_11431_12690.n12 a_11431_12690.n11 0.643357
R6610 a_11431_12690.n14 a_11431_12690.n13 0.643357
R6611 a_11431_12690.n4 a_11431_12690.n2 0.34425
R6612 a_11431_12690.n6 a_11431_12690.n4 0.34425
R6613 a_11431_12690.n8 a_11431_12690.n6 0.34425
R6614 a_11431_12690.n10 a_11431_12690.n8 0.34425
R6615 a_11431_12690.n13 a_11431_12690.n12 0.214786
R6616 a_16900_7270.n0 a_16900_7270.t4 1028.27
R6617 a_16900_7270.n2 a_16900_7270.n1 569.734
R6618 a_16900_7270.n1 a_16900_7270.n0 465.933
R6619 a_16900_7270.n1 a_16900_7270.t5 401.668
R6620 a_16900_7270.n1 a_16900_7270.t2 385.601
R6621 a_16900_7270.n0 a_16900_7270.t3 385.601
R6622 a_16900_7270.t0 a_16900_7270.n2 211.847
R6623 a_16900_7270.n2 a_16900_7270.t1 173.055
R6624 a_17290_7270.n0 a_17290_7270.t3 605.311
R6625 a_17290_7270.t3 a_17290_7270.t0 420.202
R6626 a_17290_7270.t2 a_17290_7270.n0 240.327
R6627 a_17290_7270.n0 a_17290_7270.t1 148.734
R6628 a_16270_3380.n0 a_16270_3380.t0 663.801
R6629 a_16270_3380.t6 a_16270_3380.t4 514.134
R6630 a_16270_3380.n0 a_16270_3380.t6 479.284
R6631 a_16270_3380.n3 a_16270_3380.n2 344.8
R6632 a_16270_3380.n1 a_16270_3380.t3 289.2
R6633 a_16270_3380.t1 a_16270_3380.n3 275.454
R6634 a_16270_3380.n2 a_16270_3380.t5 241
R6635 a_16270_3380.n1 a_16270_3380.t2 112.468
R6636 a_16270_3380.n3 a_16270_3380.n0 97.9205
R6637 a_16270_3380.n2 a_16270_3380.n1 64.2672
R6638 a_13650_3080.n3 a_13650_3080.n2 919.244
R6639 a_13650_3080.n8 a_13650_3080.n7 918.702
R6640 a_13650_3080.t13 a_13650_3080.t9 819.4
R6641 a_13650_3080.n10 a_13650_3080.n9 628.734
R6642 a_13650_3080.n2 a_13650_3080.n1 520.361
R6643 a_13650_3080.n7 a_13650_3080.n6 364.178
R6644 a_13650_3080.n0 a_13650_3080.t12 337.401
R6645 a_13650_3080.n8 a_13650_3080.t13 336.25
R6646 a_13650_3080.n0 a_13650_3080.t7 305.267
R6647 a_13650_3080.n9 a_13650_3080.t0 257.534
R6648 a_13650_3080.n4 a_13650_3080.t5 192.8
R6649 a_13650_3080.n1 a_13650_3080.n0 176.733
R6650 a_13650_3080.n6 a_13650_3080.n5 176.733
R6651 a_13650_3080.n4 a_13650_3080.n3 160.667
R6652 a_13650_3080.n3 a_13650_3080.t3 144.601
R6653 a_13650_3080.n2 a_13650_3080.t14 131.976
R6654 a_13650_3080.n0 a_13650_3080.t10 128.534
R6655 a_13650_3080.n1 a_13650_3080.t4 128.534
R6656 a_13650_3080.n5 a_13650_3080.t11 112.468
R6657 a_13650_3080.n6 a_13650_3080.t6 112.468
R6658 a_13650_3080.n7 a_13650_3080.t8 112.468
R6659 a_13650_3080.n5 a_13650_3080.n4 96.4005
R6660 a_13650_3080.t2 a_13650_3080.n10 78.8005
R6661 a_13650_3080.n10 a_13650_3080.t1 78.8005
R6662 a_13650_3080.n9 a_13650_3080.n8 11.2005
R6663 a_13440_7240.t8 a_13440_7240.t4 835.467
R6664 a_13440_7240.n2 a_13440_7240.t8 560.011
R6665 a_13440_7240.n0 a_13440_7240.t6 517.347
R6666 a_13440_7240.n1 a_13440_7240.t3 514.134
R6667 a_13440_7240.n2 a_13440_7240.n1 491.791
R6668 a_13440_7240.n3 a_13440_7240.n0 363.2
R6669 a_13440_7240.n1 a_13440_7240.t7 273.134
R6670 a_13440_7240.n5 a_13440_7240.n4 244.716
R6671 a_13440_7240.n0 a_13440_7240.t5 228.148
R6672 a_13440_7240.t1 a_13440_7240.n5 221.411
R6673 a_13440_7240.n5 a_13440_7240.n3 54.3734
R6674 a_13440_7240.n3 a_13440_7240.n2 37.6567
R6675 a_13440_7240.n4 a_13440_7240.t2 24.0005
R6676 a_13440_7240.n4 a_13440_7240.t0 24.0005
R6677 a_16510_7270.t1 a_16510_7270.n1 203.528
R6678 a_16510_7270.n0 a_16510_7270.t2 203.528
R6679 a_16510_7270.n1 a_16510_7270.t0 183.935
R6680 a_16510_7270.n0 a_16510_7270.t3 183.935
R6681 a_16510_7270.n1 a_16510_7270.n0 83.2005
R6682 a_14280_3560.n0 a_14280_3560.t0 723
R6683 a_14280_3560.t3 a_14280_3560.t2 514.134
R6684 a_14280_3560.n0 a_14280_3560.t3 335.983
R6685 a_14280_3560.t1 a_14280_3560.n0 314.921
R6686 a_14120_3110.t0 a_14120_3110.n0 531.067
R6687 a_14120_3110.n0 a_14120_3110.t1 48.0005
R6688 a_14120_3110.n0 a_14120_3110.t2 48.0005
R6689 a_17580_6090.n4 a_17580_6090.t6 297.233
R6690 a_17580_6090.t3 a_17580_6090.n5 297.233
R6691 a_17580_6090.n3 a_17580_6090.n1 257.067
R6692 a_17580_6090.n0 a_17580_6090.t2 241.928
R6693 a_17580_6090.n7 a_17580_6090.n6 237.728
R6694 a_17580_6090.t1 a_17580_6090.n7 235.528
R6695 a_17580_6090.n6 a_17580_6090.n1 226.942
R6696 a_17580_6090.n3 a_17580_6090.n2 226.942
R6697 a_17580_6090.n2 a_17580_6090.t4 220.505
R6698 a_17580_6090.n5 a_17580_6090.n4 216.9
R6699 a_17580_6090.n0 a_17580_6090.t0 145.536
R6700 a_17580_6090.n7 a_17580_6090.n0 121.6
R6701 a_17580_6090.n2 a_17580_6090.t6 92.3838
R6702 a_17580_6090.n6 a_17580_6090.t3 92.3838
R6703 a_17580_6090.t5 a_17580_6090.n3 80.3338
R6704 a_17580_6090.n4 a_17580_6090.t5 80.3338
R6705 a_17580_6090.t7 a_17580_6090.n1 80.3338
R6706 a_17580_6090.n5 a_17580_6090.t7 80.3338
R6707 V_CONT.n25 V_CONT.t13 404.683
R6708 V_CONT.n25 V_CONT.t11 403.755
R6709 V_CONT.n26 V_CONT.t9 403.755
R6710 V_CONT.n27 V_CONT.t14 396.866
R6711 V_CONT.n12 V_CONT.t8 377.567
R6712 V_CONT.n11 V_CONT.t15 297.233
R6713 V_CONT.n13 V_CONT.n11 232.001
R6714 V_CONT.n13 V_CONT.n12 228.2
R6715 V_CONT.n12 V_CONT.t10 216.9
R6716 V_CONT.n22 V_CONT.n21 158.589
R6717 V_CONT.n22 V_CONT.n20 148.901
R6718 V_CONT.n11 V_CONT.t12 136.567
R6719 V_CONT.n7 V_CONT.t4 57.056
R6720 V_CONT.n23 V_CONT.n19 49.3391
R6721 V_CONT.n20 V_CONT.t1 24.6255
R6722 V_CONT.n20 V_CONT.t2 24.6255
R6723 V_CONT.n21 V_CONT.t0 24.6255
R6724 V_CONT.n21 V_CONT.t3 24.6255
R6725 V_CONT.n14 V_CONT.n13 15.4814
R6726 V_CONT.n19 V_CONT.t5 15.0005
R6727 V_CONT.n19 V_CONT.t6 15.0005
R6728 V_CONT.n24 V_CONT.n23 11.7735
R6729 V_CONT.n17 V_CONT.n16 4.5005
R6730 V_CONT.n9 V_CONT.n5 4.5005
R6731 V_CONT.n17 V_CONT.n5 4.5005
R6732 V_CONT.n18 V_CONT.n1 4.5005
R6733 V_CONT.n18 V_CONT.n3 4.5005
R6734 V_CONT.n18 V_CONT.n17 4.5005
R6735 V_CONT.n16 V_CONT.n7 3.85552
R6736 V_CONT.n7 V_CONT.t7 3.7836
R6737 V_CONT V_CONT.n27 3.02137
R6738 V_CONT.n15 V_CONT.n14 2.2458
R6739 V_CONT.n6 V_CONT.n0 2.2458
R6740 V_CONT.n18 V_CONT.n2 2.24063
R6741 V_CONT.n16 V_CONT.n10 2.24063
R6742 V_CONT.n16 V_CONT.n8 2.24063
R6743 V_CONT.n5 V_CONT.n4 2.24063
R6744 V_CONT V_CONT.n24 1.27654
R6745 V_CONT.n27 V_CONT.n26 1.01121
R6746 V_CONT.n26 V_CONT.n25 0.929071
R6747 V_CONT.n23 V_CONT.n22 0.438
R6748 V_CONT.n24 V_CONT.n18 0.336438
R6749 V_CONT.n17 V_CONT.n6 0.0421667
R6750 V_CONT.n14 V_CONT.n2 0.0217373
R6751 V_CONT.n9 V_CONT.n2 0.0217373
R6752 V_CONT.n8 V_CONT.n6 0.0217373
R6753 V_CONT.n4 V_CONT.n1 0.0217373
R6754 V_CONT.n10 V_CONT.n1 0.0217373
R6755 V_CONT.n10 V_CONT.n9 0.0217373
R6756 V_CONT.n8 V_CONT.n3 0.0217373
R6757 V_CONT.n4 V_CONT.n3 0.0217373
R6758 V_CONT.n15 V_CONT.n5 0.0113926
R6759 V_CONT.n16 V_CONT.n15 0.0113926
R6760 V_CONT.n18 V_CONT.n0 0.0113926
R6761 V_CONT.n5 V_CONT.n0 0.0113926
R6762 a_23718_3560.n0 a_23718_3560.t1 236.867
R6763 a_23718_3560.n0 a_23718_3560.t0 237.337
R6764 a_23718_3560.t2 a_23718_3560.n0 209.882
R6765 a_12360_3440.n3 a_12360_3440.t6 772.196
R6766 a_12360_3440.n1 a_12360_3440.t0 756.067
R6767 a_12360_3440.n4 a_12360_3440.n3 607.465
R6768 a_12360_3440.n0 a_12360_3440.t2 514.134
R6769 a_12360_3440.t6 a_12360_3440.t3 514.134
R6770 a_12360_3440.n1 a_12360_3440.n0 438.507
R6771 a_12360_3440.n2 a_12360_3440.t4 289.2
R6772 a_12360_3440.n0 a_12360_3440.t5 273.134
R6773 a_12360_3440.t1 a_12360_3440.n4 233
R6774 a_12360_3440.n3 a_12360_3440.n2 208.868
R6775 a_12360_3440.n2 a_12360_3440.t7 176.733
R6776 a_12360_3440.n4 a_12360_3440.n1 31.7872
R6777 a_13360_7270.t0 a_13360_7270.t1 39.4005
R6778 a_11580_15080.t0 a_11580_15080.n129 172.969
R6779 a_11580_15080.n119 a_11580_15080.n118 83.5719
R6780 a_11580_15080.n121 a_11580_15080.n120 83.5719
R6781 a_11580_15080.n123 a_11580_15080.n122 83.5719
R6782 a_11580_15080.n109 a_11580_15080.n108 83.5719
R6783 a_11580_15080.n101 a_11580_15080.n11 83.5719
R6784 a_11580_15080.n94 a_11580_15080.n12 83.5719
R6785 a_11580_15080.n96 a_11580_15080.n95 83.5719
R6786 a_11580_15080.n88 a_11580_15080.n16 83.5719
R6787 a_11580_15080.n83 a_11580_15080.n17 83.5719
R6788 a_11580_15080.n75 a_11580_15080.n74 83.5719
R6789 a_11580_15080.n73 a_11580_15080.n72 83.5719
R6790 a_11580_15080.n71 a_11580_15080.n70 83.5719
R6791 a_11580_15080.n41 a_11580_15080.n40 83.5719
R6792 a_11580_15080.n48 a_11580_15080.n47 83.5719
R6793 a_11580_15080.n34 a_11580_15080.n31 83.5719
R6794 a_11580_15080.n53 a_11580_15080.n30 83.5719
R6795 a_11580_15080.n60 a_11580_15080.n59 83.5719
R6796 a_11580_15080.n28 a_11580_15080.n26 83.5719
R6797 a_11580_15080.n119 a_11580_15080.n117 73.3165
R6798 a_11580_15080.n103 a_11580_15080.n11 73.3165
R6799 a_11580_15080.n90 a_11580_15080.n16 73.3165
R6800 a_11580_15080.n76 a_11580_15080.n75 73.3165
R6801 a_11580_15080.n47 a_11580_15080.n46 73.3165
R6802 a_11580_15080.n59 a_11580_15080.n58 73.3165
R6803 a_11580_15080.n122 a_11580_15080.n6 73.19
R6804 a_11580_15080.n108 a_11580_15080.n107 73.19
R6805 a_11580_15080.n95 a_11580_15080.n93 73.19
R6806 a_11580_15080.n71 a_11580_15080.n23 73.19
R6807 a_11580_15080.n40 a_11580_15080.n35 73.19
R6808 a_11580_15080.n55 a_11580_15080.n30 73.19
R6809 a_11580_15080.n84 a_11580_15080.t4 65.0299
R6810 a_11580_15080.t3 a_11580_15080.n24 65.0299
R6811 a_11580_15080.n111 a_11580_15080.t1 36.6639
R6812 a_11580_15080.t8 a_11580_15080.n39 36.6639
R6813 a_11580_15080.n121 a_11580_15080.n119 26.074
R6814 a_11580_15080.n94 a_11580_15080.n11 26.074
R6815 a_11580_15080.n83 a_11580_15080.n16 26.074
R6816 a_11580_15080.n75 a_11580_15080.n73 26.074
R6817 a_11580_15080.n47 a_11580_15080.n34 26.074
R6818 a_11580_15080.n59 a_11580_15080.n28 26.074
R6819 a_11580_15080.n122 a_11580_15080.t6 25.7843
R6820 a_11580_15080.n108 a_11580_15080.t1 25.7843
R6821 a_11580_15080.n95 a_11580_15080.t7 25.7843
R6822 a_11580_15080.t2 a_11580_15080.n71 25.7843
R6823 a_11580_15080.n40 a_11580_15080.t8 25.7843
R6824 a_11580_15080.t5 a_11580_15080.n30 25.7843
R6825 a_11580_15080.n77 a_11580_15080.n65 9.3005
R6826 a_11580_15080.n65 a_11580_15080.n21 9.3005
R6827 a_11580_15080.n65 a_11580_15080.n22 9.3005
R6828 a_11580_15080.n81 a_11580_15080.n65 9.3005
R6829 a_11580_15080.n67 a_11580_15080.n21 9.3005
R6830 a_11580_15080.n67 a_11580_15080.n22 9.3005
R6831 a_11580_15080.n67 a_11580_15080.n19 9.3005
R6832 a_11580_15080.n81 a_11580_15080.n67 9.3005
R6833 a_11580_15080.n82 a_11580_15080.n21 9.3005
R6834 a_11580_15080.n82 a_11580_15080.n20 9.3005
R6835 a_11580_15080.n82 a_11580_15080.n22 9.3005
R6836 a_11580_15080.n82 a_11580_15080.n19 9.3005
R6837 a_11580_15080.n82 a_11580_15080.n81 9.3005
R6838 a_11580_15080.n81 a_11580_15080.n69 9.3005
R6839 a_11580_15080.n69 a_11580_15080.n19 9.3005
R6840 a_11580_15080.n69 a_11580_15080.n22 9.3005
R6841 a_11580_15080.n69 a_11580_15080.n20 9.3005
R6842 a_11580_15080.n81 a_11580_15080.n64 9.3005
R6843 a_11580_15080.n64 a_11580_15080.n19 9.3005
R6844 a_11580_15080.n64 a_11580_15080.n22 9.3005
R6845 a_11580_15080.n64 a_11580_15080.n20 9.3005
R6846 a_11580_15080.n77 a_11580_15080.n64 9.3005
R6847 a_11580_15080.n80 a_11580_15080.n21 9.3005
R6848 a_11580_15080.n80 a_11580_15080.n20 9.3005
R6849 a_11580_15080.n80 a_11580_15080.n22 9.3005
R6850 a_11580_15080.n81 a_11580_15080.n80 9.3005
R6851 a_11580_15080.n128 a_11580_15080.n3 9.3005
R6852 a_11580_15080.n128 a_11580_15080.n4 9.3005
R6853 a_11580_15080.n128 a_11580_15080.n2 9.3005
R6854 a_11580_15080.n128 a_11580_15080.n5 9.3005
R6855 a_11580_15080.n128 a_11580_15080.n127 9.3005
R6856 a_11580_15080.n115 a_11580_15080.n4 9.3005
R6857 a_11580_15080.n115 a_11580_15080.n2 9.3005
R6858 a_11580_15080.n115 a_11580_15080.n5 9.3005
R6859 a_11580_15080.n127 a_11580_15080.n115 9.3005
R6860 a_11580_15080.n113 a_11580_15080.n4 9.3005
R6861 a_11580_15080.n113 a_11580_15080.n2 9.3005
R6862 a_11580_15080.n113 a_11580_15080.n5 9.3005
R6863 a_11580_15080.n124 a_11580_15080.n113 9.3005
R6864 a_11580_15080.n127 a_11580_15080.n113 9.3005
R6865 a_11580_15080.n127 a_11580_15080.n126 9.3005
R6866 a_11580_15080.n126 a_11580_15080.n124 9.3005
R6867 a_11580_15080.n126 a_11580_15080.n5 9.3005
R6868 a_11580_15080.n126 a_11580_15080.n2 9.3005
R6869 a_11580_15080.n127 a_11580_15080.n7 9.3005
R6870 a_11580_15080.n124 a_11580_15080.n7 9.3005
R6871 a_11580_15080.n7 a_11580_15080.n5 9.3005
R6872 a_11580_15080.n7 a_11580_15080.n2 9.3005
R6873 a_11580_15080.n7 a_11580_15080.n3 9.3005
R6874 a_11580_15080.n4 a_11580_15080.n0 9.3005
R6875 a_11580_15080.n2 a_11580_15080.n0 9.3005
R6876 a_11580_15080.n5 a_11580_15080.n0 9.3005
R6877 a_11580_15080.n124 a_11580_15080.n0 9.3005
R6878 a_11580_15080.n127 a_11580_15080.n0 9.3005
R6879 a_11580_15080.n79 a_11580_15080.n19 4.64654
R6880 a_11580_15080.n66 a_11580_15080.n20 4.64654
R6881 a_11580_15080.n77 a_11580_15080.n18 4.64654
R6882 a_11580_15080.n68 a_11580_15080.n21 4.64654
R6883 a_11580_15080.n78 a_11580_15080.n77 4.64654
R6884 a_11580_15080.n124 a_11580_15080.n1 4.64654
R6885 a_11580_15080.n114 a_11580_15080.n3 4.64654
R6886 a_11580_15080.n116 a_11580_15080.n4 4.64654
R6887 a_11580_15080.n125 a_11580_15080.n3 4.64654
R6888 a_11580_15080.n107 a_11580_15080.n106 2.36206
R6889 a_11580_15080.n93 a_11580_15080.n92 2.36206
R6890 a_11580_15080.n44 a_11580_15080.n35 2.36206
R6891 a_11580_15080.n56 a_11580_15080.n55 2.36206
R6892 a_11580_15080.n104 a_11580_15080.n103 2.19742
R6893 a_11580_15080.n91 a_11580_15080.n90 2.19742
R6894 a_11580_15080.n46 a_11580_15080.n45 2.19742
R6895 a_11580_15080.n58 a_11580_15080.n57 2.19742
R6896 a_11580_15080.n111 a_11580_15080.n110 1.80838
R6897 a_11580_15080.n39 a_11580_15080.n37 1.80838
R6898 a_11580_15080.n84 a_11580_15080.n17 1.56363
R6899 a_11580_15080.n26 a_11580_15080.n24 1.56363
R6900 a_11580_15080.n27 a_11580_15080.n25 1.5505
R6901 a_11580_15080.n62 a_11580_15080.n61 1.5505
R6902 a_11580_15080.n33 a_11580_15080.n32 1.5505
R6903 a_11580_15080.n50 a_11580_15080.n49 1.5505
R6904 a_11580_15080.n52 a_11580_15080.n51 1.5505
R6905 a_11580_15080.n54 a_11580_15080.n29 1.5505
R6906 a_11580_15080.n43 a_11580_15080.n42 1.5505
R6907 a_11580_15080.n37 a_11580_15080.n36 1.5505
R6908 a_11580_15080.n89 a_11580_15080.n15 1.5505
R6909 a_11580_15080.n87 a_11580_15080.n86 1.5505
R6910 a_11580_15080.n102 a_11580_15080.n10 1.5505
R6911 a_11580_15080.n100 a_11580_15080.n99 1.5505
R6912 a_11580_15080.n98 a_11580_15080.n97 1.5505
R6913 a_11580_15080.n14 a_11580_15080.n13 1.5505
R6914 a_11580_15080.n110 a_11580_15080.n8 1.5505
R6915 a_11580_15080.n105 a_11580_15080.n9 1.5505
R6916 a_11580_15080.n124 a_11580_15080.n123 1.25468
R6917 a_11580_15080.n109 a_11580_15080.n9 1.25468
R6918 a_11580_15080.n96 a_11580_15080.n14 1.25468
R6919 a_11580_15080.n70 a_11580_15080.n19 1.25468
R6920 a_11580_15080.n42 a_11580_15080.n41 1.25468
R6921 a_11580_15080.n54 a_11580_15080.n53 1.25468
R6922 a_11580_15080.n117 a_11580_15080.n4 1.19225
R6923 a_11580_15080.n103 a_11580_15080.n102 1.19225
R6924 a_11580_15080.n90 a_11580_15080.n89 1.19225
R6925 a_11580_15080.n76 a_11580_15080.n21 1.19225
R6926 a_11580_15080.n46 a_11580_15080.n33 1.19225
R6927 a_11580_15080.n58 a_11580_15080.n27 1.19225
R6928 a_11580_15080.n120 a_11580_15080.n5 1.07024
R6929 a_11580_15080.n97 a_11580_15080.n12 1.07024
R6930 a_11580_15080.n72 a_11580_15080.n22 1.07024
R6931 a_11580_15080.n52 a_11580_15080.n31 1.07024
R6932 a_11580_15080.n39 a_11580_15080.n38 1.04968
R6933 a_11580_15080.n112 a_11580_15080.n111 1.04968
R6934 a_11580_15080.n124 a_11580_15080.n6 1.0237
R6935 a_11580_15080.n107 a_11580_15080.n9 1.0237
R6936 a_11580_15080.n93 a_11580_15080.n14 1.0237
R6937 a_11580_15080.n23 a_11580_15080.n19 1.0237
R6938 a_11580_15080.n42 a_11580_15080.n35 1.0237
R6939 a_11580_15080.n55 a_11580_15080.n54 1.0237
R6940 a_11580_15080.n118 a_11580_15080.n4 0.959578
R6941 a_11580_15080.n102 a_11580_15080.n101 0.959578
R6942 a_11580_15080.n89 a_11580_15080.n88 0.959578
R6943 a_11580_15080.n74 a_11580_15080.n21 0.959578
R6944 a_11580_15080.n48 a_11580_15080.n33 0.959578
R6945 a_11580_15080.n60 a_11580_15080.n27 0.959578
R6946 a_11580_15080.n118 a_11580_15080.n2 0.885803
R6947 a_11580_15080.n101 a_11580_15080.n100 0.885803
R6948 a_11580_15080.n88 a_11580_15080.n87 0.885803
R6949 a_11580_15080.n74 a_11580_15080.n20 0.885803
R6950 a_11580_15080.n49 a_11580_15080.n48 0.885803
R6951 a_11580_15080.n61 a_11580_15080.n60 0.885803
R6952 a_11580_15080.n127 a_11580_15080.n6 0.812055
R6953 a_11580_15080.n81 a_11580_15080.n23 0.812055
R6954 a_11580_15080.n120 a_11580_15080.n2 0.77514
R6955 a_11580_15080.n100 a_11580_15080.n12 0.77514
R6956 a_11580_15080.n87 a_11580_15080.n17 0.77514
R6957 a_11580_15080.n72 a_11580_15080.n20 0.77514
R6958 a_11580_15080.n49 a_11580_15080.n31 0.77514
R6959 a_11580_15080.n61 a_11580_15080.n26 0.77514
R6960 a_11580_15080.n117 a_11580_15080.n3 0.647417
R6961 a_11580_15080.n77 a_11580_15080.n76 0.647417
R6962 a_11580_15080.n123 a_11580_15080.n5 0.590702
R6963 a_11580_15080.n110 a_11580_15080.n109 0.590702
R6964 a_11580_15080.n97 a_11580_15080.n96 0.590702
R6965 a_11580_15080.n70 a_11580_15080.n22 0.590702
R6966 a_11580_15080.n41 a_11580_15080.n37 0.590702
R6967 a_11580_15080.n53 a_11580_15080.n52 0.590702
R6968 a_11580_15080.n63 a_11580_15080.n24 0.530034
R6969 a_11580_15080.n85 a_11580_15080.n84 0.530034
R6970 a_11580_15080.t6 a_11580_15080.n121 0.290206
R6971 a_11580_15080.t7 a_11580_15080.n94 0.290206
R6972 a_11580_15080.t4 a_11580_15080.n83 0.290206
R6973 a_11580_15080.n73 a_11580_15080.t2 0.290206
R6974 a_11580_15080.n34 a_11580_15080.t5 0.290206
R6975 a_11580_15080.n28 a_11580_15080.t3 0.290206
R6976 a_11580_15080.n57 a_11580_15080.n56 0.154071
R6977 a_11580_15080.n45 a_11580_15080.n44 0.154071
R6978 a_11580_15080.n92 a_11580_15080.n91 0.154071
R6979 a_11580_15080.n106 a_11580_15080.n104 0.154071
R6980 a_11580_15080.n85 a_11580_15080.n82 0.137464
R6981 a_11580_15080.n113 a_11580_15080.n112 0.137464
R6982 a_11580_15080.n64 a_11580_15080.n63 0.134964
R6983 a_11580_15080.n38 a_11580_15080.n7 0.134964
R6984 a_11580_15080.n62 a_11580_15080.n25 0.0183571
R6985 a_11580_15080.n57 a_11580_15080.n25 0.0183571
R6986 a_11580_15080.n56 a_11580_15080.n29 0.0183571
R6987 a_11580_15080.n51 a_11580_15080.n29 0.0183571
R6988 a_11580_15080.n51 a_11580_15080.n50 0.0183571
R6989 a_11580_15080.n50 a_11580_15080.n32 0.0183571
R6990 a_11580_15080.n45 a_11580_15080.n32 0.0183571
R6991 a_11580_15080.n44 a_11580_15080.n43 0.0183571
R6992 a_11580_15080.n43 a_11580_15080.n36 0.0183571
R6993 a_11580_15080.n86 a_11580_15080.n15 0.0183571
R6994 a_11580_15080.n91 a_11580_15080.n15 0.0183571
R6995 a_11580_15080.n92 a_11580_15080.n13 0.0183571
R6996 a_11580_15080.n98 a_11580_15080.n13 0.0183571
R6997 a_11580_15080.n99 a_11580_15080.n98 0.0183571
R6998 a_11580_15080.n99 a_11580_15080.n10 0.0183571
R6999 a_11580_15080.n104 a_11580_15080.n10 0.0183571
R7000 a_11580_15080.n106 a_11580_15080.n105 0.0183571
R7001 a_11580_15080.n105 a_11580_15080.n8 0.0183571
R7002 a_11580_15080.n38 a_11580_15080.n36 0.0106786
R7003 a_11580_15080.n112 a_11580_15080.n8 0.0106786
R7004 a_11580_15080.n129 a_11580_15080.n0 0.0106786
R7005 a_11580_15080.n69 a_11580_15080.n68 0.00992001
R7006 a_11580_15080.n80 a_11580_15080.n78 0.00992001
R7007 a_11580_15080.n79 a_11580_15080.n65 0.00992001
R7008 a_11580_15080.n67 a_11580_15080.n66 0.00992001
R7009 a_11580_15080.n82 a_11580_15080.n18 0.00992001
R7010 a_11580_15080.n66 a_11580_15080.n65 0.00992001
R7011 a_11580_15080.n67 a_11580_15080.n18 0.00992001
R7012 a_11580_15080.n78 a_11580_15080.n69 0.00992001
R7013 a_11580_15080.n68 a_11580_15080.n64 0.00992001
R7014 a_11580_15080.n80 a_11580_15080.n79 0.00992001
R7015 a_11580_15080.n126 a_11580_15080.n116 0.00992001
R7016 a_11580_15080.n125 a_11580_15080.n0 0.00992001
R7017 a_11580_15080.n115 a_11580_15080.n1 0.00992001
R7018 a_11580_15080.n114 a_11580_15080.n113 0.00992001
R7019 a_11580_15080.n128 a_11580_15080.n1 0.00992001
R7020 a_11580_15080.n115 a_11580_15080.n114 0.00992001
R7021 a_11580_15080.n126 a_11580_15080.n125 0.00992001
R7022 a_11580_15080.n116 a_11580_15080.n7 0.00992001
R7023 a_11580_15080.n63 a_11580_15080.n62 0.00817857
R7024 a_11580_15080.n86 a_11580_15080.n85 0.00817857
R7025 a_11580_15080.n129 a_11580_15080.n128 0.00817857
R7026 a_20810_11490.n1 a_20810_11490.t6 401.668
R7027 a_20810_11490.n5 a_20810_11490.n4 297.394
R7028 a_20810_11490.n3 a_20810_11490.t2 252.248
R7029 a_20810_11490.n2 a_20810_11490.n1 208.868
R7030 a_20810_11490.n4 a_20810_11490.n0 195.582
R7031 a_20810_11490.n1 a_20810_11490.t7 192.8
R7032 a_20810_11490.n2 a_20810_11490.t0 192.8
R7033 a_20810_11490.n4 a_20810_11490.n3 161.3
R7034 a_20810_11490.n0 a_20810_11490.t4 60.0005
R7035 a_20810_11490.n0 a_20810_11490.t5 60.0005
R7036 a_20810_11490.n3 a_20810_11490.n2 59.4472
R7037 a_20810_11490.n5 a_20810_11490.t1 49.2505
R7038 a_20810_11490.t3 a_20810_11490.n5 49.2505
R7039 a_14860_6060.n1 a_14860_6060.t4 562.333
R7040 a_14860_6060.t0 a_14860_6060.n4 500.086
R7041 a_14860_6060.t0 a_14860_6060.n4 461.389
R7042 a_14860_6060.n2 a_14860_6060.n1 453.315
R7043 a_14860_6060.n0 a_14860_6060.t5 417.733
R7044 a_14860_6060.n2 a_14860_6060.n0 388.639
R7045 a_14860_6060.n0 a_14860_6060.t3 369.534
R7046 a_14860_6060.n1 a_14860_6060.t2 224.934
R7047 a_14860_6060.n3 a_14860_6060.t1 172.458
R7048 a_14860_6060.n4 a_14860_6060.n3 43.2699
R7049 a_14860_6060.n3 a_14860_6060.n2 13.4217
R7050 a_14340_6060.n0 a_14340_6060.t3 517.347
R7051 a_14340_6060.n2 a_14340_6060.n0 417.574
R7052 a_14340_6060.n2 a_14340_6060.n1 244.716
R7053 a_14340_6060.n0 a_14340_6060.t4 228.148
R7054 a_14340_6060.t2 a_14340_6060.n2 221.411
R7055 a_14340_6060.n1 a_14340_6060.t0 24.0005
R7056 a_14340_6060.n1 a_14340_6060.t1 24.0005
R7057 a_20830_3320.n0 a_20830_3320.t1 713.933
R7058 a_20830_3320.t0 a_20830_3320.n0 337
R7059 a_20830_3320.n0 a_20830_3320.t2 314.233
R7060 a_21130_3020.t0 a_21130_3020.t1 96.0005
R7061 a_23718_2840.n0 a_23718_2840.t0 135.569
R7062 a_23718_2840.t1 a_23718_2840.n0 135.492
R7063 a_23718_2840.t2 a_23718_2840.n0 80.7139
R7064 a_19910_3400.t5 a_19910_3400.t4 1012.2
R7065 a_19910_3400.n0 a_19910_3400.t1 663.801
R7066 a_19910_3400.n2 a_19910_3400.n1 431.401
R7067 a_19910_3400.t2 a_19910_3400.t3 401.668
R7068 a_19910_3400.n0 a_19910_3400.t5 361.692
R7069 a_19910_3400.n1 a_19910_3400.t6 353.467
R7070 a_19910_3400.t0 a_19910_3400.n2 298.921
R7071 a_19910_3400.n1 a_19910_3400.t2 257.067
R7072 a_19910_3400.n2 a_19910_3400.n0 67.2005
R7073 a_19210_3370.n4 a_19210_3370.t1 752.333
R7074 a_19210_3370.t2 a_19210_3370.n5 752.333
R7075 a_19210_3370.n0 a_19210_3370.t4 514.134
R7076 a_19210_3370.n3 a_19210_3370.n2 366.856
R7077 a_19210_3370.n5 a_19210_3370.t0 254.333
R7078 a_19210_3370.n3 a_19210_3370.t7 190.123
R7079 a_19210_3370.n4 a_19210_3370.n3 187.201
R7080 a_19210_3370.n2 a_19210_3370.n1 176.733
R7081 a_19210_3370.n1 a_19210_3370.n0 176.733
R7082 a_19210_3370.n0 a_19210_3370.t6 112.468
R7083 a_19210_3370.n1 a_19210_3370.t3 112.468
R7084 a_19210_3370.n2 a_19210_3370.t5 112.468
R7085 a_19210_3370.n5 a_19210_3370.n4 70.4005
R7086 a_17400_3080.n1 a_17400_3080.n0 701.467
R7087 a_17400_3080.n1 a_17400_3080.t1 694.201
R7088 a_17400_3080.n0 a_17400_3080.t3 321.334
R7089 a_17400_3080.t0 a_17400_3080.n1 314.921
R7090 a_17400_3080.n0 a_17400_3080.t2 144.601
R7091 a_16960_3370.n0 a_16960_3370.t1 685.134
R7092 a_16960_3370.n1 a_16960_3370.t0 663.801
R7093 a_16960_3370.n0 a_16960_3370.t3 534.268
R7094 a_16960_3370.t2 a_16960_3370.n1 362.921
R7095 a_16960_3370.n1 a_16960_3370.n0 91.7338
R7096 a_19120_3150.n0 a_19120_3150.t3 750.201
R7097 a_19120_3150.n1 a_19120_3150.t4 349.433
R7098 a_19120_3150.n0 a_19120_3150.t1 276.733
R7099 a_19120_3150.n2 a_19120_3150.n1 206.333
R7100 a_19120_3150.n1 a_19120_3150.n0 48.0005
R7101 a_19120_3150.t2 a_19120_3150.n2 48.0005
R7102 a_19120_3150.n2 a_19120_3150.t0 48.0005
R7103 a_18610_3400.t5 a_18610_3400.t2 1012.2
R7104 a_18610_3400.n0 a_18610_3400.t0 663.801
R7105 a_18610_3400.n2 a_18610_3400.n1 431.401
R7106 a_18610_3400.t6 a_18610_3400.t3 401.668
R7107 a_18610_3400.n0 a_18610_3400.t5 361.692
R7108 a_18610_3400.t1 a_18610_3400.n2 298.921
R7109 a_18610_3400.n1 a_18610_3400.t6 257.067
R7110 a_18610_3400.n1 a_18610_3400.t4 208.868
R7111 a_18610_3400.n2 a_18610_3400.n0 67.2005
R7112 a_23198_3560.n0 a_23198_3560.t0 236.867
R7113 a_23198_3560.n0 a_23198_3560.t2 237.337
R7114 a_23198_3560.t1 a_23198_3560.n0 209.882
R7115 a_12620_3080.n4 a_12620_3080.t0 777.4
R7116 a_12620_3080.t6 a_12620_3080.t10 514.134
R7117 a_12620_3080.n3 a_12620_3080.n2 364.178
R7118 a_12620_3080.n0 a_12620_3080.t11 353.467
R7119 a_12620_3080.t4 a_12620_3080.n5 353.467
R7120 a_12620_3080.n6 a_12620_3080.t4 318.702
R7121 a_12620_3080.n6 a_12620_3080.t6 307.909
R7122 a_12620_3080.n5 a_12620_3080.t9 289.2
R7123 a_12620_3080.n4 a_12620_3080.n3 257.079
R7124 a_12620_3080.t1 a_12620_3080.n7 233
R7125 a_12620_3080.n0 a_12620_3080.t3 192.8
R7126 a_12620_3080.n2 a_12620_3080.n1 176.733
R7127 a_12620_3080.n1 a_12620_3080.t8 112.468
R7128 a_12620_3080.n2 a_12620_3080.t2 112.468
R7129 a_12620_3080.n3 a_12620_3080.t5 112.468
R7130 a_12620_3080.n5 a_12620_3080.t7 112.468
R7131 a_12620_3080.n1 a_12620_3080.n0 96.4005
R7132 a_12620_3080.n7 a_12620_3080.n6 38.2642
R7133 a_12620_3080.n7 a_12620_3080.n4 21.3338
R7134 a_12490_3240.n2 a_12490_3240.t3 761.4
R7135 a_12490_3240.n1 a_12490_3240.t4 349.433
R7136 a_12490_3240.t2 a_12490_3240.n2 254.333
R7137 a_12490_3240.n1 a_12490_3240.n0 206.333
R7138 a_12490_3240.n2 a_12490_3240.n1 70.4005
R7139 a_12490_3240.n0 a_12490_3240.t0 48.0005
R7140 a_12490_3240.n0 a_12490_3240.t1 48.0005
R7141 a_13960_7240.n4 a_13960_7240.n0 1319.38
R7142 a_13960_7240.n0 a_13960_7240.t4 562.333
R7143 a_13960_7240.n2 a_13960_7240.t6 388.813
R7144 a_13960_7240.n2 a_13960_7240.t5 356.68
R7145 a_13960_7240.n3 a_13960_7240.n2 232
R7146 a_13960_7240.n0 a_13960_7240.t3 224.934
R7147 a_13960_7240.t1 a_13960_7240.n4 221.411
R7148 a_13960_7240.n3 a_13960_7240.n1 157.278
R7149 a_13960_7240.n4 a_13960_7240.n3 90.64
R7150 a_13960_7240.n1 a_13960_7240.t0 24.0005
R7151 a_13960_7240.n1 a_13960_7240.t2 24.0005
R7152 a_14340_7240.n0 a_14340_7240.t4 517.347
R7153 a_14340_7240.n2 a_14340_7240.n0 417.574
R7154 a_14340_7240.n2 a_14340_7240.n1 244.716
R7155 a_14340_7240.n0 a_14340_7240.t3 228.148
R7156 a_14340_7240.t2 a_14340_7240.n2 221.411
R7157 a_14340_7240.n1 a_14340_7240.t0 24.0005
R7158 a_14340_7240.n1 a_14340_7240.t1 24.0005
R7159 a_13540_3080.n2 a_13540_3080.t3 723.534
R7160 a_13540_3080.n1 a_13540_3080.t4 553.534
R7161 a_13540_3080.t2 a_13540_3080.n2 254.333
R7162 a_13540_3080.n1 a_13540_3080.n0 206.333
R7163 a_13540_3080.n2 a_13540_3080.n1 70.4005
R7164 a_13540_3080.n0 a_13540_3080.t0 48.0005
R7165 a_13540_3080.n0 a_13540_3080.t1 48.0005
R7166 a_19930_11490.n3 a_19930_11490.t6 377.567
R7167 a_19930_11490.n2 a_19930_11490.t9 297.233
R7168 a_19930_11490.n4 a_19930_11490.n2 231.575
R7169 a_19930_11490.n4 a_19930_11490.n3 228.778
R7170 a_19930_11490.n3 a_19930_11490.t8 216.9
R7171 a_19930_11490.n0 a_19930_11490.n5 153.401
R7172 a_19930_11490.n6 a_19930_11490.n0 153.4
R7173 a_19930_11490.n2 a_19930_11490.t7 136.567
R7174 a_19930_11490.n0 a_19930_11490.n1 54.9641
R7175 a_19930_11490.n5 a_19930_11490.t0 24.6255
R7176 a_19930_11490.n5 a_19930_11490.t2 24.6255
R7177 a_19930_11490.t3 a_19930_11490.n6 24.6255
R7178 a_19930_11490.n6 a_19930_11490.t1 24.6255
R7179 a_19930_11490.n0 a_19930_11490.n4 21.3599
R7180 a_19930_11490.n1 a_19930_11490.t5 15.0005
R7181 a_19930_11490.n1 a_19930_11490.t4 15.0005
R7182 a_19830_3020.t0 a_19830_3020.t1 96.0005
R7183 a_19690_10220.n1 a_19690_10220.t0 476.896
R7184 a_19690_10220.n7 a_19690_10220.t11 317.317
R7185 a_19690_10220.n2 a_19690_10220.t10 317.317
R7186 a_19690_10220.n8 a_19690_10220.n7 257.067
R7187 a_19690_10220.n6 a_19690_10220.n5 257.067
R7188 a_19690_10220.n3 a_19690_10220.n2 257.067
R7189 a_19690_10220.n4 a_19690_10220.n1 152
R7190 a_19690_10220.n10 a_19690_10220.n9 152
R7191 a_19690_10220.n1 a_19690_10220.n0 123.469
R7192 a_19690_10220.n11 a_19690_10220.n10 117.781
R7193 a_19690_10220.n9 a_19690_10220.n8 85.6894
R7194 a_19690_10220.n9 a_19690_10220.n6 85.6894
R7195 a_19690_10220.n5 a_19690_10220.n4 85.6894
R7196 a_19690_10220.n4 a_19690_10220.n3 85.6894
R7197 a_19690_10220.n7 a_19690_10220.t9 60.2505
R7198 a_19690_10220.n8 a_19690_10220.t5 60.2505
R7199 a_19690_10220.n6 a_19690_10220.t7 60.2505
R7200 a_19690_10220.n5 a_19690_10220.t1 60.2505
R7201 a_19690_10220.n2 a_19690_10220.t12 60.2505
R7202 a_19690_10220.n3 a_19690_10220.t3 60.2505
R7203 a_19690_10220.n10 a_19690_10220.n1 56.0005
R7204 a_19690_10220.n0 a_19690_10220.t4 24.0005
R7205 a_19690_10220.n0 a_19690_10220.t2 24.0005
R7206 a_19690_10220.t8 a_19690_10220.n11 24.0005
R7207 a_19690_10220.n11 a_19690_10220.t6 24.0005
R7208 a_12520_10060.n4 a_12520_10060.n3 314.526
R7209 a_12520_10060.n5 a_12520_10060.t11 287.762
R7210 a_12520_10060.n6 a_12520_10060.t8 287.762
R7211 a_12520_10060.n5 a_12520_10060.t10 287.589
R7212 a_12520_10060.n7 a_12520_10060.t12 287.012
R7213 a_12520_10060.n8 a_12520_10060.t9 287.012
R7214 a_12520_10060.n2 a_12520_10060.n0 107.079
R7215 a_12520_10060.n2 a_12520_10060.n1 104.829
R7216 a_12520_10060.t0 a_12520_10060.n10 49.8165
R7217 a_12520_10060.n10 a_12520_10060.t3 44.8391
R7218 a_12520_10060.n3 a_12520_10060.t2 39.4005
R7219 a_12520_10060.n3 a_12520_10060.t1 39.4005
R7220 a_12520_10060.n0 a_12520_10060.t6 13.1338
R7221 a_12520_10060.n0 a_12520_10060.t7 13.1338
R7222 a_12520_10060.n1 a_12520_10060.t4 13.1338
R7223 a_12520_10060.n1 a_12520_10060.t5 13.1338
R7224 a_12520_10060.n10 a_12520_10060.n9 11.8755
R7225 a_12520_10060.n9 a_12520_10060.n4 10.7505
R7226 a_12520_10060.n9 a_12520_10060.n8 6.78086
R7227 a_12520_10060.n4 a_12520_10060.n2 2.0005
R7228 a_12520_10060.n7 a_12520_10060.n6 0.579071
R7229 a_12520_10060.n8 a_12520_10060.n7 0.282643
R7230 a_12520_10060.n6 a_12520_10060.n5 0.2755
R7231 a_21720_3150.n2 a_21720_3150.t3 750.201
R7232 a_21720_3150.n1 a_21720_3150.t4 349.433
R7233 a_21720_3150.t2 a_21720_3150.n2 276.733
R7234 a_21720_3150.n1 a_21720_3150.n0 206.333
R7235 a_21720_3150.n0 a_21720_3150.t1 48.0005
R7236 a_21720_3150.n0 a_21720_3150.t0 48.0005
R7237 a_21720_3150.n2 a_21720_3150.n1 48.0005
R7238 a_19244_9974.n0 a_19244_9974.t0 477.969
R7239 a_19244_9974.n8 a_19244_9974.t10 377.567
R7240 a_19244_9974.n1 a_19244_9974.t9 377.567
R7241 a_19244_9974.n9 a_19244_9974.n8 257.067
R7242 a_19244_9974.n7 a_19244_9974.n6 257.067
R7243 a_19244_9974.n2 a_19244_9974.n1 257.067
R7244 a_19244_9974.n5 a_19244_9974.n4 161.3
R7245 a_19244_9974.n11 a_19244_9974.n10 161.3
R7246 a_19244_9974.n8 a_19244_9974.t12 120.501
R7247 a_19244_9974.n9 a_19244_9974.t3 120.501
R7248 a_19244_9974.n7 a_19244_9974.t5 120.501
R7249 a_19244_9974.n6 a_19244_9974.t7 120.501
R7250 a_19244_9974.n1 a_19244_9974.t11 120.501
R7251 a_19244_9974.n2 a_19244_9974.t1 120.501
R7252 a_19244_9974.n4 a_19244_9974.n3 119.237
R7253 a_19244_9974.n12 a_19244_9974.n11 119.237
R7254 a_19244_9974.n10 a_19244_9974.n9 85.6894
R7255 a_19244_9974.n10 a_19244_9974.n7 85.6894
R7256 a_19244_9974.n6 a_19244_9974.n5 85.6894
R7257 a_19244_9974.n5 a_19244_9974.n2 85.6894
R7258 a_19244_9974.n3 a_19244_9974.t2 19.7005
R7259 a_19244_9974.n3 a_19244_9974.t8 19.7005
R7260 a_19244_9974.t6 a_19244_9974.n12 19.7005
R7261 a_19244_9974.n12 a_19244_9974.t4 19.7005
R7262 a_19244_9974.n4 a_19244_9974.n0 5.1255
R7263 a_19244_9974.n11 a_19244_9974.n0 4.5005
R7264 a_23198_2840.n0 a_23198_2840.t0 135.569
R7265 a_23198_2840.t1 a_23198_2840.n0 135.492
R7266 a_23198_2840.t2 a_23198_2840.n0 80.7139
R7267 a_15300_6090.t0 a_15300_6090.t1 48.0005
R7268 a_23280_5000.n1 a_23280_5000.t1 247.257
R7269 a_23280_5000.n0 a_23280_5000.t2 240.543
R7270 a_23280_5000.n0 a_23280_5000.t5 198.746
R7271 a_23280_5000.n0 a_23280_5000.t3 197.934
R7272 a_23280_5000.n0 a_23280_5000.t4 197.934
R7273 a_23280_5000.t0 a_23280_5000.n1 140.6
R7274 a_23280_5000.n1 a_23280_5000.n0 6.1255
R7275 a_13360_6090.n2 a_13360_6090.n0 1319.38
R7276 a_13360_6090.t6 a_13360_6090.t5 1188.93
R7277 a_13360_6090.t5 a_13360_6090.t3 835.467
R7278 a_13360_6090.n0 a_13360_6090.t4 562.333
R7279 a_13360_6090.n2 a_13360_6090.n1 247.917
R7280 a_13360_6090.n0 a_13360_6090.t6 224.934
R7281 a_13360_6090.t1 a_13360_6090.n2 221.411
R7282 a_13360_6090.n1 a_13360_6090.t2 24.0005
R7283 a_13360_6090.n1 a_13360_6090.t0 24.0005
R7284 a_14260_6510.t0 a_14260_6510.t1 39.4005
R7285 a_15740_6090.t1 a_15740_6090.n2 500.086
R7286 a_15740_6090.n1 a_15740_6090.n0 473.334
R7287 a_15740_6090.n0 a_15740_6090.t2 465.933
R7288 a_15740_6090.t1 a_15740_6090.n2 461.389
R7289 a_15740_6090.n0 a_15740_6090.t3 321.334
R7290 a_15740_6090.n1 a_15740_6090.t0 177.577
R7291 a_15740_6090.n2 a_15740_6090.n1 48.3898
R7292 a_15920_7240.n0 a_15920_7240.t3 465.933
R7293 a_15920_7240.n1 a_15920_7240.n0 431.824
R7294 a_15920_7240.n0 a_15920_7240.t2 321.334
R7295 a_15920_7240.t1 a_15920_7240.n1 288.37
R7296 a_15920_7240.n1 a_15920_7240.t0 177.577
R7297 a_20420_3150.n0 a_20420_3150.t3 750.201
R7298 a_20420_3150.n1 a_20420_3150.t4 349.433
R7299 a_20420_3150.n0 a_20420_3150.t1 276.733
R7300 a_20420_3150.n2 a_20420_3150.n1 206.333
R7301 a_20420_3150.n1 a_20420_3150.n0 48.0005
R7302 a_20420_3150.t2 a_20420_3150.n2 48.0005
R7303 a_20420_3150.n2 a_20420_3150.t0 48.0005
R7304 a_19790_10270.n7 a_19790_10270.n5 482.582
R7305 a_19790_10270.n10 a_19790_10270.t4 304.634
R7306 a_19790_10270.n3 a_19790_10270.t2 304.634
R7307 a_19790_10270.t6 a_19790_10270.n10 279.134
R7308 a_19790_10270.n3 a_19790_10270.t3 277
R7309 a_19790_10270.n8 a_19790_10270.n1 204.201
R7310 a_19790_10270.n4 a_19790_10270.n2 204.201
R7311 a_19790_10270.n9 a_19790_10270.n0 204.201
R7312 a_19790_10270.n7 a_19790_10270.n6 120.981
R7313 a_19790_10270.n8 a_19790_10270.n4 74.6672
R7314 a_19790_10270.n9 a_19790_10270.n8 74.6672
R7315 a_19790_10270.n1 a_19790_10270.t0 60.0005
R7316 a_19790_10270.n1 a_19790_10270.t7 60.0005
R7317 a_19790_10270.t3 a_19790_10270.n2 60.0005
R7318 a_19790_10270.n2 a_19790_10270.t1 60.0005
R7319 a_19790_10270.n0 a_19790_10270.t8 60.0005
R7320 a_19790_10270.n0 a_19790_10270.t5 60.0005
R7321 a_19790_10270.n8 a_19790_10270.n7 28.5443
R7322 a_19790_10270.n5 a_19790_10270.t12 24.0005
R7323 a_19790_10270.n5 a_19790_10270.t10 24.0005
R7324 a_19790_10270.n6 a_19790_10270.t11 24.0005
R7325 a_19790_10270.n6 a_19790_10270.t9 24.0005
R7326 a_19790_10270.n4 a_19790_10270.n3 16.0005
R7327 a_19790_10270.n10 a_19790_10270.n9 16.0005
R7328 a_23224_12716.t1 a_23224_12716.t0 51.4199
R7329 a_19530_3320.n0 a_19530_3320.t0 713.933
R7330 a_19530_3320.t1 a_19530_3320.n0 337
R7331 a_19530_3320.n0 a_19530_3320.t2 314.233
R7332 a_24238_2840.n0 a_24238_2840.t1 135.569
R7333 a_24238_2840.t0 a_24238_2840.n0 135.492
R7334 a_24238_2840.t2 a_24238_2840.n0 80.7139
R7335 a_19960_10960.t0 a_19960_10960.n6 857.211
R7336 a_19960_10960.n2 a_19960_10960.n0 297.988
R7337 a_19960_10960.n3 a_19960_10960.n2 264.61
R7338 a_19960_10960.n3 a_19960_10960.t7 208.868
R7339 a_19960_10960.n4 a_19960_10960.t8 208.868
R7340 a_19960_10960.n5 a_19960_10960.t5 208.868
R7341 a_19960_10960.n6 a_19960_10960.t6 208.868
R7342 a_19960_10960.n6 a_19960_10960.n5 208.868
R7343 a_19960_10960.n5 a_19960_10960.n4 208.868
R7344 a_19960_10960.n4 a_19960_10960.n3 208.868
R7345 a_19960_10960.n2 a_19960_10960.n1 195.035
R7346 a_19960_10960.n1 a_19960_10960.t4 60.0005
R7347 a_19960_10960.n1 a_19960_10960.t3 60.0005
R7348 a_19960_10960.n0 a_19960_10960.t1 49.2505
R7349 a_19960_10960.n0 a_19960_10960.t2 49.2505
R7350 a_13880_6510.t0 a_13880_6510.t1 39.4005
R7351 a_14860_3240.n0 a_14860_3240.t0 761.4
R7352 a_14860_3240.n1 a_14860_3240.t4 350.349
R7353 a_14860_3240.n0 a_14860_3240.t2 254.333
R7354 a_14860_3240.n2 a_14860_3240.n1 206.333
R7355 a_14860_3240.n1 a_14860_3240.n0 70.4005
R7356 a_14860_3240.n2 a_14860_3240.t1 48.0005
R7357 a_14860_3240.t3 a_14860_3240.n2 48.0005
R7358 a_13360_7890.n2 a_13360_7890.n0 1319.38
R7359 a_13360_7890.t6 a_13360_7890.t5 1188.93
R7360 a_13360_7890.t5 a_13360_7890.t3 835.467
R7361 a_13360_7890.n0 a_13360_7890.t4 562.333
R7362 a_13360_7890.n2 a_13360_7890.n1 247.917
R7363 a_13360_7890.n0 a_13360_7890.t6 224.934
R7364 a_13360_7890.t0 a_13360_7890.n2 221.411
R7365 a_13360_7890.n1 a_13360_7890.t1 24.0005
R7366 a_13360_7890.n1 a_13360_7890.t2 24.0005
R7367 a_14260_7270.t0 a_14260_7270.t1 39.4005
R7368 a_15380_3110.n0 a_15380_3110.t0 663.801
R7369 a_15380_3110.t1 a_15380_3110.n0 397.053
R7370 a_15380_3110.n0 a_15380_3110.t2 348.851
R7371 a_15490_3110.t0 a_15490_3110.t1 96.0005
R7372 a_15260_7240.t1 a_15260_7240.n2 500.086
R7373 a_15260_7240.n1 a_15260_7240.n0 473.334
R7374 a_15260_7240.n0 a_15260_7240.t2 465.933
R7375 a_15260_7240.t1 a_15260_7240.n2 461.389
R7376 a_15260_7240.n0 a_15260_7240.t3 321.334
R7377 a_15260_7240.n1 a_15260_7240.t0 177.577
R7378 a_15260_7240.n2 a_15260_7240.n1 48.3899
R7379 a_22130_3320.n0 a_22130_3320.t0 713.933
R7380 a_22130_3320.t1 a_22130_3320.n0 337
R7381 a_22130_3320.n0 a_22130_3320.t2 314.233
R7382 a_13880_7270.t0 a_13880_7270.t1 39.4005
R7383 a_22430_3020.t0 a_22430_3020.t1 96.0005
R7384 a_11160_14080.n0 a_11160_14080.t7 238.322
R7385 a_11160_14080.n0 a_11160_14080.t6 238.322
R7386 a_11160_14080.n4 a_11160_14080.n0 168.8
R7387 a_11160_14080.n1 a_11160_14080.t1 130.001
R7388 a_11160_14080.n3 a_11160_14080.n2 105.171
R7389 a_11160_14080.n5 a_11160_14080.n4 105.171
R7390 a_11160_14080.n1 a_11160_14080.t0 81.7085
R7391 a_11160_14080.n3 a_11160_14080.n1 48.2927
R7392 a_11160_14080.n2 a_11160_14080.t2 13.1338
R7393 a_11160_14080.n2 a_11160_14080.t4 13.1338
R7394 a_11160_14080.n5 a_11160_14080.t3 13.1338
R7395 a_11160_14080.t5 a_11160_14080.n5 13.1338
R7396 a_11160_14080.n4 a_11160_14080.n3 3.3755
R7397 a_17430_3110.t0 a_17430_3110.t1 96.0005
R7398 a_13240_14080.t0 a_13240_14080.t1 178.194
R7399 a_15570_3080.t2 a_15570_3080.n2 755.534
R7400 a_15570_3080.n2 a_15570_3080.t1 685.134
R7401 a_15570_3080.n1 a_15570_3080.n0 389.733
R7402 a_15570_3080.n1 a_15570_3080.t0 340.2
R7403 a_15570_3080.n0 a_15570_3080.t3 321.334
R7404 a_15570_3080.n0 a_15570_3080.t4 144.601
R7405 a_15570_3080.n2 a_15570_3080.n1 19.2005
R7406 a_14230_3430.t0 a_14230_3430.t1 157.601
R7407 a_15590_7240.t1 a_15590_7240.n2 500.086
R7408 a_15590_7240.n1 a_15590_7240.n0 473.334
R7409 a_15590_7240.n0 a_15590_7240.t3 465.933
R7410 a_15590_7240.t1 a_15590_7240.n2 461.389
R7411 a_15590_7240.n0 a_15590_7240.t2 321.334
R7412 a_15590_7240.n1 a_15590_7240.t0 177.577
R7413 a_15590_7240.n2 a_15590_7240.n1 48.3899
R7414 a_15300_6510.n1 a_15300_6510.n0 481.334
R7415 a_15300_6510.n0 a_15300_6510.t3 465.933
R7416 a_15300_6510.n0 a_15300_6510.t4 321.334
R7417 a_15300_6510.n2 a_15300_6510.n1 226.888
R7418 a_15300_6510.n1 a_15300_6510.t1 172.458
R7419 a_15300_6510.n2 a_15300_6510.t2 19.7005
R7420 a_15300_6510.t0 a_15300_6510.n2 19.7005
R7421 a_14992_19436.t0 a_14992_19436.t1 56.7426
R7422 a_17580_7270.t4 a_17580_7270.t5 377.567
R7423 a_17580_7270.n2 a_17580_7270.n1 237.353
R7424 a_17580_7270.t2 a_17580_7270.n3 229.127
R7425 a_17580_7270.n0 a_17580_7270.t3 220.505
R7426 a_17580_7270.n1 a_17580_7270.n0 196.817
R7427 a_17580_7270.n3 a_17580_7270.t0 158.335
R7428 a_17580_7270.n2 a_17580_7270.t1 151.935
R7429 a_17580_7270.n3 a_17580_7270.n2 121.6
R7430 a_17580_7270.t5 a_17580_7270.n0 92.3838
R7431 a_17580_7270.n1 a_17580_7270.t4 92.3838
R7432 a_13960_6060.n4 a_13960_6060.n0 1319.38
R7433 a_13960_6060.n0 a_13960_6060.t3 562.333
R7434 a_13960_6060.n2 a_13960_6060.t5 388.813
R7435 a_13960_6060.n2 a_13960_6060.t6 356.68
R7436 a_13960_6060.n3 a_13960_6060.n2 232
R7437 a_13960_6060.n0 a_13960_6060.t4 224.934
R7438 a_13960_6060.t0 a_13960_6060.n4 221.411
R7439 a_13960_6060.n3 a_13960_6060.n1 157.278
R7440 a_13960_6060.n4 a_13960_6060.n3 90.64
R7441 a_13960_6060.n1 a_13960_6060.t1 24.0005
R7442 a_13960_6060.n1 a_13960_6060.t2 24.0005
R7443 a_14780_6510.t0 a_14780_6510.t1 39.4005
R7444 a_14780_7270.t0 a_14780_7270.t1 39.4005
R7445 a_13870_3370.n1 a_13870_3370.t2 685.134
R7446 a_13870_3370.n0 a_13870_3370.t1 685.134
R7447 a_13870_3370.n0 a_13870_3370.t3 534.268
R7448 a_13870_3370.t0 a_13870_3370.n1 340.521
R7449 a_13870_3370.n1 a_13870_3370.n0 105.6
R7450 a_23224_9624.t1 a_23224_9624.t0 12.4028
R7451 a_23310_2840.n0 a_23310_2840.t3 537.245
R7452 a_23310_2840.n0 a_23310_2840.t2 386.62
R7453 a_23310_2840.t0 a_23310_2840.n1 236.581
R7454 a_23310_2840.n1 a_23310_2840.t1 135.5
R7455 a_23310_2840.n1 a_23310_2840.n0 3.08327
R7456 a_13010_3110.n0 a_13010_3110.t0 663.801
R7457 a_13010_3110.t1 a_13010_3110.n0 397.053
R7458 a_13010_3110.n0 a_13010_3110.t2 355.378
R7459 a_13120_3110.t0 a_13120_3110.t1 96.0005
R7460 a_18530_3110.t0 a_18530_3110.t1 96.0005
R7461 a_14450_3110.t0 a_14450_3110.t1 96.0005
R7462 a_17320_3110.t0 a_17320_3110.t1 96.0005
C0 VDPWR V_CONT 1.54611f
C1 ua[0] V_CONT 0.05859f
C2 VDPWR ua[0] 0.359818f
C3 ua[1] V_CONT 1.57191f
C4 VDPWR ua[1] 1.51925f
C5 ua[0] ua[1] 0.146073f
C6 I_IN V_CONT 0.036539f
C7 VDPWR I_IN 7.59812f
C8 ua[1] VGND 7.74088f
C9 ua[0] VGND 13.2231f
C10 VDPWR VGND 0.184473p
C11 I_IN VGND 8.42436f
C12 V_CONT VGND 38.928825f
C13 a_14992_19436.t1 VGND 2.19829f
C14 a_11160_14080.t3 VGND 0.041974f
C15 a_11160_14080.t6 VGND 0.015773f
C16 a_11160_14080.t7 VGND 0.015773f
C17 a_11160_14080.n0 VGND 0.051851f
C18 a_11160_14080.t0 VGND 1.67319f
C19 a_11160_14080.t1 VGND 0.043984f
C20 a_11160_14080.n1 VGND 1.51846f
C21 a_11160_14080.t2 VGND 0.041974f
C22 a_11160_14080.t4 VGND 0.041974f
C23 a_11160_14080.n2 VGND 0.103398f
C24 a_11160_14080.n3 VGND 2.32471f
C25 a_11160_14080.n4 VGND 1.18157f
C26 a_11160_14080.n5 VGND 0.103398f
C27 a_11160_14080.t5 VGND 0.041974f
C28 a_23280_5000.n0 VGND 1.03279f
C29 a_23280_5000.t5 VGND 0.49412f
C30 a_23280_5000.t4 VGND 0.493385f
C31 a_23280_5000.t3 VGND 0.493385f
C32 a_23280_5000.t2 VGND 0.093787f
C33 a_23280_5000.t1 VGND 0.487749f
C34 a_23280_5000.n1 VGND 0.832478f
C35 a_23280_5000.t0 VGND 0.072303f
C36 a_19244_9974.t4 VGND 0.037557f
C37 a_19244_9974.t0 VGND 0.07205f
C38 a_19244_9974.n0 VGND 1.121f
C39 a_19244_9974.t5 VGND 0.103656f
C40 a_19244_9974.t7 VGND 0.103656f
C41 a_19244_9974.t1 VGND 0.103656f
C42 a_19244_9974.t11 VGND 0.103656f
C43 a_19244_9974.t9 VGND 0.142523f
C44 a_19244_9974.n1 VGND 0.079812f
C45 a_19244_9974.n2 VGND 0.056635f
C46 a_19244_9974.t2 VGND 0.037557f
C47 a_19244_9974.t8 VGND 0.037557f
C48 a_19244_9974.n3 VGND 0.077646f
C49 a_19244_9974.n4 VGND 0.282214f
C50 a_19244_9974.n5 VGND 0.025445f
C51 a_19244_9974.n6 VGND 0.056635f
C52 a_19244_9974.n7 VGND 0.056635f
C53 a_19244_9974.t3 VGND 0.103656f
C54 a_19244_9974.t12 VGND 0.103656f
C55 a_19244_9974.t10 VGND 0.142523f
C56 a_19244_9974.n8 VGND 0.079812f
C57 a_19244_9974.n9 VGND 0.056635f
C58 a_19244_9974.n10 VGND 0.025445f
C59 a_19244_9974.n11 VGND 0.275179f
C60 a_19244_9974.n12 VGND 0.077646f
C61 a_19244_9974.t6 VGND 0.037557f
C62 a_12520_10060.t6 VGND 0.041299f
C63 a_12520_10060.t7 VGND 0.041299f
C64 a_12520_10060.n0 VGND 0.110485f
C65 a_12520_10060.t4 VGND 0.041299f
C66 a_12520_10060.t5 VGND 0.041299f
C67 a_12520_10060.n1 VGND 0.10021f
C68 a_12520_10060.n2 VGND 1.1329f
C69 a_12520_10060.t2 VGND 0.013766f
C70 a_12520_10060.t1 VGND 0.013766f
C71 a_12520_10060.n3 VGND 0.038807f
C72 a_12520_10060.n4 VGND 0.801094f
C73 a_12520_10060.t10 VGND 0.022789f
C74 a_12520_10060.t11 VGND 0.022325f
C75 a_12520_10060.n5 VGND 0.173944f
C76 a_12520_10060.t8 VGND 0.022325f
C77 a_12520_10060.n6 VGND 0.092865f
C78 a_12520_10060.t12 VGND 0.022626f
C79 a_12520_10060.n7 VGND 0.093528f
C80 a_12520_10060.t9 VGND 0.022626f
C81 a_12520_10060.n8 VGND 0.319446f
C82 a_12520_10060.n9 VGND 0.49355f
C83 a_12520_10060.t3 VGND 3.03225f
C84 a_12520_10060.n10 VGND 4.07807f
C85 a_12520_10060.t0 VGND 0.127426f
C86 a_19930_11490.n0 VGND 1.15801f
C87 a_19930_11490.t5 VGND 0.019782f
C88 a_19930_11490.t4 VGND 0.019782f
C89 a_19930_11490.n1 VGND 0.067671f
C90 a_19930_11490.n2 VGND 0.020139f
C91 a_19930_11490.t6 VGND 0.011563f
C92 a_19930_11490.n3 VGND 0.022197f
C93 a_19930_11490.n4 VGND 0.593f
C94 a_19930_11490.t0 VGND 0.019782f
C95 a_19930_11490.t2 VGND 0.019782f
C96 a_19930_11490.n5 VGND 0.044818f
C97 a_19930_11490.t1 VGND 0.019782f
C98 a_19930_11490.n6 VGND 0.044818f
C99 a_19930_11490.t3 VGND 0.019782f
C100 V_CONT.t7 VGND 7.27996f
C101 V_CONT.t4 VGND 0.026525f
C102 V_CONT.n7 VGND 0.613127f
C103 V_CONT.n13 VGND 0.090296f
C104 V_CONT.n14 VGND 0.348368f
C105 V_CONT.n16 VGND 0.712123f
C106 V_CONT.n18 VGND 0.07073f
C107 V_CONT.n22 VGND 0.039505f
C108 V_CONT.n23 VGND 0.046376f
C109 V_CONT.n24 VGND 0.372467f
C110 V_CONT.n25 VGND 0.017043f
C111 V_CONT.n26 VGND 0.0106f
C112 V_CONT.n27 VGND 0.020036f
C113 a_13440_7240.t5 VGND 0.028262f
C114 a_13440_7240.t6 VGND 0.064454f
C115 a_13440_7240.n0 VGND 0.162805f
C116 a_13440_7240.t7 VGND 0.029978f
C117 a_13440_7240.t3 VGND 0.063823f
C118 a_13440_7240.n1 VGND 0.09612f
C119 a_13440_7240.t4 VGND 0.063823f
C120 a_13440_7240.t8 VGND 0.092852f
C121 a_13440_7240.n2 VGND 1.17335f
C122 a_13440_7240.n3 VGND 0.254916f
C123 a_13440_7240.t2 VGND 0.025787f
C124 a_13440_7240.t0 VGND 0.025787f
C125 a_13440_7240.n4 VGND 0.137692f
C126 a_13440_7240.n5 VGND 0.244629f
C127 a_13440_7240.t1 VGND 0.135725f
C128 a_17290_7270.t1 VGND 0.034319f
C129 a_17290_7270.t0 VGND 1.73994f
C130 a_17290_7270.t3 VGND 0.042516f
C131 a_17290_7270.n0 VGND 0.102101f
C132 a_17290_7270.t2 VGND 0.08112f
C133 a_11431_12690.t10 VGND 0.019608f
C134 a_11431_12690.t7 VGND 0.019608f
C135 a_11431_12690.n0 VGND 0.043211f
C136 a_11431_12690.t1 VGND 0.019608f
C137 a_11431_12690.t4 VGND 0.019608f
C138 a_11431_12690.n1 VGND 0.042942f
C139 a_11431_12690.n2 VGND 0.500119f
C140 a_11431_12690.t9 VGND 0.019608f
C141 a_11431_12690.t3 VGND 0.019608f
C142 a_11431_12690.n3 VGND 0.042942f
C143 a_11431_12690.n4 VGND 0.263919f
C144 a_11431_12690.t8 VGND 0.019608f
C145 a_11431_12690.t2 VGND 0.019608f
C146 a_11431_12690.n5 VGND 0.042942f
C147 a_11431_12690.n6 VGND 0.263919f
C148 a_11431_12690.t6 VGND 0.019608f
C149 a_11431_12690.t5 VGND 0.019608f
C150 a_11431_12690.n7 VGND 0.042942f
C151 a_11431_12690.n8 VGND 0.263919f
C152 a_11431_12690.t0 VGND 0.019608f
C153 a_11431_12690.t11 VGND 0.019608f
C154 a_11431_12690.n9 VGND 0.042942f
C155 a_11431_12690.n10 VGND 1.22448f
C156 a_11431_12690.t13 VGND 0.030146f
C157 a_11431_12690.t16 VGND 0.030088f
C158 a_11431_12690.n11 VGND 0.211627f
C159 a_11431_12690.t15 VGND 0.030088f
C160 a_11431_12690.n12 VGND 0.131578f
C161 a_11431_12690.t17 VGND 0.030088f
C162 a_11431_12690.n13 VGND 0.131578f
C163 a_11431_12690.t14 VGND 0.030088f
C164 a_11431_12690.n14 VGND 0.596207f
C165 a_11431_12690.n15 VGND 3.87358f
C166 a_11431_12690.t12 VGND 2.59536f
C167 a_17574_18026.t1 VGND 0.304962f
C168 a_17574_18026.t4 VGND 0.321329f
C169 a_17574_18026.t9 VGND 0.321329f
C170 a_17574_18026.t2 VGND 0.321329f
C171 a_17574_18026.t5 VGND 0.321329f
C172 a_17574_18026.t20 VGND 0.321329f
C173 a_17574_18026.t17 VGND 0.321329f
C174 a_17574_18026.t10 VGND 0.321329f
C175 a_17574_18026.t14 VGND 0.306067f
C176 a_17574_18026.t7 VGND 0.147435f
C177 a_17574_18026.n0 VGND 0.190169f
C178 a_17574_18026.t13 VGND 0.334291f
C179 a_17574_18026.t18 VGND 0.307353f
C180 a_17574_18026.t16 VGND 0.321329f
C181 a_17574_18026.t19 VGND 0.321329f
C182 a_17574_18026.t3 VGND 0.321329f
C183 a_17574_18026.t12 VGND 0.321329f
C184 a_17574_18026.t8 VGND 0.321329f
C185 a_17574_18026.t15 VGND 0.321329f
C186 a_17574_18026.t11 VGND 0.321329f
C187 a_17574_18026.t6 VGND 0.937937f
C188 a_17574_18026.t0 VGND 0.173184f
C189 a_10840_11590.t5 VGND 0.02f
C190 a_10840_11590.t19 VGND 0.02f
C191 a_10840_11590.t22 VGND 0.032283f
C192 a_10840_11590.n0 VGND 0.036051f
C193 a_10840_11590.n1 VGND 0.024627f
C194 a_10840_11590.t13 VGND 0.025389f
C195 a_10840_11590.n2 VGND 0.039854f
C196 a_10840_11590.t6 VGND 0.016667f
C197 a_10840_11590.t14 VGND 0.016667f
C198 a_10840_11590.n3 VGND 0.034125f
C199 a_10840_11590.n4 VGND 0.176664f
C200 a_10840_11590.n5 VGND 0.017774f
C201 a_10840_11590.t4 VGND 0.031554f
C202 a_10840_11590.n6 VGND 0.019781f
C203 a_10840_11590.n7 VGND 0.511999f
C204 a_10840_11590.n8 VGND 0.172226f
C205 a_10840_11590.t7 VGND 0.02f
C206 a_10840_11590.t21 VGND 0.02f
C207 a_10840_11590.t17 VGND 0.032283f
C208 a_10840_11590.n9 VGND 0.036051f
C209 a_10840_11590.n10 VGND 0.024627f
C210 a_10840_11590.t11 VGND 0.025389f
C211 a_10840_11590.n11 VGND 0.039854f
C212 a_10840_11590.t8 VGND 0.016667f
C213 a_10840_11590.t12 VGND 0.016667f
C214 a_10840_11590.n12 VGND 0.034125f
C215 a_10840_11590.n13 VGND 0.221004f
C216 a_10840_11590.n14 VGND 0.242013f
C217 a_10840_11590.t15 VGND 0.02f
C218 a_10840_11590.t20 VGND 0.02f
C219 a_10840_11590.t18 VGND 0.032283f
C220 a_10840_11590.n15 VGND 0.036051f
C221 a_10840_11590.n16 VGND 0.024627f
C222 a_10840_11590.t9 VGND 0.025389f
C223 a_10840_11590.n17 VGND 0.039854f
C224 a_10840_11590.n18 VGND 0.176664f
C225 a_10840_11590.t10 VGND 0.016667f
C226 a_10840_11590.n19 VGND 0.034125f
C227 a_10840_11590.t16 VGND 0.016667f
C228 a_9573_16817.t5 VGND 0.08597f
C229 a_9573_16817.t2 VGND 0.08597f
C230 a_9573_16817.n0 VGND 0.239812f
C231 a_9573_16817.t4 VGND 0.08597f
C232 a_9573_16817.t1 VGND 0.08597f
C233 a_9573_16817.n1 VGND 0.215848f
C234 a_9573_16817.n2 VGND 2.65072f
C235 a_9573_16817.t3 VGND 0.08597f
C236 a_9573_16817.t6 VGND 0.08597f
C237 a_9573_16817.n3 VGND 0.215848f
C238 a_9573_16817.n4 VGND 2.27334f
C239 a_9573_16817.t10 VGND 0.047438f
C240 a_9573_16817.t7 VGND 0.046472f
C241 a_9573_16817.n5 VGND 0.362088f
C242 a_9573_16817.t9 VGND 0.046472f
C243 a_9573_16817.n6 VGND 0.193312f
C244 a_9573_16817.t8 VGND 0.047098f
C245 a_9573_16817.n7 VGND 0.194692f
C246 a_9573_16817.t11 VGND 0.047098f
C247 a_9573_16817.n8 VGND 0.89305f
C248 a_9573_16817.n9 VGND 2.97974f
C249 a_9573_16817.t0 VGND 1.33115f
C250 a_13880_11590.n0 VGND 0.019256f
C251 a_13880_11590.t0 VGND 0.034183f
C252 a_13880_11590.n1 VGND 0.021429f
C253 a_13880_11590.n2 VGND 0.554666f
C254 a_13880_11590.n3 VGND 0.186578f
C255 a_13880_11590.t4 VGND 0.027505f
C256 a_13880_11590.t10 VGND 0.021667f
C257 a_13880_11590.t22 VGND 0.021667f
C258 a_13880_11590.t19 VGND 0.034973f
C259 a_13880_11590.n4 VGND 0.039055f
C260 a_13880_11590.n5 VGND 0.02668f
C261 a_13880_11590.n6 VGND 0.043175f
C262 a_13880_11590.t5 VGND 0.018056f
C263 a_13880_11590.t11 VGND 0.018056f
C264 a_13880_11590.n7 VGND 0.036969f
C265 a_13880_11590.n8 VGND 0.191386f
C266 a_13880_11590.t12 VGND 0.027505f
C267 a_13880_11590.t6 VGND 0.021667f
C268 a_13880_11590.t18 VGND 0.021667f
C269 a_13880_11590.t20 VGND 0.034973f
C270 a_13880_11590.n9 VGND 0.039055f
C271 a_13880_11590.n10 VGND 0.02668f
C272 a_13880_11590.n11 VGND 0.043175f
C273 a_13880_11590.t13 VGND 0.018056f
C274 a_13880_11590.t7 VGND 0.018056f
C275 a_13880_11590.n12 VGND 0.036969f
C276 a_13880_11590.n13 VGND 0.191386f
C277 a_13880_11590.n14 VGND 0.26218f
C278 a_13880_11590.t14 VGND 0.027505f
C279 a_13880_11590.t8 VGND 0.021667f
C280 a_13880_11590.t17 VGND 0.021667f
C281 a_13880_11590.t21 VGND 0.034973f
C282 a_13880_11590.n15 VGND 0.039055f
C283 a_13880_11590.n16 VGND 0.02668f
C284 a_13880_11590.n17 VGND 0.043175f
C285 a_13880_11590.n18 VGND 0.239421f
C286 a_13880_11590.t9 VGND 0.018056f
C287 a_13880_11590.n19 VGND 0.036969f
C288 a_13880_11590.t15 VGND 0.018056f
C289 PFET_GATE.t17 VGND 0.026779f
C290 PFET_GATE.t27 VGND 0.026747f
C291 PFET_GATE.n0 VGND 0.139892f
C292 PFET_GATE.t21 VGND 0.026747f
C293 PFET_GATE.n1 VGND 0.073346f
C294 PFET_GATE.t12 VGND 0.026747f
C295 PFET_GATE.n2 VGND 0.073346f
C296 PFET_GATE.t23 VGND 0.026747f
C297 PFET_GATE.n3 VGND 0.073346f
C298 PFET_GATE.t15 VGND 0.026747f
C299 PFET_GATE.n4 VGND 0.073346f
C300 PFET_GATE.t26 VGND 0.026747f
C301 PFET_GATE.n5 VGND 0.073346f
C302 PFET_GATE.t28 VGND 0.026747f
C303 PFET_GATE.n6 VGND 0.073346f
C304 PFET_GATE.t19 VGND 0.026747f
C305 PFET_GATE.n7 VGND 0.073346f
C306 PFET_GATE.t10 VGND 0.026747f
C307 PFET_GATE.n8 VGND 0.181639f
C308 PFET_GATE.t14 VGND 0.026747f
C309 PFET_GATE.n9 VGND 0.181639f
C310 PFET_GATE.t25 VGND 0.026747f
C311 PFET_GATE.n10 VGND 0.073346f
C312 PFET_GATE.t20 VGND 0.026747f
C313 PFET_GATE.n11 VGND 0.073346f
C314 PFET_GATE.t11 VGND 0.026747f
C315 PFET_GATE.n12 VGND 0.073346f
C316 PFET_GATE.t22 VGND 0.026747f
C317 PFET_GATE.n13 VGND 0.073346f
C318 PFET_GATE.t13 VGND 0.026747f
C319 PFET_GATE.n14 VGND 0.073346f
C320 PFET_GATE.t24 VGND 0.026747f
C321 PFET_GATE.n15 VGND 0.073346f
C322 PFET_GATE.t16 VGND 0.026747f
C323 PFET_GATE.n16 VGND 0.073346f
C324 PFET_GATE.t18 VGND 0.026747f
C325 PFET_GATE.n17 VGND 0.073346f
C326 PFET_GATE.t29 VGND 0.026747f
C327 PFET_GATE.n18 VGND 0.829525f
C328 PFET_GATE.t7 VGND 0.234008f
C329 PFET_GATE.t9 VGND 0.01547f
C330 PFET_GATE.t5 VGND 0.01547f
C331 PFET_GATE.n19 VGND 0.033417f
C332 PFET_GATE.n20 VGND 0.763672f
C333 PFET_GATE.t1 VGND 0.01547f
C334 PFET_GATE.t3 VGND 0.01547f
C335 PFET_GATE.n21 VGND 0.033417f
C336 PFET_GATE.n22 VGND 0.337871f
C337 PFET_GATE.t6 VGND 0.01547f
C338 PFET_GATE.t2 VGND 0.01547f
C339 PFET_GATE.n23 VGND 0.033417f
C340 PFET_GATE.n24 VGND 0.330909f
C341 PFET_GATE.t4 VGND 0.01547f
C342 PFET_GATE.t8 VGND 0.01547f
C343 PFET_GATE.n25 VGND 0.033417f
C344 PFET_GATE.n26 VGND 0.76477f
C345 PFET_GATE.n27 VGND 2.03706f
C346 PFET_GATE.t0 VGND 0.906421f
C347 a_19440_11540.t7 VGND 0.032027f
C348 a_19440_11540.n0 VGND 0.178495f
C349 a_19440_11540.t0 VGND 0.021157f
C350 a_19440_11540.t12 VGND 0.021157f
C351 a_19440_11540.n1 VGND 0.0506f
C352 a_19440_11540.t9 VGND 0.021157f
C353 a_19440_11540.t5 VGND 0.021157f
C354 a_19440_11540.n2 VGND 0.0506f
C355 a_19440_11540.t6 VGND 0.085694f
C356 a_19440_11540.t4 VGND 0.032027f
C357 a_19440_11540.n3 VGND 0.150205f
C358 a_19440_11540.n4 VGND 0.14861f
C359 a_19440_11540.n5 VGND 0.149118f
C360 a_19440_11540.t2 VGND 0.052891f
C361 a_19440_11540.t10 VGND 0.052891f
C362 a_19440_11540.n6 VGND 0.109442f
C363 a_19440_11540.t3 VGND 0.052891f
C364 a_19440_11540.t11 VGND 0.052891f
C365 a_19440_11540.n7 VGND 0.158354f
C366 a_19440_11540.n8 VGND 1.17815f
C367 a_19440_11540.n9 VGND 0.051715f
C368 a_19440_11540.n10 VGND 0.147792f
C369 a_19440_11540.t1 VGND 0.021157f
C370 a_19440_11540.n11 VGND 0.050792f
C371 a_19440_11540.t8 VGND 0.109026f
C372 a_17290_6090.t0 VGND 0.023659f
C373 a_17290_6090.t2 VGND 2.0362f
C374 a_17290_6090.n0 VGND 0.026464f
C375 a_17290_6090.n1 VGND 0.060553f
C376 a_17290_6090.t1 VGND 0.044187f
C377 a_17450_6090.t10 VGND 3.04931f
C378 a_17450_6090.t12 VGND 3.0506f
C379 a_17450_6090.n2 VGND 0.038153f
C380 a_17450_6090.n3 VGND 0.034141f
C381 a_17450_6090.n4 VGND 0.019754f
C382 a_17450_6090.t13 VGND 0.040996f
C383 a_17450_6090.t11 VGND 0.040996f
C384 a_17450_6090.t14 VGND 0.017908f
C385 a_17450_6090.n5 VGND 0.021587f
C386 a_17450_6090.n6 VGND 0.021587f
C387 a_17450_6090.t15 VGND 0.017908f
C388 a_17450_6090.n7 VGND 0.019754f
C389 a_17450_6090.t0 VGND 0.038298f
C390 a_17450_6090.t9 VGND 0.012094f
C391 a_17450_6090.n9 VGND 0.059495f
C392 a_17450_6090.n10 VGND 0.724568f
C393 a_17450_6090.n11 VGND 0.343525f
C394 a_17450_6090.n12 VGND 0.034843f
C395 a_17450_6090.n13 VGND 0.012508f
C396 a_17450_6090.n14 VGND 0.048726f
C397 a_11880_10030.t9 VGND 0.13799f
C398 a_11880_10030.t30 VGND 0.138771f
C399 a_11880_10030.n0 VGND 0.061848f
C400 a_11880_10030.t32 VGND 0.139054f
C401 a_11880_10030.t33 VGND 0.139653f
C402 a_11880_10030.n1 VGND 0.175709f
C403 a_11880_10030.t22 VGND 0.139653f
C404 a_11880_10030.n2 VGND 0.09625f
C405 a_11880_10030.t49 VGND 0.139653f
C406 a_11880_10030.n3 VGND 0.09625f
C407 a_11880_10030.t40 VGND 0.139653f
C408 a_11880_10030.n4 VGND 0.09625f
C409 a_11880_10030.t29 VGND 0.139653f
C410 a_11880_10030.n5 VGND 0.09625f
C411 a_11880_10030.n6 VGND 0.02722f
C412 a_11880_10030.n7 VGND 0.018146f
C413 a_11880_10030.t24 VGND 0.138651f
C414 a_11880_10030.t31 VGND 0.139653f
C415 a_11880_10030.n8 VGND 0.175357f
C416 a_11880_10030.t43 VGND 0.139653f
C417 a_11880_10030.n9 VGND 0.09625f
C418 a_11880_10030.t18 VGND 0.139653f
C419 a_11880_10030.n10 VGND 0.09625f
C420 a_11880_10030.t27 VGND 0.139653f
C421 a_11880_10030.n11 VGND 0.09625f
C422 a_11880_10030.t26 VGND 0.139653f
C423 a_11880_10030.n12 VGND 0.09625f
C424 a_11880_10030.t37 VGND 0.139653f
C425 a_11880_10030.n13 VGND 0.09625f
C426 a_11880_10030.t45 VGND 0.138579f
C427 a_11880_10030.n14 VGND 0.091275f
C428 a_11880_10030.n15 VGND 0.02722f
C429 a_11880_10030.t19 VGND 0.137776f
C430 a_11880_10030.n16 VGND 0.056794f
C431 a_11880_10030.n17 VGND 0.096781f
C432 a_11880_10030.n18 VGND 0.377485f
C433 a_11880_10030.t7 VGND 0.010081f
C434 a_11880_10030.t11 VGND 0.010081f
C435 a_11880_10030.n19 VGND 0.021777f
C436 a_11880_10030.n20 VGND 0.20524f
C437 a_11880_10030.t3 VGND 0.010081f
C438 a_11880_10030.t4 VGND 0.010081f
C439 a_11880_10030.n21 VGND 0.021777f
C440 a_11880_10030.n22 VGND 0.220176f
C441 a_11880_10030.t8 VGND 0.010081f
C442 a_11880_10030.t6 VGND 0.010081f
C443 a_11880_10030.n23 VGND 0.021777f
C444 a_11880_10030.n24 VGND 0.214127f
C445 a_11880_10030.t10 VGND 0.010081f
C446 a_11880_10030.t5 VGND 0.010081f
C447 a_11880_10030.n25 VGND 0.020642f
C448 a_11880_10030.t1 VGND 0.010081f
C449 a_11880_10030.t13 VGND 0.010081f
C450 a_11880_10030.n26 VGND 0.023461f
C451 a_11880_10030.t12 VGND 0.010081f
C452 a_11880_10030.t2 VGND 0.010081f
C453 a_11880_10030.n27 VGND 0.020642f
C454 a_11880_10030.n28 VGND 0.276484f
C455 a_11880_10030.n29 VGND 0.170904f
C456 a_11880_10030.n30 VGND 0.676976f
C457 a_11880_10030.t14 VGND 0.403254f
C458 a_11880_10030.t21 VGND 0.409946f
C459 a_11880_10030.t17 VGND 0.403254f
C460 a_11880_10030.n31 VGND 0.268025f
C461 a_11880_10030.t47 VGND 0.403254f
C462 a_11880_10030.n32 VGND 0.176424f
C463 a_11880_10030.t20 VGND 0.403254f
C464 a_11880_10030.n33 VGND 0.176424f
C465 a_11880_10030.t16 VGND 0.403254f
C466 a_11880_10030.n34 VGND 0.176424f
C467 a_11880_10030.t25 VGND 0.403254f
C468 a_11880_10030.n35 VGND 0.176424f
C469 a_11880_10030.t35 VGND 0.403254f
C470 a_11880_10030.n36 VGND 0.176424f
C471 a_11880_10030.t44 VGND 0.403254f
C472 a_11880_10030.n37 VGND 0.176424f
C473 a_11880_10030.t39 VGND 0.403254f
C474 a_11880_10030.n38 VGND 0.176424f
C475 a_11880_10030.n39 VGND 0.176424f
C476 a_11880_10030.t38 VGND 0.403254f
C477 a_11880_10030.n40 VGND 0.176424f
C478 a_11880_10030.t28 VGND 0.403254f
C479 a_11880_10030.n41 VGND 0.176424f
C480 a_11880_10030.t34 VGND 0.403254f
C481 a_11880_10030.n42 VGND 0.176424f
C482 a_11880_10030.t23 VGND 0.403254f
C483 a_11880_10030.n43 VGND 0.176424f
C484 a_11880_10030.t15 VGND 0.403254f
C485 a_11880_10030.n44 VGND 0.176424f
C486 a_11880_10030.t41 VGND 0.403254f
C487 a_11880_10030.n45 VGND 0.176424f
C488 a_11880_10030.t46 VGND 0.403254f
C489 a_11880_10030.n46 VGND 0.176424f
C490 a_11880_10030.t36 VGND 0.403254f
C491 a_11880_10030.n47 VGND 0.176424f
C492 a_11880_10030.t42 VGND 0.403254f
C493 a_11880_10030.n48 VGND 0.175163f
C494 a_11880_10030.t48 VGND 0.403254f
C495 a_11880_10030.n49 VGND 0.371024f
C496 a_11880_10030.n50 VGND 1.17936f
C497 a_11880_10030.t0 VGND 0.155821f
C498 VDPWR.n1 VGND 0.044215f
C499 VDPWR.t44 VGND 0.027757f
C500 VDPWR.n3 VGND 0.033774f
C501 VDPWR.t194 VGND 0.022136f
C502 VDPWR.n5 VGND 0.033774f
C503 VDPWR.t380 VGND 0.026703f
C504 VDPWR.t22 VGND 0.025298f
C505 VDPWR.t75 VGND 0.025298f
C506 VDPWR.t371 VGND 0.022136f
C507 VDPWR.n8 VGND 0.060566f
C508 VDPWR.n10 VGND 0.040734f
C509 VDPWR.n11 VGND 0.033894f
C510 VDPWR.n13 VGND 0.021251f
C511 VDPWR.t61 VGND 0.04392f
C512 VDPWR.t73 VGND 0.042163f
C513 VDPWR.t220 VGND 0.025298f
C514 VDPWR.t410 VGND 0.025298f
C515 VDPWR.t4 VGND 0.022136f
C516 VDPWR.t246 VGND 0.025298f
C517 VDPWR.t118 VGND 0.025298f
C518 VDPWR.t133 VGND 0.042163f
C519 VDPWR.t283 VGND 0.04392f
C520 VDPWR.n14 VGND 0.021251f
C521 VDPWR.n16 VGND 0.033894f
C522 VDPWR.n18 VGND 0.040734f
C523 VDPWR.n20 VGND 0.033774f
C524 VDPWR.n22 VGND 0.040734f
C525 VDPWR.n23 VGND 0.033894f
C526 VDPWR.n25 VGND 0.021251f
C527 VDPWR.t395 VGND 0.04392f
C528 VDPWR.t208 VGND 0.042163f
C529 VDPWR.t102 VGND 0.025298f
C530 VDPWR.t167 VGND 0.025298f
C531 VDPWR.t30 VGND 0.022136f
C532 VDPWR.t40 VGND 0.031622f
C533 VDPWR.t14 VGND 0.031622f
C534 VDPWR.t58 VGND 0.025298f
C535 VDPWR.t48 VGND 0.025298f
C536 VDPWR.t104 VGND 0.040757f
C537 VDPWR.t227 VGND 0.040757f
C538 VDPWR.t397 VGND 0.03092f
C539 VDPWR.t424 VGND 0.03092f
C540 VDPWR.t206 VGND 0.043568f
C541 VDPWR.t188 VGND 0.045325f
C542 VDPWR.n26 VGND 0.021251f
C543 VDPWR.n28 VGND 0.034429f
C544 VDPWR.n30 VGND 0.043412f
C545 VDPWR.n32 VGND 0.039396f
C546 VDPWR.n33 VGND 0.034015f
C547 VDPWR.n34 VGND 0.028125f
C548 VDPWR.n36 VGND 0.033507f
C549 VDPWR.n38 VGND 0.038325f
C550 VDPWR.n40 VGND 0.04823f
C551 VDPWR.n42 VGND 0.04978f
C552 VDPWR.n43 VGND 0.039248f
C553 VDPWR.n45 VGND 0.026873f
C554 VDPWR.t100 VGND 0.053055f
C555 VDPWR.t34 VGND 0.051298f
C556 VDPWR.t32 VGND 0.01546f
C557 VDPWR.t250 VGND 0.03092f
C558 VDPWR.t404 VGND 0.03092f
C559 VDPWR.t81 VGND 0.047082f
C560 VDPWR.t244 VGND 0.047082f
C561 VDPWR.t402 VGND 0.027757f
C562 VDPWR.t83 VGND 0.060785f
C563 VDPWR.n46 VGND 0.026873f
C564 VDPWR.n48 VGND 0.647049f
C565 VDPWR.n49 VGND 0.015387f
C566 VDPWR.n50 VGND 0.068671f
C567 VDPWR.n51 VGND 0.015004f
C568 VDPWR.n52 VGND 0.012047f
C569 VDPWR.n53 VGND 0.020078f
C570 VDPWR.t357 VGND 0.083456f
C571 VDPWR.t356 VGND 0.031478f
C572 VDPWR.t341 VGND 0.031478f
C573 VDPWR.n57 VGND 0.014181f
C574 VDPWR.n58 VGND 0.035365f
C575 VDPWR.n59 VGND 0.020078f
C576 VDPWR.n60 VGND 0.018739f
C577 VDPWR.t306 VGND 0.03364f
C578 VDPWR.n62 VGND 0.021281f
C579 VDPWR.n64 VGND 0.010842f
C580 VDPWR.n66 VGND 0.012047f
C581 VDPWR.n70 VGND 0.015004f
C582 VDPWR.n71 VGND 0.012047f
C583 VDPWR.t231 VGND 0.085397f
C584 VDPWR.t190 VGND 0.085397f
C585 VDPWR.t238 VGND 0.085397f
C586 VDPWR.t225 VGND 0.085397f
C587 VDPWR.t307 VGND 0.083456f
C588 VDPWR.n74 VGND 0.075693f
C589 VDPWR.n76 VGND 0.010922f
C590 VDPWR.n77 VGND 0.020078f
C591 VDPWR.t308 VGND 0.013385f
C592 VDPWR.n78 VGND 0.015387f
C593 VDPWR.n79 VGND 0.076326f
C594 VDPWR.n80 VGND 0.015387f
C595 VDPWR.n81 VGND 0.074561f
C596 VDPWR.n82 VGND 0.015387f
C597 VDPWR.n83 VGND 0.071348f
C598 VDPWR.n86 VGND 0.018739f
C599 VDPWR.n87 VGND 0.018739f
C600 VDPWR.n88 VGND 0.018182f
C601 VDPWR.n89 VGND 0.028674f
C602 VDPWR.n90 VGND 0.017638f
C603 VDPWR.n91 VGND 0.015387f
C604 VDPWR.n92 VGND 0.074561f
C605 VDPWR.n93 VGND 0.071348f
C606 VDPWR.n94 VGND 0.015387f
C607 VDPWR.t343 VGND 0.013385f
C608 VDPWR.n95 VGND 0.020078f
C609 VDPWR.n97 VGND 0.024405f
C610 VDPWR.n99 VGND 0.081515f
C611 VDPWR.t342 VGND 0.083456f
C612 VDPWR.t18 VGND 0.085397f
C613 VDPWR.t234 VGND 0.085397f
C614 VDPWR.t236 VGND 0.085397f
C615 VDPWR.t153 VGND 0.085397f
C616 VDPWR.t303 VGND 0.083456f
C617 VDPWR.n102 VGND 0.012047f
C618 VDPWR.n104 VGND 0.012238f
C619 VDPWR.n106 VGND 0.075693f
C620 VDPWR.n108 VGND 0.012158f
C621 VDPWR.t302 VGND 0.03364f
C622 VDPWR.n110 VGND 0.020717f
C623 VDPWR.n111 VGND 0.025649f
C624 VDPWR.n112 VGND 0.028003f
C625 VDPWR.n118 VGND 0.096125f
C626 VDPWR.n128 VGND 0.021486f
C627 VDPWR.n129 VGND 0.028213f
C628 VDPWR.t383 VGND 0.01409f
C629 VDPWR.n140 VGND 0.096125f
C630 VDPWR.n150 VGND 0.021486f
C631 VDPWR.n151 VGND 0.028213f
C632 VDPWR.t55 VGND 0.01409f
C633 VDPWR.n157 VGND 0.010563f
C634 VDPWR.n159 VGND 0.069414f
C635 VDPWR.n160 VGND 0.035928f
C636 VDPWR.n161 VGND 0.069414f
C637 VDPWR.n162 VGND 0.144328f
C638 VDPWR.n163 VGND 0.044193f
C639 VDPWR.n165 VGND 0.015625f
C640 VDPWR.n171 VGND 0.096125f
C641 VDPWR.n181 VGND 0.021486f
C642 VDPWR.n182 VGND 0.028213f
C643 VDPWR.t413 VGND 0.01409f
C644 VDPWR.n188 VGND 0.010563f
C645 VDPWR.n189 VGND 0.041816f
C646 VDPWR.t121 VGND 0.014426f
C647 VDPWR.n190 VGND 0.051402f
C648 VDPWR.n192 VGND 0.011251f
C649 VDPWR.n193 VGND 0.02327f
C650 VDPWR.n194 VGND 0.284119f
C651 VDPWR.t120 VGND 0.556208f
C652 VDPWR.t412 VGND 0.488772f
C653 VDPWR.t265 VGND 0.101486f
C654 VDPWR.t181 VGND 0.108202f
C655 VDPWR.n195 VGND 0.286548f
C656 VDPWR.t54 VGND 0.279832f
C657 VDPWR.t269 VGND 0.101486f
C658 VDPWR.t224 VGND 0.287294f
C659 VDPWR.t382 VGND 0.387287f
C660 VDPWR.t267 VGND 0.101486f
C661 VDPWR.t166 VGND 0.210793f
C662 VDPWR.n196 VGND 0.211298f
C663 VDPWR.n197 VGND 0.049205f
C664 VDPWR.n198 VGND 0.024439f
C665 VDPWR.n199 VGND 0.010563f
C666 VDPWR.n200 VGND 0.109796f
C667 VDPWR.n201 VGND 2.28944f
C668 VDPWR.n202 VGND 0.02698f
C669 VDPWR.n203 VGND 0.01332f
C670 VDPWR.t158 VGND 0.10166f
C671 VDPWR.n211 VGND 0.014724f
C672 VDPWR.n214 VGND 0.014724f
C673 VDPWR.n215 VGND 0.017622f
C674 VDPWR.n219 VGND 0.014724f
C675 VDPWR.t159 VGND 0.014123f
C676 VDPWR.n222 VGND 0.014677f
C677 VDPWR.n224 VGND 0.0208f
C678 VDPWR.n225 VGND 0.01332f
C679 VDPWR.n228 VGND 0.080913f
C680 VDPWR.t177 VGND 0.019887f
C681 VDPWR.n232 VGND 0.025087f
C682 VDPWR.n234 VGND 0.0235f
C683 VDPWR.t420 VGND 0.056016f
C684 VDPWR.t98 VGND 0.161825f
C685 VDPWR.n245 VGND 0.020078f
C686 VDPWR.n246 VGND 0.020078f
C687 VDPWR.n248 VGND 0.012158f
C688 VDPWR.n249 VGND 0.012047f
C689 VDPWR.n252 VGND 0.012047f
C690 VDPWR.n253 VGND 0.014291f
C691 VDPWR.n254 VGND 0.052515f
C692 VDPWR.n255 VGND 0.020078f
C693 VDPWR.n256 VGND 0.012047f
C694 VDPWR.t186 VGND 0.188796f
C695 VDPWR.n262 VGND 0.020078f
C696 VDPWR.n263 VGND 0.020078f
C697 VDPWR.n265 VGND 0.012158f
C698 VDPWR.n266 VGND 0.012047f
C699 VDPWR.n269 VGND 0.012047f
C700 VDPWR.n270 VGND 0.014291f
C701 VDPWR.n271 VGND 0.020078f
C702 VDPWR.n272 VGND 0.012047f
C703 VDPWR.t408 VGND 0.197095f
C704 VDPWR.n277 VGND 0.012047f
C705 VDPWR.n278 VGND 0.010842f
C706 VDPWR.t6 VGND 0.213693f
C707 VDPWR.n280 VGND 0.161825f
C708 VDPWR.n282 VGND 0.014876f
C709 VDPWR.n283 VGND 0.054803f
C710 VDPWR.n285 VGND 0.014291f
C711 VDPWR.n287 VGND 0.012047f
C712 VDPWR.n289 VGND 0.012047f
C713 VDPWR.n290 VGND 0.012158f
C714 VDPWR.n292 VGND 0.161825f
C715 VDPWR.t229 VGND 0.161825f
C716 VDPWR.n293 VGND 0.012158f
C717 VDPWR.n295 VGND 0.012047f
C718 VDPWR.n298 VGND 0.161825f
C719 VDPWR.n300 VGND 0.01576f
C720 VDPWR.n301 VGND 0.025042f
C721 VDPWR.n302 VGND 0.025106f
C722 VDPWR.n304 VGND 0.014291f
C723 VDPWR.n306 VGND 0.012047f
C724 VDPWR.n308 VGND 0.012047f
C725 VDPWR.n309 VGND 0.012158f
C726 VDPWR.n311 VGND 0.176348f
C727 VDPWR.t108 VGND 0.056016f
C728 VDPWR.t421 VGND 0.014116f
C729 VDPWR.n315 VGND 0.013036f
C730 VDPWR.n317 VGND 0.114108f
C731 VDPWR.n319 VGND 0.01332f
C732 VDPWR.n324 VGND 0.013036f
C733 VDPWR.t109 VGND 0.014116f
C734 VDPWR.n326 VGND 0.01332f
C735 VDPWR.n328 VGND 0.080913f
C736 VDPWR.t160 VGND 0.056016f
C737 VDPWR.t414 VGND 0.056016f
C738 VDPWR.t161 VGND 0.014116f
C739 VDPWR.n332 VGND 0.013036f
C740 VDPWR.n334 VGND 0.080913f
C741 VDPWR.n336 VGND 0.01332f
C742 VDPWR.t415 VGND 0.014116f
C743 VDPWR.n340 VGND 0.013036f
C744 VDPWR.n345 VGND 0.01332f
C745 VDPWR.n347 VGND 0.017342f
C746 VDPWR.n352 VGND 0.013177f
C747 VDPWR.t39 VGND 0.014116f
C748 VDPWR.n356 VGND 0.013036f
C749 VDPWR.n358 VGND 0.080913f
C750 VDPWR.t176 VGND 0.051867f
C751 VDPWR.t2 VGND 0.049793f
C752 VDPWR.t38 VGND 0.056016f
C753 VDPWR.n364 VGND 0.013036f
C754 VDPWR.t3 VGND 0.014046f
C755 VDPWR.n366 VGND 0.014529f
C756 VDPWR.n368 VGND 0.109958f
C757 VDPWR.t117 VGND 0.215767f
C758 VDPWR.t132 VGND 0.215767f
C759 VDPWR.t106 VGND 0.10166f
C760 VDPWR.t107 VGND 0.014116f
C761 VDPWR.n370 VGND 0.013036f
C762 VDPWR.t233 VGND 0.014116f
C763 VDPWR.n380 VGND 0.013036f
C764 VDPWR.n382 VGND 0.114108f
C765 VDPWR.n384 VGND 0.01332f
C766 VDPWR.n386 VGND 0.029389f
C767 VDPWR.n387 VGND 0.02698f
C768 VDPWR.n390 VGND 0.014677f
C769 VDPWR.n393 VGND 0.014724f
C770 VDPWR.t172 VGND 0.014123f
C771 VDPWR.n396 VGND 0.017622f
C772 VDPWR.n398 VGND 0.112033f
C773 VDPWR.t42 VGND 0.10166f
C774 VDPWR.t171 VGND 0.215767f
C775 VDPWR.t11 VGND 0.215767f
C776 VDPWR.t71 VGND 0.10166f
C777 VDPWR.t72 VGND 0.014116f
C778 VDPWR.n400 VGND 0.013036f
C779 VDPWR.t178 VGND 0.014116f
C780 VDPWR.n410 VGND 0.013036f
C781 VDPWR.n412 VGND 0.122406f
C782 VDPWR.n414 VGND 0.01332f
C783 VDPWR.n416 VGND 0.71534f
C784 VDPWR.t399 VGND 0.149645f
C785 VDPWR.t173 VGND 0.157676f
C786 VDPWR.t137 VGND 0.157676f
C787 VDPWR.t384 VGND 0.157676f
C788 VDPWR.t112 VGND 0.157676f
C789 VDPWR.t377 VGND 0.157676f
C790 VDPWR.t368 VGND 0.157676f
C791 VDPWR.t56 VGND 0.157676f
C792 VDPWR.t196 VGND 0.150187f
C793 VDPWR.t122 VGND 0.072346f
C794 VDPWR.n417 VGND 0.093316f
C795 VDPWR.t376 VGND 0.164037f
C796 VDPWR.t123 VGND 0.150818f
C797 VDPWR.t142 VGND 0.157676f
C798 VDPWR.t57 VGND 0.157676f
C799 VDPWR.t388 VGND 0.157676f
C800 VDPWR.t46 VGND 0.157676f
C801 VDPWR.t422 VGND 0.157676f
C802 VDPWR.t385 VGND 0.157676f
C803 VDPWR.t47 VGND 0.157676f
C804 VDPWR.t423 VGND 0.293276f
C805 VDPWR.t426 VGND 0.316242f
C806 VDPWR.t427 VGND 0.316242f
C807 VDPWR.t431 VGND 0.300446f
C808 VDPWR.n418 VGND 0.5815f
C809 VDPWR.n419 VGND 0.307031f
C810 VDPWR.t433 VGND 0.296783f
C811 VDPWR.n420 VGND 0.533168f
C812 VDPWR.n421 VGND 0.482849f
C813 VDPWR.n422 VGND 0.019804f
C814 VDPWR.n423 VGND 0.079379f
C815 VDPWR.n424 VGND 0.010093f
C816 VDPWR.t130 VGND 0.07233f
C817 VDPWR.n431 VGND 0.083509f
C818 VDPWR.n435 VGND 0.025097f
C819 VDPWR.n436 VGND 0.012047f
C820 VDPWR.t361 VGND 0.129316f
C821 VDPWR.t16 VGND 0.113974f
C822 VDPWR.t7 VGND 0.113974f
C823 VDPWR.t12 VGND 0.113974f
C824 VDPWR.t113 VGND 0.113974f
C825 VDPWR.t351 VGND 0.225286f
C826 VDPWR.t352 VGND 0.015347f
C827 VDPWR.n441 VGND 0.091982f
C828 VDPWR.n443 VGND 0.014472f
C829 VDPWR.t363 VGND 0.011994f
C830 VDPWR.n445 VGND 0.025174f
C831 VDPWR.n447 VGND 0.014472f
C832 VDPWR.n448 VGND 0.020945f
C833 VDPWR.n449 VGND 0.019804f
C834 VDPWR.n450 VGND 0.084733f
C835 VDPWR.n451 VGND 0.019804f
C836 VDPWR.n452 VGND 0.084733f
C837 VDPWR.n453 VGND 0.017387f
C838 VDPWR.n454 VGND 0.065734f
C839 VDPWR.n455 VGND 0.01285f
C840 VDPWR.n456 VGND 0.010708f
C841 VDPWR.t346 VGND 0.016731f
C842 VDPWR.n457 VGND 0.019804f
C843 VDPWR.n458 VGND 0.077237f
C844 VDPWR.n459 VGND 0.047486f
C845 VDPWR.t344 VGND 0.033436f
C846 VDPWR.n460 VGND 0.024384f
C847 VDPWR.n462 VGND 0.012158f
C848 VDPWR.n464 VGND 0.012047f
C849 VDPWR.n467 VGND 0.012047f
C850 VDPWR.n468 VGND 0.015004f
C851 VDPWR.n470 VGND 0.010922f
C852 VDPWR.n472 VGND 0.070138f
C853 VDPWR.t313 VGND 0.07233f
C854 VDPWR.t242 VGND 0.07233f
C855 VDPWR.t36 VGND 0.056987f
C856 VDPWR.t192 VGND 0.087672f
C857 VDPWR.t378 VGND 0.056987f
C858 VDPWR.t28 VGND 0.067946f
C859 VDPWR.t369 VGND 0.076713f
C860 VDPWR.t135 VGND 0.056987f
C861 VDPWR.t348 VGND 0.087672f
C862 VDPWR.t345 VGND 0.07233f
C863 VDPWR.n473 VGND 0.094481f
C864 VDPWR.t349 VGND 0.015348f
C865 VDPWR.n474 VGND 0.039535f
C866 VDPWR.n476 VGND 0.023505f
C867 VDPWR.n477 VGND 0.028839f
C868 VDPWR.n478 VGND 0.023505f
C869 VDPWR.t315 VGND 0.011997f
C870 VDPWR.n480 VGND 0.034773f
C871 VDPWR.n481 VGND 0.094473f
C872 VDPWR.t88 VGND 0.118357f
C873 VDPWR.t67 VGND 0.111782f
C874 VDPWR.t373 VGND 0.081097f
C875 VDPWR.t85 VGND 0.063562f
C876 VDPWR.t86 VGND 0.056987f
C877 VDPWR.t60 VGND 0.087672f
C878 VDPWR.t169 VGND 0.056987f
C879 VDPWR.t394 VGND 0.076713f
C880 VDPWR.t157 VGND 0.067946f
C881 VDPWR.t317 VGND 0.056987f
C882 VDPWR.t389 VGND 0.087672f
C883 VDPWR.n485 VGND 0.012047f
C884 VDPWR.n486 VGND 0.015004f
C885 VDPWR.n487 VGND 0.012047f
C886 VDPWR.n488 VGND 0.012047f
C887 VDPWR.n490 VGND 0.025097f
C888 VDPWR.n491 VGND 0.012238f
C889 VDPWR.n493 VGND 0.18192f
C890 VDPWR.n495 VGND 0.013552f
C891 VDPWR.t316 VGND 0.033151f
C892 VDPWR.n496 VGND 0.016144f
C893 VDPWR.n497 VGND 0.071797f
C894 VDPWR.n498 VGND 0.160992f
C895 VDPWR.n500 VGND 0.071565f
C896 VDPWR.n501 VGND 0.010409f
C897 VDPWR.n502 VGND 0.010329f
C898 VDPWR.n504 VGND 0.071565f
C899 VDPWR.n506 VGND 0.071565f
C900 VDPWR.n508 VGND 0.071565f
C901 VDPWR.n510 VGND 0.071565f
C902 VDPWR.n512 VGND 0.071565f
C903 VDPWR.n514 VGND 0.071565f
C904 VDPWR.n516 VGND 0.071565f
C905 VDPWR.n518 VGND 0.071565f
C906 VDPWR.n520 VGND 0.071565f
C907 VDPWR.n521 VGND 0.010409f
C908 VDPWR.n522 VGND 0.010329f
C909 VDPWR.n524 VGND 0.071565f
C910 VDPWR.n526 VGND 0.071565f
C911 VDPWR.n528 VGND 0.071565f
C912 VDPWR.n530 VGND 0.071565f
C913 VDPWR.n532 VGND 0.071565f
C914 VDPWR.n534 VGND 0.071565f
C915 VDPWR.n536 VGND 0.071565f
C916 VDPWR.n538 VGND 0.097517f
C917 VDPWR.n539 VGND 0.031296f
C918 VDPWR.n541 VGND 0.010409f
C919 VDPWR.n542 VGND 0.032999f
C920 VDPWR.t300 VGND 0.027782f
C921 VDPWR.t277 VGND 0.022487f
C922 VDPWR.t149 VGND 0.022487f
C923 VDPWR.t179 VGND 0.022487f
C924 VDPWR.t0 VGND 0.022487f
C925 VDPWR.t182 VGND 0.022487f
C926 VDPWR.t273 VGND 0.022487f
C927 VDPWR.t281 VGND 0.022487f
C928 VDPWR.t94 VGND 0.022487f
C929 VDPWR.t240 VGND 0.022487f
C930 VDPWR.t52 VGND 0.022487f
C931 VDPWR.t96 VGND 0.022487f
C932 VDPWR.t275 VGND 0.022487f
C933 VDPWR.t271 VGND 0.022487f
C934 VDPWR.t216 VGND 0.022487f
C935 VDPWR.t151 VGND 0.022487f
C936 VDPWR.t285 VGND 0.022487f
C937 VDPWR.t248 VGND 0.022487f
C938 VDPWR.t279 VGND 0.022487f
C939 VDPWR.t324 VGND 0.034169f
C940 VDPWR.n543 VGND 0.028485f
C941 VDPWR.n544 VGND 0.010329f
C942 VDPWR.n546 VGND 0.022102f
C943 VDPWR.n547 VGND 0.072751f
C944 VDPWR.n548 VGND 0.072751f
C945 VDPWR.n549 VGND 0.029472f
C946 VDPWR.n551 VGND 0.010409f
C947 VDPWR.n552 VGND 0.034644f
C948 VDPWR.t310 VGND 0.02801f
C949 VDPWR.t261 VGND 0.022487f
C950 VDPWR.t20 VGND 0.022487f
C951 VDPWR.t291 VGND 0.022487f
C952 VDPWR.t287 VGND 0.022487f
C953 VDPWR.t251 VGND 0.022487f
C954 VDPWR.t255 VGND 0.022487f
C955 VDPWR.t253 VGND 0.022487f
C956 VDPWR.t364 VGND 0.022487f
C957 VDPWR.t69 VGND 0.022487f
C958 VDPWR.t140 VGND 0.022487f
C959 VDPWR.t65 VGND 0.022487f
C960 VDPWR.t259 VGND 0.022487f
C961 VDPWR.t263 VGND 0.022487f
C962 VDPWR.t184 VGND 0.022487f
C963 VDPWR.t289 VGND 0.022487f
C964 VDPWR.t126 VGND 0.022487f
C965 VDPWR.t50 VGND 0.022487f
C966 VDPWR.t257 VGND 0.022487f
C967 VDPWR.t294 VGND 0.033648f
C968 VDPWR.n553 VGND 0.027132f
C969 VDPWR.n554 VGND 0.010329f
C970 VDPWR.n556 VGND 0.022102f
C971 VDPWR.n557 VGND 0.277043f
C972 VDPWR.n558 VGND 0.274632f
C973 VDPWR.t296 VGND 0.038295f
C974 VDPWR.n559 VGND 0.01468f
C975 VDPWR.n560 VGND 0.031248f
C976 VDPWR.n561 VGND 0.031248f
C977 VDPWR.n562 VGND 0.031248f
C978 VDPWR.n563 VGND 0.031248f
C979 VDPWR.n564 VGND 0.031248f
C980 VDPWR.n565 VGND 0.031248f
C981 VDPWR.n566 VGND 0.031248f
C982 VDPWR.n567 VGND 0.031248f
C983 VDPWR.n582 VGND 0.010697f
C984 VDPWR.n591 VGND 0.010098f
C985 VDPWR.n593 VGND 0.07509f
C986 VDPWR.t297 VGND 0.079641f
C987 VDPWR.t90 VGND 0.081917f
C988 VDPWR.t92 VGND 0.081917f
C989 VDPWR.t366 VGND 0.081917f
C990 VDPWR.t400 VGND 0.081917f
C991 VDPWR.t110 VGND 0.081917f
C992 VDPWR.t197 VGND 0.081917f
C993 VDPWR.t145 VGND 0.081917f
C994 VDPWR.t212 VGND 0.081917f
C995 VDPWR.t143 VGND 0.081917f
C996 VDPWR.t138 VGND 0.081917f
C997 VDPWR.t416 VGND 0.081917f
C998 VDPWR.t418 VGND 0.081917f
C999 VDPWR.t210 VGND 0.081917f
C1000 VDPWR.t174 VGND 0.081917f
C1001 VDPWR.t147 VGND 0.081917f
C1002 VDPWR.t386 VGND 0.081917f
C1003 VDPWR.t339 VGND 0.079641f
C1004 VDPWR.n608 VGND 0.011297f
C1005 VDPWR.n610 VGND 0.07509f
C1006 VDPWR.n612 VGND 0.010697f
C1007 VDPWR.t338 VGND 0.038295f
C1008 VDPWR.n613 VGND 0.015467f
C1009 VDPWR.n614 VGND 0.153046f
C1010 VDPWR.n615 VGND 0.107421f
C1011 VDPWR.n616 VGND 0.107421f
C1012 VDPWR.n617 VGND 0.107421f
C1013 VDPWR.n618 VGND 0.107421f
C1014 VDPWR.n619 VGND 0.107421f
C1015 VDPWR.n620 VGND 0.107421f
C1016 VDPWR.n621 VGND 0.107421f
C1017 VDPWR.n622 VGND 0.090582f
C1018 VDPWR.n623 VGND 0.089327f
C1019 VDPWR.n624 VGND 0.010409f
C1020 VDPWR.n625 VGND 0.010946f
C1021 VDPWR.n626 VGND 0.034067f
C1022 VDPWR.t355 VGND 0.010623f
C1023 VDPWR.n628 VGND 0.011025f
C1024 VDPWR.n629 VGND 0.033516f
C1025 VDPWR.t354 VGND 0.027264f
C1026 VDPWR.t218 VGND 0.020613f
C1027 VDPWR.t219 VGND 0.020613f
C1028 VDPWR.t333 VGND 0.032355f
C1029 VDPWR.n630 VGND 0.026551f
C1030 VDPWR.n631 VGND 0.010329f
C1031 VDPWR.n633 VGND 0.025662f
C1032 VDPWR.n634 VGND 0.297201f
C1033 VDPWR.n635 VGND 0.270196f
C1034 VDPWR.n637 VGND 0.031696f
C1035 VDPWR.n638 VGND 0.010488f
C1036 VDPWR.n639 VGND 0.010329f
C1037 VDPWR.n642 VGND 0.031696f
C1038 VDPWR.n644 VGND 0.031696f
C1039 VDPWR.n646 VGND 0.031696f
C1040 VDPWR.n648 VGND 0.031696f
C1041 VDPWR.n650 VGND 0.031696f
C1042 VDPWR.n651 VGND 0.010488f
C1043 VDPWR.n652 VGND 0.010329f
C1044 VDPWR.n655 VGND 0.031696f
C1045 VDPWR.n657 VGND 0.031696f
C1046 VDPWR.n659 VGND 0.031696f
C1047 VDPWR.n661 VGND 0.039157f
C1048 VDPWR.n662 VGND 0.013274f
C1049 VDPWR.n663 VGND 0.017628f
C1050 VDPWR.n664 VGND 0.010488f
C1051 VDPWR.n665 VGND 0.032478f
C1052 VDPWR.t336 VGND 0.026428f
C1053 VDPWR.t200 VGND 0.020613f
C1054 VDPWR.t222 VGND 0.020613f
C1055 VDPWR.t374 VGND 0.020613f
C1056 VDPWR.t26 VGND 0.020613f
C1057 VDPWR.t128 VGND 0.020613f
C1058 VDPWR.t155 VGND 0.020613f
C1059 VDPWR.t124 VGND 0.020613f
C1060 VDPWR.t24 VGND 0.020613f
C1061 VDPWR.t406 VGND 0.020613f
C1062 VDPWR.t390 VGND 0.020613f
C1063 VDPWR.t327 VGND 0.032355f
C1064 VDPWR.n666 VGND 0.026551f
C1065 VDPWR.n667 VGND 0.010329f
C1066 VDPWR.n668 VGND 0.017628f
C1067 VDPWR.n669 VGND 0.012704f
C1068 VDPWR.n670 VGND 0.021416f
C1069 VDPWR.n671 VGND 0.021416f
C1070 VDPWR.n672 VGND 0.012704f
C1071 VDPWR.n673 VGND 0.017628f
C1072 VDPWR.n674 VGND 0.010488f
C1073 VDPWR.n675 VGND 0.032478f
C1074 VDPWR.t330 VGND 0.026428f
C1075 VDPWR.t79 VGND 0.020613f
C1076 VDPWR.t204 VGND 0.020613f
C1077 VDPWR.t115 VGND 0.020613f
C1078 VDPWR.t392 VGND 0.020613f
C1079 VDPWR.t162 VGND 0.020613f
C1080 VDPWR.t9 VGND 0.020613f
C1081 VDPWR.t164 VGND 0.020613f
C1082 VDPWR.t63 VGND 0.020613f
C1083 VDPWR.t214 VGND 0.020613f
C1084 VDPWR.t77 VGND 0.020613f
C1085 VDPWR.t321 VGND 0.032355f
C1086 VDPWR.n676 VGND 0.026551f
C1087 VDPWR.n677 VGND 0.010329f
C1088 VDPWR.n678 VGND 0.017628f
C1089 VDPWR.n679 VGND 0.012704f
C1090 VDPWR.n680 VGND 0.117109f
C1091 VDPWR.n681 VGND 2.31842f
C1092 VDPWR.n682 VGND 12.2733f
C1093 VDPWR.n683 VGND 1.85173f
C1094 VDPWR.n684 VGND 1.9729f
C1095 a_8454_18026.t18 VGND 0.270217f
C1096 a_8454_18026.t2 VGND 0.284719f
C1097 a_8454_18026.t6 VGND 0.284719f
C1098 a_8454_18026.t20 VGND 0.284719f
C1099 a_8454_18026.t3 VGND 0.284719f
C1100 a_8454_18026.t16 VGND 0.284719f
C1101 a_8454_18026.t11 VGND 0.284719f
C1102 a_8454_18026.t8 VGND 0.284719f
C1103 a_8454_18026.t9 VGND 0.271196f
C1104 a_8454_18026.t5 VGND 0.130637f
C1105 a_8454_18026.n0 VGND 0.168502f
C1106 a_8454_18026.t17 VGND 0.296204f
C1107 a_8454_18026.t4 VGND 0.272335f
C1108 a_8454_18026.t1 VGND 0.284719f
C1109 a_8454_18026.t7 VGND 0.284719f
C1110 a_8454_18026.t10 VGND 0.284719f
C1111 a_8454_18026.t15 VGND 0.284719f
C1112 a_8454_18026.t13 VGND 0.284719f
C1113 a_8454_18026.t19 VGND 0.284719f
C1114 a_8454_18026.t14 VGND 0.284719f
C1115 a_8454_18026.t12 VGND 1.3341f
C1116 a_8454_18026.t0 VGND 0.470749f
C1117 a_10710_11860.n0 VGND 1.01403f
C1118 a_10710_11860.n1 VGND 0.777726f
C1119 a_10710_11860.n2 VGND 2.14452f
C1120 a_10710_11860.n3 VGND 0.460584f
C1121 a_10710_11860.n4 VGND 0.152132f
C1122 a_10710_11860.n5 VGND 0.249616f
C1123 a_10710_11860.t19 VGND 0.021328f
C1124 a_10710_11860.n6 VGND 0.019491f
C1125 a_10710_11860.t33 VGND 0.013761f
C1126 a_10710_11860.t23 VGND 0.013761f
C1127 a_10710_11860.n7 VGND 0.026658f
C1128 a_10710_11860.n8 VGND 0.019491f
C1129 a_10710_11860.t3 VGND 0.015654f
C1130 a_10710_11860.n9 VGND 0.011231f
C1131 a_10710_11860.n10 VGND 0.010836f
C1132 a_10710_11860.n11 VGND 0.289023f
C1133 a_10710_11860.t14 VGND 0.013761f
C1134 a_10710_11860.t27 VGND 0.013761f
C1135 a_10710_11860.n12 VGND 0.025567f
C1136 a_10710_11860.t20 VGND 0.021048f
C1137 a_10710_11860.t15 VGND 0.355532f
C1138 a_10710_11860.t22 VGND 0.361432f
C1139 a_10710_11860.t18 VGND 0.355532f
C1140 a_10710_11860.t12 VGND 0.355532f
C1141 a_10710_11860.t21 VGND 0.355532f
C1142 a_10710_11860.t17 VGND 0.355532f
C1143 a_10710_11860.t25 VGND 0.355532f
C1144 a_10710_11860.t29 VGND 0.355532f
C1145 a_10710_11860.t36 VGND 0.355532f
C1146 a_10710_11860.t32 VGND 0.355532f
C1147 a_10710_11860.t31 VGND 0.355532f
C1148 a_10710_11860.t26 VGND 0.355532f
C1149 a_10710_11860.t28 VGND 0.355532f
C1150 a_10710_11860.t24 VGND 0.355532f
C1151 a_10710_11860.t16 VGND 0.355532f
C1152 a_10710_11860.t34 VGND 0.355532f
C1153 a_10710_11860.t11 VGND 0.355532f
C1154 a_10710_11860.t30 VGND 0.355532f
C1155 a_10710_11860.t35 VGND 0.355532f
C1156 a_10710_11860.t13 VGND 0.355532f
C1157 a_10710_11860.n13 VGND 0.97888f
C1158 a_10710_11860.n14 VGND 0.019491f
C1159 I_IN.t5 VGND 0.010427f
C1160 I_IN.t1 VGND 0.010427f
C1161 I_IN.n0 VGND 0.022175f
C1162 I_IN.t6 VGND 0.010427f
C1163 I_IN.t11 VGND 0.010427f
C1164 I_IN.n1 VGND 0.022089f
C1165 I_IN.n2 VGND 0.491704f
C1166 I_IN.t8 VGND 0.010427f
C1167 I_IN.t17 VGND 0.010427f
C1168 I_IN.n3 VGND 0.022089f
C1169 I_IN.n4 VGND 0.267792f
C1170 I_IN.t9 VGND 0.010427f
C1171 I_IN.t0 VGND 0.010427f
C1172 I_IN.n5 VGND 0.022089f
C1173 I_IN.n6 VGND 0.267792f
C1174 I_IN.t12 VGND 0.010427f
C1175 I_IN.t3 VGND 0.010427f
C1176 I_IN.n7 VGND 0.022089f
C1177 I_IN.n8 VGND 0.267792f
C1178 I_IN.t2 VGND 0.010427f
C1179 I_IN.t4 VGND 0.010427f
C1180 I_IN.n9 VGND 0.022089f
C1181 I_IN.n10 VGND 2.05318f
C1182 I_IN.t16 VGND 0.026069f
C1183 I_IN.t14 VGND 0.026069f
C1184 I_IN.n11 VGND 0.103772f
C1185 I_IN.t15 VGND 0.087787f
C1186 I_IN.t19 VGND 0.113398f
C1187 I_IN.t18 VGND 0.152123f
C1188 I_IN.n12 VGND 0.113824f
C1189 I_IN.n13 VGND 0.11894f
C1190 I_IN.t13 VGND 0.126512f
C1191 I_IN.n14 VGND 0.061648f
C1192 I_IN.n15 VGND 0.167906f
C1193 I_IN.t10 VGND 0.09234f
C1194 I_IN.t7 VGND 0.075732f
C1195 I_IN.n16 VGND 0.159906f
C1196 I_IN.n17 VGND 0.619209f
C1197 a_13750_11850.n0 VGND 0.594039f
C1198 a_13750_11850.n1 VGND 0.475232f
C1199 a_13750_11850.n2 VGND 0.299302f
C1200 a_13750_11850.n3 VGND 0.475232f
C1201 a_13750_11850.n4 VGND 0.846873f
C1202 a_13750_11850.n5 VGND 0.793313f
C1203 a_13750_11850.n6 VGND 2.30308f
C1204 a_13750_11850.n7 VGND 0.116175f
C1205 a_13750_11850.t4 VGND 0.011957f
C1206 a_13750_11850.t13 VGND 0.010511f
C1207 a_13750_11850.t18 VGND 0.010511f
C1208 a_13750_11850.n8 VGND 0.019555f
C1209 a_13750_11850.t21 VGND 0.271561f
C1210 a_13750_11850.t30 VGND 0.276068f
C1211 a_13750_11850.t23 VGND 0.271561f
C1212 a_13750_11850.t19 VGND 0.271561f
C1213 a_13750_11850.t28 VGND 0.271561f
C1214 a_13750_11850.t22 VGND 0.271561f
C1215 a_13750_11850.t33 VGND 0.271561f
C1216 a_13750_11850.t12 VGND 0.271561f
C1217 a_13750_11850.t17 VGND 0.271561f
C1218 a_13750_11850.t14 VGND 0.271561f
C1219 a_13750_11850.t29 VGND 0.271561f
C1220 a_13750_11850.t20 VGND 0.271561f
C1221 a_13750_11850.t26 VGND 0.271561f
C1222 a_13750_11850.t16 VGND 0.271561f
C1223 a_13750_11850.t11 VGND 0.271561f
C1224 a_13750_11850.t31 VGND 0.271561f
C1225 a_13750_11850.t34 VGND 0.271561f
C1226 a_13750_11850.t27 VGND 0.271561f
C1227 a_13750_11850.t32 VGND 0.271561f
C1228 a_13750_11850.t35 VGND 0.271561f
C1229 a_13750_11850.t24 VGND 0.016321f
C1230 a_13750_11850.n9 VGND 0.014381f
C1231 a_13750_11850.t15 VGND 0.016062f
C1232 a_13750_11850.n10 VGND 0.014381f
C1233 a_13750_11850.t36 VGND 0.010511f
C1234 a_13750_11850.t25 VGND 0.010511f
C1235 a_13750_11850.n11 VGND 0.020019f
C1236 a_13750_11850.n12 VGND 0.014381f
C1237 a_13750_11850.n14 VGND 0.22076f
C1238 a_10354_16286.t2 VGND 0.049617f
C1239 a_10354_16286.t5 VGND 0.049617f
C1240 a_10354_16286.n0 VGND 0.123425f
C1241 a_10354_16286.t4 VGND 0.049617f
C1242 a_10354_16286.t3 VGND 0.049617f
C1243 a_10354_16286.n1 VGND 0.11861f
C1244 a_10354_16286.n2 VGND 1.69171f
C1245 a_10354_16286.t10 VGND 0.025428f
C1246 a_10354_16286.t7 VGND 0.025379f
C1247 a_10354_16286.n3 VGND 0.178506f
C1248 a_10354_16286.t6 VGND 0.025379f
C1249 a_10354_16286.n4 VGND 0.110986f
C1250 a_10354_16286.t8 VGND 0.025379f
C1251 a_10354_16286.n5 VGND 0.110986f
C1252 a_10354_16286.t9 VGND 0.025379f
C1253 a_10354_16286.n6 VGND 0.371616f
C1254 a_10354_16286.n7 VGND 0.875787f
C1255 a_10354_16286.t1 VGND 0.144357f
C1256 a_10354_16286.n8 VGND 2.20679f
C1257 a_10354_16286.t0 VGND 0.441816f
.ends

