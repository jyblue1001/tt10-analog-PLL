* PEX produced on Mon Sep  1 08:25:58 PM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from project_magic.ext - technology: sky130A

.subckt project_magic ua[0] ua[1] VDPWR VGND
X0 VDPWR.t343 VDPWR.t340 VDPWR.t342 VDPWR.t341 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X1 VDPWR.t379 a_19190_29050.t11 a_14348_27710.t8 VDPWR.t378 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X2 a_19190_31850.t10 a_19190_31610.t17 VDPWR.t222 VDPWR.t221 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X3 w_13193_29093.t277 a_26300_25010.t3 a_26300_25670.t1 w_13193_29093.t276 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X4 a_18974_25970.t8 a_18974_25060.t8 sky130_fd_pr__res_generic_po w=0.33 l=2.4
X5 a_18180_33430.t8 VDPWR.t428 w_13193_29093.t268 w_13193_29093.t267 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X6 a_14348_27710.t14 VDPWR.t185 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7 a_26640_21760.t0 a_25860_20180.t3 VDPWR.t123 VDPWR.t122 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X8 a_23100_30460.t1 a_24280_30060.t2 VDPWR.t235 VDPWR.t234 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X9 w_13193_29093.t53 w_13193_29093.t104 a_14730_30630.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X10 w_13193_29093.t252 a_19910_25340.t3 a_19910_25340.t4 w_13193_29093.t4 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X11 a_20480_25210.t12 a_19910_24200.t6 a_19040_22530.t2 VDPWR.t251 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X12 VDPWR.t366 a_18974_25970.t9 a_20480_25210.t3 VDPWR.t365 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X13 VDPWR.t263 a_26320_28790.t2 a_26420_30200.t2 VDPWR.t262 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X14 a_19190_29050.t12 a_13532_27710.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X15 a_19940_23090.t6 a_23100_27770.t2 a_23130_27670.t0 w_13193_29093.t150 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X16 a_23100_30980.t1 a_23100_30570.t3 a_23550_30490.t0 VDPWR.t86 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X17 a_19250_24340.t10 a_18974_25060.t9 w_13193_29093.t279 w_13193_29093.t13 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X18 VDPWR.t409 a_19190_29290.t17 a_19190_29050.t10 VDPWR.t408 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X19 a_17540_31010.t5 a_14348_27710.t15 VDPWR.t187 VDPWR.t186 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X20 VDPWR.t339 VDPWR.t337 a_14348_27710.t13 VDPWR.t338 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X21 VDPWR.t37 a_14348_27710.t16 a_14730_30630.t7 VDPWR.t36 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X22 a_14348_27710.t9 VDPWR.t429 w_13193_29093.t266 w_13193_29093.t265 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1.01 ps=6.15 w=2.5 l=5
X23 a_14348_27710.t17 VDPWR.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X24 a_26420_26340.t0 a_26390_26310.t3 a_26420_26230.t0 w_13193_29093.t132 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X25 a_14730_30630.t6 a_14348_27710.t18 VDPWR.t381 VDPWR.t380 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X26 a_19190_29290.t13 a_14730_30630.t8 a_18180_28430.t4 w_13193_29093.t22 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X27 VDPWR.t383 a_14348_27710.t19 a_14990_33500.t4 VDPWR.t382 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X28 w_13193_29093.t103 w_13193_29093.t100 w_13193_29093.t102 w_13193_29093.t101 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X29 a_26310_26200.t0 a_26390_27520.t2 w_13193_29093.t255 w_13193_29093.t254 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X30 a_24310_31390.t0 a_24280_30570.t3 VDPWR.t248 VDPWR.t178 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X31 a_14990_33500.t3 a_14348_27710.t20 VDPWR.t64 VDPWR.t63 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X32 a_24280_31090.t0 a_23100_30050.t3 w_13193_29093.t288 w_13193_29093.t287 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X33 VDPWR.t350 a_24280_31090.t3 a_24310_31010.t0 VDPWR.t245 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X34 w_13193_29093.t217 a_26390_26310.t4 a_26390_28180.t2 w_13193_29093.t216 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X35 a_25860_21760.t0 V_CONT.t8 w_13193_29093.t151 w_13193_29093.t140 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X36 a_19940_24490.t1 V_CONT.t9 a_19250_24340.t13 w_13193_29093.t4 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X37 VDPWR.t128 a_23100_29610.t3 a_23100_29280.t1 VDPWR.t127 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X38 a_22190_29430.t10 a_14558_34050.t10 VDPWR.t345 VDPWR.t344 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X39 w_13193_29093.t280 a_18974_25060.t10 a_19250_24340.t9 w_13193_29093.t13 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X40 VDPWR.t387 a_19190_29290.t18 a_19190_29050.t8 VDPWR.t386 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X41 w_13193_29093.t142 a_23100_30570.t4 a_23100_30980.t0 w_13193_29093.t141 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X42 VDPWR.t360 a_23130_27670.t3 V_CONT.t3 VDPWR.t359 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X43 a_19190_29290.t11 a_19190_29290.t10 VDPWR.t109 VDPWR.t108 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X44 VDPWR.t105 a_19190_31610.t18 a_19190_31850.t9 VDPWR.t104 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X45 a_14348_27710.t21 VDPWR.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X46 a_26300_22300.t0 a_26300_23070.t4 w_13193_29093.t301 w_13193_29093.t300 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X47 w_13193_29093.t249 a_26390_27520.t3 a_26420_27440.t1 w_13193_29093.t248 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X48 w_13193_29093.t20 a_26310_26200.t3 a_26390_29930.t3 w_13193_29093.t19 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X49 a_14348_27710.t22 VDPWR.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X50 a_20480_25210.t9 a_20480_25210.t7 a_20480_25210.t8 VDPWR.t247 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X51 VDPWR.t220 a_14558_34050.t11 a_14140_28370.t10 VDPWR.t219 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X52 a_26310_26200.t2 a_26390_27520.t4 VDPWR.t352 VDPWR.t351 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X53 a_26390_31270.t3 a_26310_26200.t4 w_13193_29093.t290 w_13193_29093.t289 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X54 w_13193_29093.t112 a_19040_22530.t5 a_19940_23090.t4 w_13193_29093.t111 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X55 w_13193_29093.t53 w_13193_29093.t99 a_13370_29270.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X56 a_24280_31990.t0 a_26320_28790.t3 VDPWR.t259 VDPWR.t258 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X57 w_13193_29093.t51 a_23100_29610.t4 a_23100_29280.t0 w_13193_29093.t50 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X58 VDPWR.t40 a_19190_31610.t19 a_19190_31850.t8 VDPWR.t39 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X59 a_26640_21160.t1 w_13193_29093.t313 VDPWR.t67 VDPWR.t66 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X60 a_19910_24200.t4 a_19940_23090.t10 VDPWR.t362 VDPWR.t361 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X61 a_22190_29430.t0 a_24280_27770.t2 a_24310_27670.t2 VDPWR.t97 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X62 a_24280_29730.t1 a_23130_29200.t2 VDPWR.t208 VDPWR.t207 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X63 a_26300_23600.t1 a_26300_24370.t4 w_13193_29093.t251 w_13193_29093.t250 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X64 a_14558_34050.t9 a_19190_31850.t11 VDPWR.t204 VDPWR.t203 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X65 w_13193_29093.t247 a_26390_30500.t2 a_26420_30420.t1 w_13193_29093.t246 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X66 w_13193_29093.t264 VDPWR.t430 a_14558_34050.t1 w_13193_29093.t263 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X67 a_14348_27710.t23 VDPWR.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X68 VDPWR.t336 VDPWR.t334 a_14348_27710.t12 VDPWR.t335 sky130_fd_pr__pfet_01v8 ad=0.45 pd=2.9 as=0.2 ps=1.4 w=1 l=0.15
X69 a_25860_21760.t1 ua[1].t2 a_26400_21130.t1 w_13193_29093.t140 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X70 a_26420_27220.t1 a_26390_27520.t5 VDPWR.t257 VDPWR.t256 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X71 VDPWR.t92 a_19940_24490.t4 a_19940_24490.t5 VDPWR.t91 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X72 a_26390_32300.t3 a_26320_28790.t4 w_13193_29093.t8 w_13193_29093.t7 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X73 a_26320_28790.t0 a_26310_26200.t5 VDPWR.t83 VDPWR.t82 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X74 VDPWR.t119 ua[0].t0 a_23550_31910.t0 VDPWR.t118 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X75 a_14348_27710.t7 a_19190_29050.t13 VDPWR.t399 VDPWR.t398 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X76 VDPWR.t141 a_23100_29280.t2 a_23130_29200.t1 VDPWR.t140 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X77 a_19190_31850.t4 a_14140_28370.t13 a_18180_33430.t5 w_13193_29093.t139 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X78 VDPWR.t206 a_19190_29290.t8 a_19190_29290.t9 VDPWR.t205 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X79 a_26300_24900.t0 a_26300_25670.t4 w_13193_29093.t106 w_13193_29093.t105 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X80 a_24280_30980.t1 a_24280_30570.t4 a_24310_30490.t0 VDPWR.t86 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X81 a_26640_20560.t2 a_26400_20530.t2 ua[1].t1 VDPWR.t59 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X82 a_14348_27710.t24 VDPWR.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X83 a_22190_29430.t9 a_14558_34050.t12 VDPWR.t354 VDPWR.t353 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X84 w_13193_29093.t98 w_13193_29093.t96 w_13193_29093.t97 w_13193_29093.t4 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X85 a_26740_30530.t1 a_26390_30500.t3 VDPWR.t212 VDPWR.t211 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X86 a_18974_25970.t7 a_18974_25970.t6 VDPWR.t161 VDPWR.t160 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X87 a_23100_30460.t0 a_24280_30060.t3 w_13193_29093.t225 w_13193_29093.t224 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X88 a_14140_28370.t12 VDPWR.t331 VDPWR.t333 VDPWR.t332 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X89 w_13193_29093.t95 w_13193_29093.t93 w_13193_29093.t94 w_13193_29093.t4 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X90 VDPWR.t369 a_23100_30050.t4 a_23100_29610.t0 VDPWR.t368 sky130_fd_pr__pfet_01v8 ad=0.805 pd=5 as=0.4 ps=2.4 w=2 l=0.15
X91 w_13193_29093.t163 ua[0].t1 a_23020_31090.t0 w_13193_29093.t162 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X92 a_19190_29050.t14 a_13532_27710.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X93 VDPWR.t330 VDPWR.t327 VDPWR.t329 VDPWR.t328 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X94 a_19190_31610.t14 a_19190_31610.t13 VDPWR.t28 VDPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X95 w_13193_29093.t155 a_23100_29280.t3 a_23130_29200.t0 w_13193_29093.t154 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X96 w_13193_29093.t135 ua[1].t3 a_26300_22410.t0 w_13193_29093.t134 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X97 w_13193_29093.t190 a_26390_26310.t5 a_26390_26970.t2 w_13193_29093.t189 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X98 VDPWR.t192 a_19190_31850.t12 a_14558_34050.t8 VDPWR.t191 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X99 a_14348_27710.t25 VDPWR.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X100 V_CONT.t7 a_25350_8708.t1 w_13193_29093.t245 sky130_fd_pr__res_xhigh_po_0p35 l=7.52
X101 a_19190_29050.t15 a_13532_27710.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X102 w_13193_29093.t294 a_24280_27770.t3 a_24310_27670.t1 w_13193_29093.t293 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X103 a_18180_28430.t7 a_14990_33500.t6 a_19190_29050.t3 w_13193_29093.t215 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X104 VDPWR.t326 VDPWR.t323 VDPWR.t325 VDPWR.t324 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0 ps=0 w=2.5 l=0.5
X105 a_23100_30050.t0 a_24280_30570.t5 w_13193_29093.t46 w_13193_29093.t45 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X106 VDPWR.t322 VDPWR.t320 a_14140_28370.t11 VDPWR.t321 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X107 a_19190_31850.t13 a_13742_34050.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X108 a_23100_29610.t2 a_23020_29890.t3 VDPWR.t397 VDPWR.t396 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X109 w_13193_29093.t239 a_24280_31090.t4 a_24280_30570.t2 w_13193_29093.t238 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X110 a_19190_29050.t16 a_13532_27710.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X111 VDPWR.t50 a_19190_29050.t17 a_14348_27710.t6 VDPWR.t49 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X112 w_13193_29093.t175 a_23100_30050.t5 a_23130_29970.t0 w_13193_29093.t174 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X113 a_18180_33430.t4 a_14140_28370.t14 a_19190_31850.t3 w_13193_29093.t133 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X114 w_13193_29093.t121 a_26300_22300.t2 a_26300_23710.t0 w_13193_29093.t120 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X115 a_19190_29050.t0 a_19190_29290.t19 VDPWR.t152 VDPWR.t151 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X116 a_14348_27710.t26 VDPWR.t188 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X117 w_13193_29093.t42 a_26390_26310.t6 a_26390_28180.t1 w_13193_29093.t41 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X118 a_18180_28430.t8 a_14990_33500.t7 a_19190_29050.t6 w_13193_29093.t218 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X119 a_13532_33810.t1 a_14610_33690.t1 w_13193_29093.t253 sky130_fd_pr__res_xhigh_po_0p35 l=3.35
X120 a_19190_29050.t18 a_13532_27710.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X121 a_19910_25340.t2 a_19910_25340.t1 w_13193_29093.t38 w_13193_29093.t4 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X122 a_19190_31850.t14 a_13742_34050.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X123 a_19040_22530.t3 a_19910_24200.t7 a_20480_25210.t11 VDPWR.t177 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X124 V_CONT.t2 a_23130_27670.t4 VDPWR.t7 VDPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X125 a_26300_23070.t2 a_26300_22410.t3 w_13193_29093.t167 w_13193_29093.t166 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X126 a_23130_29970.t1 a_23020_29890.t4 a_23100_29610.t1 w_13193_29093.t128 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X127 a_26640_21760.t1 w_13193_29093.t314 VDPWR.t69 VDPWR.t68 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X128 a_19190_31850.t15 a_13742_34050.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X129 a_18974_25060.t7 a_18974_25060.t6 w_13193_29093.t28 w_13193_29093.t13 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X130 VDPWR.t230 a_19190_31610.t11 a_19190_31610.t12 VDPWR.t229 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X131 w_13193_29093.t123 a_26300_23600.t2 a_26300_25010.t1 w_13193_29093.t122 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X132 a_24280_30060.t0 a_24280_29730.t2 VDPWR.t393 VDPWR.t392 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X133 VDPWR.t416 a_24280_31990.t2 a_24310_31910.t1 VDPWR.t118 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X134 a_19190_29050.t19 a_13532_27710.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X135 a_19190_31850.t7 a_19190_31610.t20 VDPWR.t42 VDPWR.t41 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X136 V_CONT.t6 a_24310_27670.t3 w_13193_29093.t159 w_13193_29093.t158 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X137 a_22190_29430.t15 a_24310_27960.t3 a_24310_27670.t0 w_13193_29093.t199 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X138 a_24280_29730.t0 a_23130_29200.t3 w_13193_29093.t232 w_13193_29093.t231 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X139 VDPWR.t395 a_26420_27220.t3 a_26390_28180.t3 VDPWR.t394 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X140 a_26390_29240.t0 a_26320_28790.t5 w_13193_29093.t177 w_13193_29093.t176 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X141 a_19250_24340.t11 a_19910_24200.t8 a_19940_24230.t4 w_13193_29093.t4 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X142 VDPWR.t319 VDPWR.t316 VDPWR.t318 VDPWR.t317 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X143 a_22190_29430.t8 a_14558_34050.t13 VDPWR.t265 VDPWR.t264 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X144 a_19190_29050.t20 a_13532_27710.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X145 a_14140_28370.t9 a_14558_34050.t14 VDPWR.t143 VDPWR.t142 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X146 a_19190_31850.t16 a_13742_34050.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X147 w_13193_29093.t92 w_13193_29093.t90 w_13193_29093.t91 w_13193_29093.t13 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0 ps=0 w=1.25 l=0.5
X148 a_23020_29890.t2 a_23020_31090.t3 a_23550_31390.t1 VDPWR.t124 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X149 a_13370_29270.t8 a_14990_33500.t5 w_13193_29093.t278 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X150 a_19190_29290.t7 a_19190_29290.t6 VDPWR.t3 VDPWR.t2 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X151 a_18180_28430.t9 a_14990_33500.t8 a_19190_29050.t7 w_13193_29093.t219 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X152 a_19190_31850.t6 a_19190_31610.t21 VDPWR.t356 VDPWR.t355 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X153 a_19190_29050.t21 a_13532_27710.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X154 a_26420_27330.t0 a_26390_26310.t7 a_26420_27220.t0 w_13193_29093.t230 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X155 VDPWR.t315 VDPWR.t313 a_14610_33930.t6 VDPWR.t314 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X156 w_13193_29093.t44 a_26310_26200.t6 a_26390_29930.t2 w_13193_29093.t43 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X157 w_13193_29093.t18 a_22190_29430.t18 a_19910_24200.t1 w_13193_29093.t17 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X158 a_19190_29290.t15 a_14730_30630.t9 a_18180_28430.t3 w_13193_29093.t23 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X159 a_13532_33810.t0 a_14610_33930.t0 w_13193_29093.t27 sky130_fd_pr__res_xhigh_po_0p35 l=3.35
X160 a_14610_33930.t4 a_14348_27710.t27 VDPWR.t190 VDPWR.t189 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X161 a_18180_33430.t10 a_14610_33930.t7 a_19190_31610.t16 w_13193_29093.t295 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X162 a_20480_25210.t13 V_CONT.t10 a_19910_25340.t5 VDPWR.t250 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X163 VDPWR.t232 a_14348_27710.t28 a_17540_31010.t4 VDPWR.t231 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X164 a_26420_29270.t0 a_26390_29240.t3 w_13193_29093.t198 w_13193_29093.t197 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X165 VDPWR.t242 a_14558_34050.t15 a_22190_29430.t7 VDPWR.t241 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X166 w_13193_29093.t292 a_24280_30570.t6 a_24280_30980.t0 w_13193_29093.t291 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X167 VDPWR.t267 a_14558_34050.t16 a_14140_28370.t8 VDPWR.t266 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X168 a_14348_27710.t29 VDPWR.t233 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X169 a_19940_23090.t3 a_19040_22530.t6 w_13193_29093.t184 w_13193_29093.t183 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X170 VDPWR.t163 a_26320_28790.t6 a_26390_29240.t2 VDPWR.t162 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X171 a_26330_22330.t1 a_26300_22300.t3 w_13193_29093.t153 w_13193_29093.t152 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X172 w_13193_29093.t234 a_23020_31090.t4 a_23020_29890.t1 w_13193_29093.t233 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X173 VDPWR.t238 a_19940_23090.t11 a_19910_24200.t3 VDPWR.t237 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X174 a_14558_34050.t7 a_19190_31850.t17 VDPWR.t44 VDPWR.t43 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X175 a_19190_29050.t22 a_13532_27710.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X176 a_26390_27410.t1 a_26390_26970.t4 w_13193_29093.t309 w_13193_29093.t308 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X177 a_26300_24370.t0 a_26300_23710.t3 w_13193_29093.t30 w_13193_29093.t29 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X178 a_18180_33430.t2 a_14140_28370.t15 a_19190_31850.t2 w_13193_29093.t107 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X179 a_14730_30630.t3 a_17540_31010.t6 a_14348_27710.t2 VDPWR.t236 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X180 w_13193_29093.t315 a_25350_8708.t0 sky130_fd_pr__cap_mim_m3_1 l=69.8 w=60
X181 a_26640_21160.t2 a_26400_21130.t2 a_26400_20530.t1 VDPWR.t66 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X182 a_19250_24340.t6 a_19250_24340.t4 a_19250_24340.t5 w_13193_29093.t4 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X183 a_19190_31610.t0 a_14610_33930.t8 a_18180_33430.t3 w_13193_29093.t130 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X184 a_19940_24490.t3 a_19940_24490.t2 VDPWR.t20 VDPWR.t19 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X185 a_14348_27710.t30 VDPWR.t376 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X186 VDPWR.t424 a_26390_29240.t4 a_26420_29380.t0 VDPWR.t423 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X187 a_19190_31850.t18 a_13742_34050.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X188 VDPWR.t46 a_18974_25970.t10 a_20480_25210.t2 VDPWR.t45 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X189 a_26330_23630.t1 a_26300_23600.t3 w_13193_29093.t161 w_13193_29093.t160 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X190 w_13193_29093.t53 w_13193_29093.t75 a_13370_29270.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X191 VDPWR.t62 a_26300_22300.t4 a_26330_22440.t1 VDPWR.t61 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X192 a_19190_29290.t12 a_14730_30630.t10 a_18180_28430.t2 w_13193_29093.t210 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X193 a_26300_25670.t3 a_26300_25010.t4 w_13193_29093.t275 w_13193_29093.t274 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X194 VDPWR.t358 a_19190_31610.t22 a_19190_31850.t5 VDPWR.t357 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X195 VDPWR.t375 ua[1].t4 a_26300_22410.t2 VDPWR.t374 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X196 a_18180_28430.t1 a_14730_30630.t11 a_19190_29290.t14 w_13193_29093.t211 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X197 w_13193_29093.t270 a_19040_22530.t7 a_19940_23090.t2 w_13193_29093.t269 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X198 a_22190_29430.t17 VDPWR.t310 VDPWR.t312 VDPWR.t311 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X199 w_13193_29093.t244 a_14610_33690.t0 w_13193_29093.t243 sky130_fd_pr__res_xhigh_po_0p35 l=3.35
X200 VDPWR.t198 a_19940_24230.t5 a_19940_23090.t7 VDPWR.t197 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X201 w_13193_29093.t89 w_13193_29093.t86 w_13193_29093.t88 w_13193_29093.t87 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X202 a_18974_25970.t5 a_18974_25970.t4 VDPWR.t150 VDPWR.t149 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X203 w_13193_29093.t226 a_18974_25060.t11 a_19250_24340.t8 w_13193_29093.t13 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X204 VDPWR.t155 a_23100_27770.t3 a_23130_27960.t2 VDPWR.t32 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X205 a_26330_24930.t0 a_26300_24900.t2 w_13193_29093.t165 w_13193_29093.t164 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X206 VDPWR.t96 a_26300_23600.t4 a_26330_23740.t1 VDPWR.t95 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X207 w_13193_29093.t53 w_13193_29093.t76 a_13370_29270.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X208 VDPWR.t364 a_19190_31850.t19 a_14558_34050.t6 VDPWR.t363 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X209 a_26300_22300.t1 a_26300_22410.t4 VDPWR.t74 VDPWR.t73 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X210 a_19190_31610.t1 a_14610_33930.t9 a_18180_33430.t6 w_13193_29093.t170 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X211 VDPWR.t71 a_26300_22300.t5 a_26300_23710.t2 VDPWR.t70 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X212 a_23100_30050.t2 a_24280_31090.t5 a_24310_31390.t1 VDPWR.t124 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X213 a_24280_30060.t1 a_24280_29730.t3 w_13193_29093.t303 w_13193_29093.t302 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X214 w_13193_29093.t157 a_24280_31990.t3 a_24280_31090.t2 w_13193_29093.t156 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X215 a_18180_33430.t9 a_14610_33930.t10 a_19190_31610.t15 w_13193_29093.t286 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X216 a_19940_23090.t12 a_18460_22530.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X217 a_26390_27520.t1 a_26390_28180.t4 w_13193_29093.t173 w_13193_29093.t172 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X218 a_19940_23090.t13 a_21386_22530.t1 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X219 VDPWR.t244 a_14558_34050.t17 a_22190_29430.t6 VDPWR.t243 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X220 a_18974_25060.t5 a_18974_25060.t4 w_13193_29093.t182 w_13193_29093.t13 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X221 w_13193_29093.t194 a_23100_27770.t4 a_23130_27960.t1 w_13193_29093.t193 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X222 VDPWR.t309 VDPWR.t307 a_14558_34050.t3 VDPWR.t308 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X223 a_26300_23600.t0 a_26300_23710.t4 VDPWR.t111 VDPWR.t110 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X224 a_18180_28430.t0 a_14730_30630.t12 a_19190_29290.t16 w_13193_29093.t310 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X225 a_19190_31610.t10 a_19190_31610.t9 VDPWR.t157 VDPWR.t156 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X226 a_26390_30500.t0 a_26390_29930.t4 w_13193_29093.t119 w_13193_29093.t118 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X227 VDPWR.t90 a_26300_23600.t5 a_26300_25010.t0 VDPWR.t89 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X228 a_19190_29050.t2 a_14990_33500.t9 a_18180_28430.t6 w_13193_29093.t202 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X229 a_26420_31640.t0 a_24280_31990.t4 w_13193_29093.t283 w_13193_29093.t282 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X230 a_26390_29240.t1 a_26320_28790.t7 VDPWR.t11 VDPWR.t10 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X231 a_19190_29050.t23 a_13532_27710.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X232 VDPWR.t306 VDPWR.t303 VDPWR.t305 VDPWR.t304 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X233 a_20480_25210.t6 a_20480_25210.t4 a_20480_25210.t5 VDPWR.t249 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X234 a_13742_34050.t0 a_14558_34050.t0 w_13193_29093.t214 sky130_fd_pr__res_high_po_0p35 l=2.05
X235 a_14140_28370.t7 a_14558_34050.t18 VDPWR.t165 VDPWR.t164 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X236 VDPWR.t126 a_26390_27520.t6 a_26310_26200.t1 VDPWR.t125 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X237 w_13193_29093.t188 a_26310_26200.t7 a_26390_31270.t2 w_13193_29093.t187 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X238 a_14348_27710.t31 VDPWR.t377 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X239 VDPWR.t144 a_23100_28450.t2 a_23100_27770.t0 VDPWR.t58 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X240 a_23550_31010.t1 a_23100_30980.t3 a_23100_30570.t2 VDPWR.t216 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X241 VDPWR.t24 a_23130_27670.t5 V_CONT.t1 VDPWR.t23 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X242 a_19940_24230.t2 a_21386_22530.t0 w_13193_29093.t213 sky130_fd_pr__res_xhigh_po_0p35 l=1.14
X243 a_24310_27670.t4 a_24310_27960.t2 sky130_fd_pr__cap_mim_m3_1 l=2.7 w=3.8
X244 a_26300_24900.t1 a_26300_25010.t5 VDPWR.t391 VDPWR.t390 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X245 w_13193_29093.t85 w_13193_29093.t82 w_13193_29093.t84 w_13193_29093.t83 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X246 a_26420_30420.t0 a_24280_31990.t5 w_13193_29093.t34 w_13193_29093.t33 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X247 a_26640_21760.t2 ua[1].t5 a_26400_21130.t0 VDPWR.t68 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X248 w_13193_29093.t81 w_13193_29093.t78 w_13193_29093.t80 w_13193_29093.t79 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X249 a_18180_33430.t7 a_14610_33930.t11 a_19190_31610.t2 w_13193_29093.t212 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X250 a_19190_29050.t24 a_13532_27710.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X251 w_13193_29093.t285 a_26300_24900.t3 a_26390_26310.t2 w_13193_29093.t284 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X252 VDPWR.t57 a_26300_24900.t4 a_26330_25040.t0 VDPWR.t56 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X253 a_19190_31850.t0 a_14140_28370.t16 a_18180_33430.t0 w_13193_29093.t21 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X254 a_19940_24230.t3 a_19910_24200.t9 a_19250_24340.t12 w_13193_29093.t4 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X255 VDPWR.t52 a_24280_31990.t6 a_26420_31750.t0 VDPWR.t51 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X256 w_13193_29093.t53 w_13193_29093.t77 a_13370_29270.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X257 a_14348_27710.t32 VDPWR.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X258 w_13193_29093.t10 a_26320_28790.t8 a_26390_32300.t2 w_13193_29093.t9 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X259 w_13193_29093.t147 a_23100_28450.t3 a_23100_27770.t1 w_13193_29093.t146 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X260 a_23100_30570.t1 a_23100_30980.t4 w_13193_29093.t229 w_13193_29093.t228 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X261 a_19190_31850.t20 a_13742_34050.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X262 a_26300_22410.t1 ua[1].t6 VDPWR.t418 VDPWR.t417 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X263 a_14730_30630.t5 a_14348_27710.t33 VDPWR.t133 VDPWR.t132 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X264 a_26390_27410.t0 a_26390_26310.t8 VDPWR.t22 VDPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X265 a_19190_29050.t1 a_14990_33500.t10 a_18180_28430.t5 w_13193_29093.t149 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X266 VDPWR.t33 a_24280_27770.t4 a_24310_27960.t1 VDPWR.t32 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X267 VDPWR.t181 a_19190_31610.t7 a_19190_31610.t8 VDPWR.t180 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X268 a_19190_29050.t25 a_13532_27710.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X269 a_19910_24200.t2 a_22190_29430.t19 w_13193_29093.t221 w_13193_29093.t220 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X270 a_19190_31850.t21 a_13742_34050.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X271 a_19910_25340.t0 V_CONT.t11 a_20480_25210.t10 VDPWR.t81 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X272 VDPWR.t261 a_26310_26200.t8 a_26420_26340.t1 VDPWR.t260 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X273 VDPWR.t427 a_14558_34050.t19 a_22190_29430.t5 VDPWR.t426 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X274 w_13193_29093.t53 w_13193_29093.t74 a_13370_29270.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X275 a_26420_30200.t0 a_24280_31990.t7 a_26740_30530.t0 VDPWR.t12 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X276 VDPWR.t171 a_14558_34050.t20 a_14140_28370.t6 VDPWR.t170 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X277 VDPWR.t18 a_26300_24900.t5 a_26390_26310.t0 VDPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X278 VDPWR.t148 a_23020_29890.t5 a_23100_28450.t1 VDPWR.t147 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X279 a_19190_31850.t22 a_13742_34050.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X280 a_26300_23710.t1 a_26300_22300.t6 VDPWR.t88 VDPWR.t87 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X281 w_13193_29093.t73 w_13193_29093.t70 w_13193_29093.t72 w_13193_29093.t71 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X282 a_19910_24200.t0 a_19940_23090.t14 VDPWR.t1 VDPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X283 a_26390_26970.t1 a_26390_26310.t9 w_13193_29093.t204 w_13193_29093.t203 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X284 a_19190_29050.t26 a_13532_27710.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X285 a_19190_31850.t23 a_13742_34050.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X286 w_13193_29093.t1 a_22190_29430.t13 a_22190_29430.t14 w_13193_29093.t0 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X287 w_13193_29093.t26 a_14140_28370.t0 w_13193_29093.t25 sky130_fd_pr__res_xhigh_po_0p35 l=1
X288 a_19190_31850.t1 a_14140_28370.t17 a_18180_33430.t1 w_13193_29093.t47 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X289 VDPWR.t176 a_19940_24490.t6 a_19940_24230.t1 VDPWR.t175 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X290 a_22190_29430.t4 a_14558_34050.t21 VDPWR.t218 VDPWR.t217 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X291 a_26420_30310.t1 a_26310_26200.t9 a_26420_30200.t1 w_13193_29093.t148 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X292 w_13193_29093.t12 a_24280_31090.t6 a_23100_30050.t1 w_13193_29093.t11 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X293 a_18460_22530.t1 a_19040_22530.t4 w_13193_29093.t281 sky130_fd_pr__res_xhigh_po_0p35 l=0.86
X294 a_25860_20560.t2 VDPWR.t431 w_13193_29093.t262 w_13193_29093.t129 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X295 w_13193_29093.t53 w_13193_29093.t58 a_13370_29270.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X296 a_19190_29050.t27 a_13532_27710.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X297 w_13193_29093.t169 a_23020_29890.t6 a_23100_28450.t0 w_13193_29093.t168 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X298 VDPWR.t146 a_18974_25970.t2 a_18974_25970.t3 VDPWR.t145 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X299 a_26300_25010.t2 a_26300_23600.t6 VDPWR.t210 VDPWR.t209 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X300 a_24310_28480.t2 w_13193_29093.t316 a_24280_27770.t0 VDPWR.t58 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X301 a_24310_31010.t1 a_24280_30980.t3 a_24280_30570.t1 VDPWR.t216 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X302 a_19190_29050.t28 a_13532_27710.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X303 a_26390_28180.t0 a_26390_26310.t10 w_13193_29093.t181 w_13193_29093.t180 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X304 a_19190_31850.t24 a_13742_34050.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X305 a_14558_34050.t5 a_19190_31850.t25 VDPWR.t401 VDPWR.t400 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X306 a_19940_23090.t1 a_19040_22530.t8 w_13193_29093.t186 w_13193_29093.t185 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X307 a_19940_23090.t0 a_19940_24230.t6 VDPWR.t9 VDPWR.t8 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X308 a_19190_29050.t29 a_13532_27710.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X309 a_20480_25210.t1 a_18974_25970.t11 VDPWR.t48 VDPWR.t47 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X310 a_19190_31850.t26 a_13742_34050.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X311 a_23550_30490.t1 a_23100_30460.t2 VDPWR.t425 VDPWR.t223 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X312 w_13193_29093.t127 a_26300_22410.t5 a_26300_23070.t1 w_13193_29093.t126 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X313 w_13193_29093.t14 a_18974_25060.t2 a_18974_25060.t3 w_13193_29093.t13 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X314 a_14348_27710.t34 VDPWR.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X315 VDPWR.t302 VDPWR.t299 VDPWR.t301 VDPWR.t300 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X316 a_19190_31850.t27 a_13742_34050.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X317 a_26420_26230.t1 a_26310_26200.t10 w_13193_29093.t299 w_13193_29093.t298 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X318 a_26640_20560.t0 a_25860_20180.t4 VDPWR.t99 VDPWR.t98 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X319 w_13193_29093.t40 a_26310_26200.t11 a_26390_31270.t1 w_13193_29093.t39 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X320 VDPWR.t298 VDPWR.t295 VDPWR.t297 VDPWR.t296 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X321 a_26390_27520.t0 a_26390_26310.t11 VDPWR.t154 VDPWR.t153 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X322 a_24280_31990.t1 a_26390_32300.t4 w_13193_29093.t307 w_13193_29093.t306 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X323 VDPWR.t255 a_14558_34050.t22 a_22190_29430.t3 VDPWR.t254 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X324 a_19250_24340.t7 a_18974_25060.t12 w_13193_29093.t227 w_13193_29093.t13 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X325 VDPWR.t167 a_14558_34050.t23 a_14140_28370.t5 VDPWR.t166 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X326 a_14348_27710.t35 VDPWR.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X327 a_23100_30980.t2 a_23100_30460.t3 w_13193_29093.t144 w_13193_29093.t143 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X328 VDPWR.t367 a_23100_30050.t6 a_24310_28480.t1 VDPWR.t147 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X329 a_19190_31850.t28 a_13742_34050.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X330 a_26420_27440.t0 a_26390_27410.t2 a_26420_27330.t1 w_13193_29093.t237 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X331 a_26390_29930.t1 a_26310_26200.t12 w_13193_29093.t16 w_13193_29093.t15 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X332 VDPWR.t113 a_19940_24230.t7 a_19940_23090.t5 VDPWR.t112 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X333 a_26390_26310.t1 a_26300_24900.t6 VDPWR.t35 VDPWR.t34 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X334 w_13193_29093.t137 a_26320_28790.t9 a_26390_32300.t1 w_13193_29093.t136 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X335 w_13193_29093.t114 a_24280_27770.t5 a_24310_27960.t0 w_13193_29093.t113 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X336 a_26420_29380.t1 a_26310_26200.t13 a_26420_29270.t1 w_13193_29093.t205 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X337 VDPWR.t194 a_26420_30200.t3 a_26390_31270.t0 VDPWR.t193 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X338 a_14140_28370.t4 a_14558_34050.t24 VDPWR.t347 VDPWR.t346 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X339 a_25860_20560.t0 V_CONT.t12 w_13193_29093.t256 w_13193_29093.t129 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X340 w_13193_29093.t32 V_CONT.t13 a_25860_20180.t0 w_13193_29093.t31 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X341 w_13193_29093.t110 a_19910_25340.t6 a_19040_22530.t1 w_13193_29093.t4 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X342 a_26330_22440.t0 a_26300_22410.t6 a_26330_22330.t0 w_13193_29093.t115 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X343 VDPWR.t130 a_19190_29050.t30 a_14348_27710.t5 VDPWR.t129 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X344 w_13193_29093.t305 a_26300_23710.t5 a_26300_24370.t3 w_13193_29093.t304 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X345 a_14348_27710.t1 a_17540_31010.t7 a_14730_30630.t0 VDPWR.t72 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X346 VDPWR.t385 a_26390_27410.t3 a_26420_27220.t2 VDPWR.t384 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X347 VDPWR.t294 VDPWR.t291 VDPWR.t293 VDPWR.t292 sky130_fd_pr__pfet_01v8 ad=1.25 pd=6 as=0 ps=0 w=2.5 l=0.5
X348 a_26390_29930.t0 a_26420_29380.t2 VDPWR.t76 VDPWR.t75 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X349 a_14348_27710.t36 VDPWR.t182 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X350 a_23550_31910.t1 a_23020_29890.t7 a_23020_31090.t2 VDPWR.t174 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X351 a_26330_23740.t0 a_26300_23710.t6 a_26330_23630.t0 w_13193_29093.t145 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X352 a_14610_33930.t3 a_14348_27710.t37 VDPWR.t184 VDPWR.t183 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X353 a_26300_23070.t3 a_26330_22440.t2 VDPWR.t202 VDPWR.t201 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X354 VDPWR.t420 a_14348_27710.t38 a_14990_33500.t2 VDPWR.t419 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X355 w_13193_29093.t273 a_26300_25010.t6 a_26300_25670.t2 w_13193_29093.t272 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X356 a_24310_30490.t1 a_23100_30460.t4 VDPWR.t224 VDPWR.t223 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X357 a_14990_33500.t1 a_14348_27710.t39 VDPWR.t422 VDPWR.t421 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X358 VDPWR.t214 a_14348_27710.t40 a_14730_30630.t4 VDPWR.t213 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X359 w_13193_29093.t69 w_13193_29093.t66 w_13193_29093.t68 w_13193_29093.t67 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X360 a_13382_33380.t0 a_14990_33500.t0 w_13193_29093.t6 sky130_fd_pr__res_xhigh_po_0p35 l=6
X361 a_25860_20560.t1 a_26400_20530.t3 ua[1].t0 w_13193_29093.t129 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X362 a_24280_30570.t0 a_24280_30980.t4 w_13193_29093.t125 w_13193_29093.t124 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X363 a_24310_28480.t3 VDPWR.t432 a_24280_27770.t1 w_13193_29093.t261 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X364 VDPWR.t173 a_14558_34050.t25 a_22190_29430.t2 VDPWR.t172 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X365 w_13193_29093.t65 w_13193_29093.t63 w_13193_29093.t64 w_13193_29093.t4 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X366 VDPWR.t403 a_18974_25970.t0 a_18974_25970.t1 VDPWR.t402 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X367 a_17540_31010.t1 a_17540_31010.t0 a_17540_28930.t0 w_13193_29093.t37 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X368 a_25860_21160.t1 VDPWR.t433 w_13193_29093.t260 w_13193_29093.t195 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X369 w_13193_29093.t62 w_13193_29093.t60 w_13193_29093.t61 w_13193_29093.t13 sky130_fd_pr__nfet_01v8 ad=0.625 pd=3.5 as=0 ps=0 w=1.25 l=0.5
X370 a_13532_27710.t0 a_14348_27710.t0 w_13193_29093.t5 sky130_fd_pr__res_high_po_0p35 l=2.05
X371 a_19190_29290.t5 a_19190_29290.t4 VDPWR.t411 VDPWR.t410 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X372 a_23020_31090.t1 a_23020_29890.t8 w_13193_29093.t209 w_13193_29093.t208 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X373 a_19190_29050.t4 a_19190_29290.t20 VDPWR.t226 VDPWR.t225 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X374 a_14348_27710.t41 VDPWR.t215 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X375 w_13193_29093.t36 a_24310_27670.t5 V_CONT.t4 w_13193_29093.t35 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X376 a_13382_28490.t1 a_14990_28610.t1 w_13193_29093.t242 sky130_fd_pr__res_xhigh_po_0p35 l=6
X377 a_26640_21160.t0 a_25860_20180.t5 VDPWR.t101 VDPWR.t100 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X378 a_26300_24370.t1 a_26330_23740.t2 VDPWR.t78 VDPWR.t77 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X379 VDPWR.t290 VDPWR.t287 VDPWR.t289 VDPWR.t288 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X380 VDPWR.t30 a_14348_27710.t42 a_14610_33930.t2 VDPWR.t29 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X381 a_22190_29430.t12 a_22190_29430.t11 w_13193_29093.t117 w_13193_29093.t116 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X382 a_19190_31850.t29 a_13742_34050.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X383 a_19940_24230.t0 a_19940_24490.t7 VDPWR.t137 VDPWR.t136 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X384 a_23130_27670.t6 a_23130_27960.t0 sky130_fd_pr__cap_mim_m3_1 l=5.2 w=6.3
X385 a_14140_28370.t3 a_14558_34050.t26 VDPWR.t349 VDPWR.t348 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X386 a_19250_24340.t0 V_CONT.t14 a_19940_24490.t0 w_13193_29093.t4 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X387 w_13193_29093.t171 a_18974_25060.t0 a_18974_25060.t1 w_13193_29093.t13 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X388 a_14348_27710.t43 VDPWR.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X389 a_14558_34050.t2 VDPWR.t284 VDPWR.t286 VDPWR.t285 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X390 VDPWR.t405 a_25860_20180.t1 a_25860_20180.t2 VDPWR.t404 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X391 VDPWR.t283 VDPWR.t280 VDPWR.t282 VDPWR.t281 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X392 a_26330_25040.t1 a_26300_25010.t7 a_26330_24930.t1 w_13193_29093.t271 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X393 w_13193_29093.t192 a_23100_30050.t7 a_24310_28480.t0 w_13193_29093.t191 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X394 a_26420_31750.t1 a_26320_28790.t10 a_26420_31640.t1 w_13193_29093.t138 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X395 a_19190_31850.t30 a_13742_34050.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X396 w_13193_29093.t297 a_14990_33260.t1 w_13193_29093.t296 sky130_fd_pr__res_xhigh_po_0p35 l=6
X397 a_26320_28790.t1 a_26390_31270.t4 w_13193_29093.t312 w_13193_29093.t311 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X398 a_19190_29050.t31 a_13532_27710.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X399 w_13193_29093.t109 a_26300_22410.t7 a_26300_23070.t0 w_13193_29093.t108 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X400 VDPWR.t107 a_19190_29290.t2 a_19190_29290.t3 VDPWR.t106 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X401 VDPWR.t407 a_19190_29290.t21 a_19190_29050.t9 VDPWR.t406 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X402 VDPWR.t413 a_19940_23090.t15 a_19910_24200.t5 VDPWR.t412 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X403 a_14348_27710.t11 VDPWR.t277 VDPWR.t279 VDPWR.t278 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X404 w_13193_29093.t179 a_14990_28610.t0 w_13193_29093.t178 sky130_fd_pr__res_xhigh_po_0p35 l=6
X405 a_24310_31910.t0 a_23100_30050.t8 a_24280_31090.t1 VDPWR.t174 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X406 a_19190_31850.t31 a_13742_34050.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X407 w_13193_29093.t57 w_13193_29093.t54 w_13193_29093.t56 w_13193_29093.t55 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X408 a_26300_25670.t0 a_26330_25040.t2 VDPWR.t115 VDPWR.t114 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X409 a_26390_32300.t0 a_26420_31750.t2 VDPWR.t85 VDPWR.t84 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X410 a_19190_29050.t32 a_13532_27710.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X411 a_26390_30500.t1 a_26310_26200.t14 VDPWR.t94 VDPWR.t93 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X412 a_25860_21160.t0 V_CONT.t15 w_13193_29093.t196 w_13193_29093.t195 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X413 VDPWR.t26 a_23100_27770.t5 a_23130_27670.t1 VDPWR.t25 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X414 VDPWR.t169 a_14558_34050.t27 a_14140_28370.t2 VDPWR.t168 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X415 a_14348_27710.t44 VDPWR.t372 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X416 a_19190_31610.t6 a_19190_31610.t5 VDPWR.t371 VDPWR.t370 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X417 a_26640_20560.t1 w_13193_29093.t317 VDPWR.t60 VDPWR.t59 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X418 a_23550_31390.t0 a_23100_30570.t5 VDPWR.t179 VDPWR.t178 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X419 a_19190_29050.t33 a_13532_27710.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X420 w_13193_29093.t259 VDPWR.t434 a_18180_28430.t10 w_13193_29093.t258 sky130_fd_pr__nfet_01v8 ad=1.01 pd=6.15 as=1 ps=5.8 w=2.5 l=5
X421 a_14348_27710.t4 a_19190_29050.t34 VDPWR.t415 VDPWR.t414 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X422 VDPWR.t200 a_19190_31850.t32 a_14558_34050.t4 VDPWR.t199 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X423 VDPWR.t246 a_23020_31090.t5 a_23550_31010.t0 VDPWR.t245 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X424 w_13193_29093.t318 V_CONT.t5 sky130_fd_pr__cap_mim_m3_1 l=13.8 w=60
X425 a_19190_31850.t33 a_13742_34050.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X426 w_13193_29093.t53 w_13193_29093.t59 a_13370_29270.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X427 a_14348_27710.t45 VDPWR.t373 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X428 a_19940_23090.t9 a_19940_24230.t8 VDPWR.t240 VDPWR.t239 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X429 a_26390_26970.t3 a_26420_26340.t2 VDPWR.t103 VDPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X430 a_22190_29430.t1 a_14558_34050.t28 VDPWR.t253 VDPWR.t252 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X431 a_24280_30980.t2 a_23100_30460.t5 w_13193_29093.t49 w_13193_29093.t48 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X432 a_13382_33380.t1 a_14990_33260.t0 w_13193_29093.t24 sky130_fd_pr__res_xhigh_po_0p35 l=6
X433 a_14140_28370.t1 a_14558_34050.t29 VDPWR.t139 VDPWR.t138 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X434 a_19190_31850.t34 a_13742_34050.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X435 a_25860_21760.t2 VDPWR.t435 w_13193_29093.t257 w_13193_29093.t140 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X436 a_19040_22530.t0 a_19910_25340.t7 w_13193_29093.t241 w_13193_29093.t4 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X437 a_19190_29050.t35 a_13532_27710.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X438 a_19190_29050.t5 a_19190_29290.t22 VDPWR.t228 VDPWR.t227 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X439 a_14348_27710.t3 a_19190_29050.t36 VDPWR.t389 VDPWR.t388 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X440 V_CONT.t0 a_23130_27670.t7 VDPWR.t196 VDPWR.t195 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X441 VDPWR.t14 a_14348_27710.t46 a_17540_31010.t3 VDPWR.t13 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X442 a_23020_29890.t0 a_23100_30570.t6 w_13193_29093.t201 w_13193_29093.t200 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X443 a_19190_31850.t35 a_13742_34050.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X444 w_13193_29093.t223 a_26390_26310.t12 a_26390_26970.t0 w_13193_29093.t222 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X445 a_17540_31010.t2 a_14348_27710.t47 VDPWR.t16 VDPWR.t15 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X446 w_13193_29093.t236 a_26300_23710.t7 a_26300_24370.t2 w_13193_29093.t235 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X447 VDPWR.t54 a_14348_27710.t48 a_14610_33930.t1 VDPWR.t53 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X448 VDPWR.t5 a_19190_29290.t0 a_19190_29290.t1 VDPWR.t4 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X449 w_13193_29093.t207 a_23020_31090.t6 a_23100_30570.t0 w_13193_29093.t206 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X450 w_13193_29093.t53 w_13193_29093.t52 a_13370_29270.t0 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X451 a_14348_27710.t49 VDPWR.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X452 a_14610_33930.t5 VDPWR.t274 VDPWR.t276 VDPWR.t275 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X453 a_13382_28490.t0 a_14730_30630.t2 w_13193_29093.t131 sky130_fd_pr__res_xhigh_po_0p35 l=6
X454 a_14348_27710.t10 VDPWR.t271 VDPWR.t273 VDPWR.t272 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X455 a_17540_28930.t0 a_17540_28930.t1 w_13193_29093.t3 w_13193_29093.t2 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X456 VDPWR.t270 VDPWR.t268 a_22190_29430.t16 VDPWR.t269 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X457 a_25860_21160.t2 a_26400_21130.t3 a_26400_20530.t0 w_13193_29093.t195 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X458 a_19190_31850.t36 a_13742_34050.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X459 a_26420_30420.t2 a_26320_28790.t11 a_26420_30310.t0 w_13193_29093.t240 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X460 a_19940_23090.t8 a_23130_27960.t3 a_23130_27670.t2 VDPWR.t97 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X461 a_19250_24340.t3 a_19250_24340.t1 a_19250_24340.t2 w_13193_29093.t4 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X462 a_20480_25210.t0 a_18974_25970.t12 VDPWR.t80 VDPWR.t79 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X463 VDPWR.t159 a_19190_31610.t3 a_19190_31610.t4 VDPWR.t158 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
R0 VDPWR.t93 VDPWR.t262 2804.76
R1 VDPWR.t82 VDPWR.t51 2533.33
R2 VDPWR.t384 VDPWR.t21 2307.14
R3 VDPWR.t390 VDPWR.t17 2216.67
R4 VDPWR.t110 VDPWR.t89 2216.67
R5 VDPWR.t70 VDPWR.t73 2216.67
R6 VDPWR.t351 VDPWR.t153 2126.19
R7 VDPWR.t423 VDPWR.t10 1538.1
R8 VDPWR.t12 VDPWR.t193 1492.86
R9 VDPWR.t394 VDPWR.t256 1492.86
R10 VDPWR.t68 VDPWR.t374 1317.78
R11 VDPWR.t84 VDPWR.n22 1289.29
R12 VDPWR.n252 VDPWR.t75 1289.29
R13 VDPWR.t162 VDPWR.t125 1130.95
R14 VDPWR.t34 VDPWR.t260 1130.95
R15 VDPWR.t209 VDPWR.t56 1130.95
R16 VDPWR.t95 VDPWR.t87 1130.95
R17 VDPWR.t417 VDPWR.t61 1130.95
R18 VDPWR.n251 VDPWR.t102 927.381
R19 VDPWR.t114 VDPWR.n106 927.381
R20 VDPWR.n206 VDPWR.t77 927.381
R21 VDPWR.n205 VDPWR.t201 927.381
R22 VDPWR.n949 VDPWR.n300 831.25
R23 VDPWR.n339 VDPWR.n338 831.25
R24 VDPWR.n326 VDPWR.n325 831.25
R25 VDPWR.n332 VDPWR.n331 831.25
R26 VDPWR.n148 VDPWR.n146 831.25
R27 VDPWR.n154 VDPWR.n144 831.25
R28 VDPWR.n867 VDPWR.n866 782
R29 VDPWR.n868 VDPWR.n842 782
R30 VDPWR.n62 VDPWR.t352 733.134
R31 VDPWR.n56 VDPWR.t126 733.134
R32 VDPWR.n575 VDPWR.t286 708.125
R33 VDPWR.t286 VDPWR.n552 708.125
R34 VDPWR.n572 VDPWR.t309 708.125
R35 VDPWR.t309 VDPWR.n553 708.125
R36 VDPWR.n601 VDPWR.t279 708.125
R37 VDPWR.t279 VDPWR.n548 708.125
R38 VDPWR.t339 VDPWR.n549 708.125
R39 VDPWR.n598 VDPWR.t339 708.125
R40 VDPWR.n779 VDPWR.t273 708.125
R41 VDPWR.t273 VDPWR.n772 708.125
R42 VDPWR.n807 VDPWR.t333 708.125
R43 VDPWR.t333 VDPWR.n791 708.125
R44 VDPWR.n825 VDPWR.t312 708.125
R45 VDPWR.t312 VDPWR.n786 708.125
R46 VDPWR.t336 VDPWR.n773 694.444
R47 VDPWR.n776 VDPWR.t336 694.444
R48 VDPWR.n253 VDPWR.t94 663.801
R49 VDPWR.n21 VDPWR.t259 663.801
R50 VDPWR.n250 VDPWR.t22 663.801
R51 VDPWR.n105 VDPWR.t391 663.801
R52 VDPWR.n207 VDPWR.t111 663.801
R53 VDPWR.n204 VDPWR.t74 663.801
R54 VDPWR.n574 VDPWR.t285 657.76
R55 VDPWR.n600 VDPWR.t278 657.76
R56 VDPWR.n243 VDPWR.n88 654.333
R57 VDPWR.n237 VDPWR.n91 654.333
R58 VDPWR.n97 VDPWR.n96 654.333
R59 VDPWR.n100 VDPWR.n99 654.333
R60 VDPWR.n117 VDPWR.n116 654.333
R61 VDPWR.n125 VDPWR.n124 654.333
R62 VDPWR.n197 VDPWR.n135 654.333
R63 VDPWR.n191 VDPWR.n190 654.333
R64 VDPWR.n77 VDPWR.n28 654.333
R65 VDPWR.n70 VDPWR.n31 654.333
R66 VDPWR.n54 VDPWR.n37 654.333
R67 VDPWR.n47 VDPWR.n40 654.333
R68 VDPWR.n7 VDPWR.n6 654.333
R69 VDPWR.n11 VDPWR.n10 654.333
R70 VDPWR.n265 VDPWR.n15 653.115
R71 VDPWR.n778 VDPWR.t272 640.794
R72 VDPWR.n806 VDPWR.t332 640.794
R73 VDPWR.n824 VDPWR.t311 640.794
R74 VDPWR.n22 VDPWR.t258 610.715
R75 VDPWR.n252 VDPWR.t93 610.715
R76 VDPWR.t21 VDPWR.n251 610.715
R77 VDPWR.n106 VDPWR.t390 610.715
R78 VDPWR.n206 VDPWR.t110 610.715
R79 VDPWR.t73 VDPWR.n205 610.715
R80 VDPWR.n755 VDPWR.n710 587.407
R81 VDPWR.n756 VDPWR.n753 587.407
R82 VDPWR.n743 VDPWR.n742 587.407
R83 VDPWR.n744 VDPWR.n718 587.407
R84 VDPWR.n338 VDPWR.n337 585
R85 VDPWR.n336 VDPWR.n300 585
R86 VDPWR.n331 VDPWR.n330 585
R87 VDPWR.n329 VDPWR.n325 585
R88 VDPWR.n746 VDPWR.n744 585
R89 VDPWR.n743 VDPWR.n720 585
R90 VDPWR.n757 VDPWR.n756 585
R91 VDPWR.n755 VDPWR.n713 585
R92 VDPWR.n869 VDPWR.n868 585
R93 VDPWR.n867 VDPWR.n862 585
R94 VDPWR.n662 VDPWR.n661 585
R95 VDPWR.n639 VDPWR.n637 585
R96 VDPWR.n151 VDPWR.n144 585
R97 VDPWR.n150 VDPWR.n146 585
R98 VDPWR.t335 VDPWR.n777 557.783
R99 VDPWR.t308 VDPWR.n573 540.818
R100 VDPWR.t338 VDPWR.n599 540.818
R101 VDPWR.n160 VDPWR.t435 537.492
R102 VDPWR.n170 VDPWR.t433 537.491
R103 VDPWR.n155 VDPWR.t431 537.491
R104 VDPWR.t321 VDPWR.n805 523.855
R105 VDPWR.t269 VDPWR.n823 523.855
R106 VDPWR.t51 VDPWR.t84 497.62
R107 VDPWR.t193 VDPWR.t82 497.62
R108 VDPWR.t211 VDPWR.t12 497.62
R109 VDPWR.t262 VDPWR.t211 497.62
R110 VDPWR.t75 VDPWR.t423 497.62
R111 VDPWR.t10 VDPWR.t162 497.62
R112 VDPWR.t125 VDPWR.t351 497.62
R113 VDPWR.t153 VDPWR.t394 497.62
R114 VDPWR.t256 VDPWR.t384 497.62
R115 VDPWR.t260 VDPWR.t102 497.62
R116 VDPWR.t17 VDPWR.t34 497.62
R117 VDPWR.t56 VDPWR.t114 497.62
R118 VDPWR.t89 VDPWR.t209 497.62
R119 VDPWR.t77 VDPWR.t95 497.62
R120 VDPWR.t87 VDPWR.t70 497.62
R121 VDPWR.t61 VDPWR.t201 497.62
R122 VDPWR.t374 VDPWR.t417 497.62
R123 VDPWR.t246 VDPWR.n301 465.079
R124 VDPWR.n335 VDPWR.t246 465.079
R125 VDPWR.n327 VDPWR.t350 465.079
R126 VDPWR.t350 VDPWR.n324 465.079
R127 VDPWR.n149 VDPWR.t405 465.079
R128 VDPWR.t405 VDPWR.n143 465.079
R129 VDPWR.n385 VDPWR.t141 464.281
R130 VDPWR.t141 VDPWR.n384 464.281
R131 VDPWR.n401 VDPWR.t128 464.281
R132 VDPWR.t128 VDPWR.n400 464.281
R133 VDPWR.t393 VDPWR.n407 464.281
R134 VDPWR.n408 VDPWR.t393 464.281
R135 VDPWR.t208 VDPWR.n391 464.281
R136 VDPWR.n392 VDPWR.t208 464.281
R137 VDPWR.t119 VDPWR.n318 464.281
R138 VDPWR.n319 VDPWR.t119 464.281
R139 VDPWR.t416 VDPWR.n308 464.281
R140 VDPWR.n309 VDPWR.t416 464.281
R141 VDPWR.n440 VDPWR.t425 464.281
R142 VDPWR.t425 VDPWR.n439 464.281
R143 VDPWR.t224 VDPWR.n432 464.281
R144 VDPWR.n433 VDPWR.t224 464.281
R145 VDPWR.n452 VDPWR.t369 464.281
R146 VDPWR.t369 VDPWR.n451 464.281
R147 VDPWR.t235 VDPWR.n459 464.281
R148 VDPWR.n460 VDPWR.t235 464.281
R149 VDPWR.n163 VDPWR.t123 464.281
R150 VDPWR.n166 VDPWR.t123 464.281
R151 VDPWR.t101 VDPWR.n141 464.281
R152 VDPWR.n173 VDPWR.t101 464.281
R153 VDPWR.n865 VDPWR.t282 432.038
R154 VDPWR.t282 VDPWR.n863 432.038
R155 VDPWR.t367 VDPWR.n487 431.421
R156 VDPWR.n488 VDPWR.t367 431.421
R157 VDPWR.n495 VDPWR.t148 431.421
R158 VDPWR.t148 VDPWR.n494 431.421
R159 VDPWR.n508 VDPWR.t144 431.421
R160 VDPWR.t144 VDPWR.n507 431.421
R161 VDPWR.t33 VDPWR.n521 431.421
R162 VDPWR.n522 VDPWR.t33 431.421
R163 VDPWR.n529 VDPWR.t155 431.421
R164 VDPWR.t155 VDPWR.n528 431.421
R165 VDPWR.t26 VDPWR.n933 431.421
R166 VDPWR.n934 VDPWR.t26 431.421
R167 VDPWR.t301 VDPWR.n855 431.421
R168 VDPWR.n856 VDPWR.t301 431.421
R169 VDPWR.n873 VDPWR.t330 431.421
R170 VDPWR.t330 VDPWR.n848 431.421
R171 VDPWR.n781 VDPWR.t271 422.384
R172 VDPWR.n774 VDPWR.t334 422.384
R173 VDPWR.n809 VDPWR.t331 418.368
R174 VDPWR.n802 VDPWR.t320 418.368
R175 VDPWR.n827 VDPWR.t310 418.368
R176 VDPWR.n820 VDPWR.t268 418.368
R177 VDPWR.n513 VDPWR.t432 415.336
R178 VDPWR.t400 VDPWR.t308 407.144
R179 VDPWR.t180 VDPWR.t400 407.144
R180 VDPWR.t156 VDPWR.t180 407.144
R181 VDPWR.t357 VDPWR.t156 407.144
R182 VDPWR.t355 VDPWR.t357 407.144
R183 VDPWR.t363 VDPWR.t355 407.144
R184 VDPWR.t43 VDPWR.t363 407.144
R185 VDPWR.t229 VDPWR.t43 407.144
R186 VDPWR.t27 VDPWR.t229 407.144
R187 VDPWR.t39 VDPWR.t27 407.144
R188 VDPWR.t41 VDPWR.t39 407.144
R189 VDPWR.t191 VDPWR.t41 407.144
R190 VDPWR.t203 VDPWR.t191 407.144
R191 VDPWR.t158 VDPWR.t203 407.144
R192 VDPWR.t370 VDPWR.t158 407.144
R193 VDPWR.t104 VDPWR.t370 407.144
R194 VDPWR.t221 VDPWR.t104 407.144
R195 VDPWR.t199 VDPWR.t221 407.144
R196 VDPWR.t285 VDPWR.t199 407.144
R197 VDPWR.t388 VDPWR.t338 407.144
R198 VDPWR.t406 VDPWR.t388 407.144
R199 VDPWR.t225 VDPWR.t406 407.144
R200 VDPWR.t4 VDPWR.t225 407.144
R201 VDPWR.t2 VDPWR.t4 407.144
R202 VDPWR.t49 VDPWR.t2 407.144
R203 VDPWR.t398 VDPWR.t49 407.144
R204 VDPWR.t386 VDPWR.t398 407.144
R205 VDPWR.t151 VDPWR.t386 407.144
R206 VDPWR.t205 VDPWR.t151 407.144
R207 VDPWR.t108 VDPWR.t205 407.144
R208 VDPWR.t378 VDPWR.t108 407.144
R209 VDPWR.t414 VDPWR.t378 407.144
R210 VDPWR.t408 VDPWR.t414 407.144
R211 VDPWR.t227 VDPWR.t408 407.144
R212 VDPWR.t106 VDPWR.t227 407.144
R213 VDPWR.t410 VDPWR.t106 407.144
R214 VDPWR.t129 VDPWR.t410 407.144
R215 VDPWR.t278 VDPWR.t129 407.144
R216 VDPWR.n670 VDPWR.t287 384.967
R217 VDPWR.n666 VDPWR.t303 384.967
R218 VDPWR.n649 VDPWR.t316 384.967
R219 VDPWR.n644 VDPWR.t295 384.967
R220 VDPWR.n22 VDPWR.n21 382.8
R221 VDPWR.n253 VDPWR.n252 382.8
R222 VDPWR.n251 VDPWR.n250 382.8
R223 VDPWR.n106 VDPWR.n105 382.8
R224 VDPWR.n207 VDPWR.n206 382.8
R225 VDPWR.n205 VDPWR.n204 382.8
R226 VDPWR.n661 VDPWR.t323 374.878
R227 VDPWR.t72 VDPWR.t335 373.214
R228 VDPWR.t236 VDPWR.t72 373.214
R229 VDPWR.t272 VDPWR.t236 373.214
R230 VDPWR.t348 VDPWR.t321 373.214
R231 VDPWR.t166 VDPWR.t348 373.214
R232 VDPWR.t142 VDPWR.t166 373.214
R233 VDPWR.t168 VDPWR.t142 373.214
R234 VDPWR.t164 VDPWR.t168 373.214
R235 VDPWR.t219 VDPWR.t164 373.214
R236 VDPWR.t346 VDPWR.t219 373.214
R237 VDPWR.t266 VDPWR.t346 373.214
R238 VDPWR.t138 VDPWR.t266 373.214
R239 VDPWR.t170 VDPWR.t138 373.214
R240 VDPWR.t332 VDPWR.t170 373.214
R241 VDPWR.t217 VDPWR.t269 373.214
R242 VDPWR.t243 VDPWR.t217 373.214
R243 VDPWR.t344 VDPWR.t243 373.214
R244 VDPWR.t254 VDPWR.t344 373.214
R245 VDPWR.t264 VDPWR.t254 373.214
R246 VDPWR.t241 VDPWR.t264 373.214
R247 VDPWR.t252 VDPWR.t241 373.214
R248 VDPWR.t426 VDPWR.t252 373.214
R249 VDPWR.t353 VDPWR.t426 373.214
R250 VDPWR.t172 VDPWR.t353 373.214
R251 VDPWR.t311 VDPWR.t172 373.214
R252 VDPWR.n577 VDPWR.t284 370.168
R253 VDPWR.n570 VDPWR.t307 370.168
R254 VDPWR.n603 VDPWR.t277 370.168
R255 VDPWR.n596 VDPWR.t337 370.168
R256 VDPWR.n769 VDPWR.t274 360.868
R257 VDPWR.n735 VDPWR.t313 360.868
R258 VDPWR.t412 VDPWR.t300 360.346
R259 VDPWR.t361 VDPWR.t412 360.346
R260 VDPWR.t237 VDPWR.t361 360.346
R261 VDPWR.t0 VDPWR.t237 360.346
R262 VDPWR.t341 VDPWR.t0 360.346
R263 VDPWR.t359 VDPWR.t281 360.346
R264 VDPWR.t6 VDPWR.t359 360.346
R265 VDPWR.t23 VDPWR.t6 360.346
R266 VDPWR.t195 VDPWR.t23 360.346
R267 VDPWR.t328 VDPWR.t195 360.346
R268 VDPWR.n160 VDPWR.t69 359.752
R269 VDPWR.n170 VDPWR.t67 359.752
R270 VDPWR.n155 VDPWR.t60 359.752
R271 VDPWR.n638 VDPWR.t291 352.834
R272 VDPWR.n793 VDPWR.t322 351.793
R273 VDPWR.n788 VDPWR.t270 351.793
R274 VDPWR.t300 VDPWR.n859 343.966
R275 VDPWR.n872 VDPWR.t341 343.966
R276 VDPWR.t281 VDPWR.n872 343.966
R277 VDPWR.n878 VDPWR.t328 343.966
R278 VDPWR.n645 VDPWR.t297 341.752
R279 VDPWR.n650 VDPWR.t319 341.752
R280 VDPWR.n667 VDPWR.t305 341.752
R281 VDPWR.n669 VDPWR.t290 341.75
R282 VDPWR.n864 VDPWR.t340 336.329
R283 VDPWR.n864 VDPWR.t280 336.329
R284 VDPWR.n624 VDPWR.n623 322.046
R285 VDPWR.n672 VDPWR.n625 322.046
R286 VDPWR.n620 VDPWR.n619 322.046
R287 VDPWR.n648 VDPWR.n647 322.046
R288 VDPWR.n643 VDPWR.n642 322.046
R289 VDPWR.n671 VDPWR.n626 322.046
R290 VDPWR.n410 VDPWR.t397 321.649
R291 VDPWR.n831 VDPWR.t299 320.7
R292 VDPWR.n881 VDPWR.t327 320.7
R293 VDPWR.n669 VDPWR.t288 315.325
R294 VDPWR.t124 VDPWR.t174 314.113
R295 VDPWR.t216 VDPWR.t86 314.113
R296 VDPWR.n801 VDPWR.n800 301.933
R297 VDPWR.n799 VDPWR.n798 301.933
R298 VDPWR.n797 VDPWR.n796 301.933
R299 VDPWR.n795 VDPWR.n794 301.933
R300 VDPWR.n790 VDPWR.n789 301.933
R301 VDPWR.n818 VDPWR.n817 301.933
R302 VDPWR.n816 VDPWR.n815 301.933
R303 VDPWR.n814 VDPWR.n813 301.933
R304 VDPWR.n812 VDPWR.n811 301.933
R305 VDPWR.n785 VDPWR.n784 301.933
R306 VDPWR.n569 VDPWR.n568 299.231
R307 VDPWR.n567 VDPWR.n566 299.231
R308 VDPWR.n565 VDPWR.n564 299.231
R309 VDPWR.n563 VDPWR.n562 299.231
R310 VDPWR.n561 VDPWR.n560 299.231
R311 VDPWR.n559 VDPWR.n558 299.231
R312 VDPWR.n557 VDPWR.n556 299.231
R313 VDPWR.n555 VDPWR.n554 299.231
R314 VDPWR.n551 VDPWR.n550 299.231
R315 VDPWR.n594 VDPWR.n593 299.231
R316 VDPWR.n592 VDPWR.n591 299.231
R317 VDPWR.n590 VDPWR.n589 299.231
R318 VDPWR.n588 VDPWR.n587 299.231
R319 VDPWR.n586 VDPWR.n585 299.231
R320 VDPWR.n584 VDPWR.n583 299.231
R321 VDPWR.n582 VDPWR.n581 299.231
R322 VDPWR.n580 VDPWR.n579 299.231
R323 VDPWR.n547 VDPWR.n546 299.231
R324 VDPWR.n662 VDPWR.n656 290.733
R325 VDPWR.n663 VDPWR.n662 290.733
R326 VDPWR.n637 VDPWR.n636 290.733
R327 VDPWR.n637 VDPWR.n631 290.733
R328 VDPWR.t189 VDPWR.t314 251.471
R329 VDPWR.t231 VDPWR.t189 251.471
R330 VDPWR.t186 VDPWR.t231 251.471
R331 VDPWR.t36 VDPWR.t186 251.471
R332 VDPWR.t380 VDPWR.t36 251.471
R333 VDPWR.t382 VDPWR.t380 251.471
R334 VDPWR.t63 VDPWR.t382 251.471
R335 VDPWR.t29 VDPWR.t63 251.471
R336 VDPWR.t183 VDPWR.t29 251.471
R337 VDPWR.t419 VDPWR.t183 251.471
R338 VDPWR.t421 VDPWR.t419 251.471
R339 VDPWR.t213 VDPWR.t421 251.471
R340 VDPWR.t132 VDPWR.t213 251.471
R341 VDPWR.t13 VDPWR.t132 251.471
R342 VDPWR.t15 VDPWR.t13 251.471
R343 VDPWR.t53 VDPWR.t15 251.471
R344 VDPWR.t275 VDPWR.t53 251.471
R345 VDPWR.n320 VDPWR.n319 243.698
R346 VDPWR.n439 VDPWR.n344 243.698
R347 VDPWR.n451 VDPWR.n346 243.698
R348 VDPWR.n400 VDPWR.n350 243.698
R349 VDPWR.n384 VDPWR.n354 243.698
R350 VDPWR.n407 VDPWR.n351 243.698
R351 VDPWR.n391 VDPWR.n355 243.698
R352 VDPWR.n308 VDPWR.n303 243.698
R353 VDPWR.n432 VDPWR.n341 243.698
R354 VDPWR.n459 VDPWR.n347 243.698
R355 VDPWR.n311 VDPWR.n310 238.367
R356 VDPWR.n340 VDPWR.n339 238.367
R357 VDPWR.n333 VDPWR.n332 238.367
R358 VDPWR.n434 VDPWR.n342 238.367
R359 VDPWR.n461 VDPWR.n348 238.367
R360 VDPWR.n409 VDPWR.n352 238.367
R361 VDPWR.n393 VDPWR.n356 238.367
R362 VDPWR.n386 VDPWR.n353 238.367
R363 VDPWR.n402 VDPWR.n349 238.367
R364 VDPWR.n453 VDPWR.n345 238.367
R365 VDPWR.n441 VDPWR.n343 238.367
R366 VDPWR.n326 VDPWR.n322 238.367
R367 VDPWR.n949 VDPWR.n948 238.367
R368 VDPWR.n315 VDPWR.n312 238.367
R369 VDPWR.n573 VDPWR.n572 238.367
R370 VDPWR.n573 VDPWR.n553 238.367
R371 VDPWR.n599 VDPWR.n598 238.367
R372 VDPWR.n599 VDPWR.n549 238.367
R373 VDPWR.n750 VDPWR.n749 238.367
R374 VDPWR.n736 VDPWR.n715 238.367
R375 VDPWR.n768 VDPWR.n711 238.367
R376 VDPWR.n761 VDPWR.n760 238.367
R377 VDPWR.n777 VDPWR.n776 238.367
R378 VDPWR.n777 VDPWR.n773 238.367
R379 VDPWR.n805 VDPWR.n804 238.367
R380 VDPWR.n805 VDPWR.n792 238.367
R381 VDPWR.n823 VDPWR.n822 238.367
R382 VDPWR.n823 VDPWR.n787 238.367
R383 VDPWR.n168 VDPWR.n167 238.367
R384 VDPWR.n172 VDPWR.n171 238.367
R385 VDPWR.n154 VDPWR.n153 238.367
R386 VDPWR.n148 VDPWR.n147 238.367
R387 VDPWR.n178 VDPWR.n177 238.367
R388 VDPWR.n162 VDPWR.n158 238.367
R389 VDPWR.t314 VDPWR.n751 237.5
R390 VDPWR.n762 VDPWR.t275 237.5
R391 VDPWR.n494 VDPWR.n360 234.355
R392 VDPWR.n487 VDPWR.n357 234.355
R393 VDPWR.n507 VDPWR.n362 234.355
R394 VDPWR.n528 VDPWR.n366 234.355
R395 VDPWR.n521 VDPWR.n363 234.355
R396 VDPWR.n935 VDPWR.n934 234.355
R397 VDPWR.n855 VDPWR.n850 234.355
R398 VDPWR.n877 VDPWR.n873 234.355
R399 VDPWR.n631 VDPWR.n627 233.841
R400 VDPWR.n489 VDPWR.n358 230.308
R401 VDPWR.n523 VDPWR.n364 230.308
R402 VDPWR.n530 VDPWR.n365 230.308
R403 VDPWR.n509 VDPWR.n361 230.308
R404 VDPWR.n496 VDPWR.n359 230.308
R405 VDPWR.n930 VDPWR.n367 230.308
R406 VDPWR.n858 VDPWR.n857 230.308
R407 VDPWR.n880 VDPWR.n879 230.308
R408 VDPWR.n866 VDPWR.n860 230.308
R409 VDPWR.n871 VDPWR.n842 230.308
R410 VDPWR.n661 VDPWR.n652 230.308
R411 VDPWR.t32 VDPWR.t97 222.178
R412 VDPWR.n169 VDPWR.t122 219.232
R413 VDPWR.t100 VDPWR.n156 219.232
R414 VDPWR.t98 VDPWR.n142 219.232
R415 VDPWR.n142 VDPWR.t404 219.232
R416 VDPWR.n940 VDPWR.n939 199.195
R417 VDPWR.n884 VDPWR.n883 196.502
R418 VDPWR.n892 VDPWR.n891 196.502
R419 VDPWR.n900 VDPWR.n899 196.502
R420 VDPWR.n839 VDPWR.n838 196.502
R421 VDPWR.n917 VDPWR.n836 196.502
R422 VDPWR.n923 VDPWR.n833 196.502
R423 VDPWR.n664 VDPWR.n663 188.536
R424 VDPWR.n170 VDPWR.t100 185.002
R425 VDPWR.t98 VDPWR.n155 185.002
R426 VDPWR.n160 VDPWR.t122 185.002
R427 VDPWR.n668 VDPWR.n667 185.001
R428 VDPWR.n651 VDPWR.n650 185.001
R429 VDPWR.n646 VDPWR.n645 185.001
R430 VDPWR.n518 VDPWR.n517 185
R431 VDPWR.n520 VDPWR.n519 185
R432 VDPWR.n527 VDPWR.n526 185
R433 VDPWR.n525 VDPWR.n524 185
R434 VDPWR.n506 VDPWR.n505 185
R435 VDPWR.n504 VDPWR.n503 185
R436 VDPWR.n484 VDPWR.n483 185
R437 VDPWR.n486 VDPWR.n485 185
R438 VDPWR.n493 VDPWR.n492 185
R439 VDPWR.n491 VDPWR.n490 185
R440 VDPWR.n388 VDPWR.n387 185
R441 VDPWR.n390 VDPWR.n389 185
R442 VDPWR.n383 VDPWR.n382 185
R443 VDPWR.n381 VDPWR.n380 185
R444 VDPWR.n404 VDPWR.n403 185
R445 VDPWR.n406 VDPWR.n405 185
R446 VDPWR.n399 VDPWR.n398 185
R447 VDPWR.n397 VDPWR.n396 185
R448 VDPWR.n456 VDPWR.n455 185
R449 VDPWR.n458 VDPWR.n457 185
R450 VDPWR.n450 VDPWR.n449 185
R451 VDPWR.n448 VDPWR.n447 185
R452 VDPWR.n429 VDPWR.n428 185
R453 VDPWR.n431 VDPWR.n430 185
R454 VDPWR.n438 VDPWR.n437 185
R455 VDPWR.n436 VDPWR.n435 185
R456 VDPWR.n330 VDPWR.n323 185
R457 VDPWR.n329 VDPWR.n328 185
R458 VDPWR.n337 VDPWR.n334 185
R459 VDPWR.n336 VDPWR.n302 185
R460 VDPWR.n305 VDPWR.n304 185
R461 VDPWR.n307 VDPWR.n306 185
R462 VDPWR.n314 VDPWR.n313 185
R463 VDPWR.n317 VDPWR.n316 185
R464 VDPWR.n369 VDPWR.n368 185
R465 VDPWR.n932 VDPWR.n931 185
R466 VDPWR.n747 VDPWR.n717 185
R467 VDPWR.n746 VDPWR.n745 185
R468 VDPWR.n739 VDPWR.n720 185
R469 VDPWR.n741 VDPWR.n740 185
R470 VDPWR.n758 VDPWR.n752 185
R471 VDPWR.n757 VDPWR.n714 185
R472 VDPWR.n764 VDPWR.n713 185
R473 VDPWR.n766 VDPWR.n765 185
R474 VDPWR.n874 VDPWR.n849 185
R475 VDPWR.n876 VDPWR.n875 185
R476 VDPWR.n852 VDPWR.n851 185
R477 VDPWR.n854 VDPWR.n853 185
R478 VDPWR.n870 VDPWR.n869 185
R479 VDPWR.n862 VDPWR.n861 185
R480 VDPWR.n660 VDPWR.n659 185
R481 VDPWR.n658 VDPWR.n657 185
R482 VDPWR.n655 VDPWR.n654 185
R483 VDPWR.n665 VDPWR.n664 185
R484 VDPWR.n640 VDPWR.n639 185
R485 VDPWR.n641 VDPWR.n640 185
R486 VDPWR.n630 VDPWR.n629 185
R487 VDPWR.n635 VDPWR.n634 185
R488 VDPWR.n633 VDPWR.n632 185
R489 VDPWR.n152 VDPWR.n151 185
R490 VDPWR.n150 VDPWR.n145 185
R491 VDPWR.n174 VDPWR.n157 185
R492 VDPWR.n176 VDPWR.n175 185
R493 VDPWR.n165 VDPWR.n159 185
R494 VDPWR.n164 VDPWR.n161 185
R495 VDPWR.t147 VDPWR.n938 172.38
R496 VDPWR.t58 VDPWR.n937 172.38
R497 VDPWR.t97 VDPWR.n936 172.38
R498 VDPWR.n866 VDPWR.n864 166.63
R499 VDPWR.t66 VDPWR.n169 158.333
R500 VDPWR.n156 VDPWR.t59 158.333
R501 VDPWR.n316 VDPWR.n313 150
R502 VDPWR.n306 VDPWR.n304 150
R503 VDPWR.n334 VDPWR.n302 150
R504 VDPWR.n328 VDPWR.n323 150
R505 VDPWR.n437 VDPWR.n436 150
R506 VDPWR.n430 VDPWR.n429 150
R507 VDPWR.n449 VDPWR.n448 150
R508 VDPWR.n457 VDPWR.n456 150
R509 VDPWR.n398 VDPWR.n397 150
R510 VDPWR.n405 VDPWR.n404 150
R511 VDPWR.n382 VDPWR.n381 150
R512 VDPWR.n389 VDPWR.n388 150
R513 VDPWR.n740 VDPWR.n739 150
R514 VDPWR.n745 VDPWR.n717 150
R515 VDPWR.n765 VDPWR.n764 150
R516 VDPWR.n752 VDPWR.n714 150
R517 VDPWR.n161 VDPWR.n159 150
R518 VDPWR.n176 VDPWR.n157 150
R519 VDPWR.n152 VDPWR.n145 150
R520 VDPWR.t160 VDPWR.t145 145.038
R521 VDPWR.n734 VDPWR.n733 141.709
R522 VDPWR.n732 VDPWR.n731 141.709
R523 VDPWR.n730 VDPWR.n729 141.709
R524 VDPWR.n728 VDPWR.n727 141.709
R525 VDPWR.n726 VDPWR.n725 141.709
R526 VDPWR.n724 VDPWR.n723 141.709
R527 VDPWR.n722 VDPWR.n721 141.709
R528 VDPWR.n709 VDPWR.n708 141.709
R529 VDPWR.n944 VDPWR.n943 137.904
R530 VDPWR.n942 VDPWR.n941 137.904
R531 VDPWR.n939 VDPWR.t147 126.412
R532 VDPWR.n938 VDPWR.t58 126.412
R533 VDPWR.n937 VDPWR.t32 126.412
R534 VDPWR.n936 VDPWR.t25 126.412
R535 VDPWR.t179 VDPWR.n300 123.126
R536 VDPWR.n338 VDPWR.t179 123.126
R537 VDPWR.n325 VDPWR.t248 123.126
R538 VDPWR.n331 VDPWR.t248 123.126
R539 VDPWR.t276 VDPWR.n755 123.126
R540 VDPWR.n756 VDPWR.t276 123.126
R541 VDPWR.t315 VDPWR.n743 123.126
R542 VDPWR.n744 VDPWR.t315 123.126
R543 VDPWR.n146 VDPWR.t99 123.126
R544 VDPWR.t99 VDPWR.n144 123.126
R545 VDPWR.n492 VDPWR.n491 120.001
R546 VDPWR.n485 VDPWR.n484 120.001
R547 VDPWR.n505 VDPWR.n504 120.001
R548 VDPWR.n526 VDPWR.n525 120.001
R549 VDPWR.n519 VDPWR.n518 120.001
R550 VDPWR.n931 VDPWR.n368 120.001
R551 VDPWR.n853 VDPWR.n851 120.001
R552 VDPWR.n876 VDPWR.n849 120.001
R553 VDPWR.n870 VDPWR.n861 120.001
R554 VDPWR.n664 VDPWR.n654 120.001
R555 VDPWR.n659 VDPWR.n658 120.001
R556 VDPWR.n634 VDPWR.n633 120.001
R557 VDPWR.n640 VDPWR.n629 120.001
R558 VDPWR.n702 VDPWR.n608 119.737
R559 VDPWR.n695 VDPWR.n611 119.737
R560 VDPWR.n688 VDPWR.n614 119.737
R561 VDPWR.n681 VDPWR.n617 119.737
R562 VDPWR.n674 VDPWR.n622 119.737
R563 VDPWR.t304 VDPWR.n668 119.656
R564 VDPWR.t122 VDPWR.t68 109.615
R565 VDPWR.t100 VDPWR.t66 109.615
R566 VDPWR.t59 VDPWR.t98 109.615
R567 VDPWR.n665 VDPWR.n651 108.779
R568 VDPWR.n946 VDPWR.n945 107.258
R569 VDPWR.t118 VDPWR.n321 103.427
R570 VDPWR.n947 VDPWR.t178 103.427
R571 VDPWR.n947 VDPWR.t245 103.427
R572 VDPWR.t223 VDPWR.n946 103.427
R573 VDPWR.t343 VDPWR.n867 98.5005
R574 VDPWR.n868 VDPWR.t343 98.5005
R575 VDPWR.n945 VDPWR.t234 95.7666
R576 VDPWR.t81 VDPWR.t250 94.2753
R577 VDPWR.t249 VDPWR.t177 94.2753
R578 VDPWR.t402 VDPWR.n646 94.2753
R579 VDPWR.t91 VDPWR.t296 94.2753
R580 VDPWR.t136 VDPWR.t175 94.2753
R581 VDPWR.t112 VDPWR.t304 94.2753
R582 VDPWR.t239 VDPWR.t112 94.2753
R583 VDPWR.t197 VDPWR.t239 94.2753
R584 VDPWR.t8 VDPWR.t197 94.2753
R585 VDPWR.t288 VDPWR.t8 94.2753
R586 VDPWR.t392 VDPWR.t127 91.936
R587 VDPWR.t207 VDPWR.t140 91.936
R588 VDPWR.n155 VDPWR.n154 90.5056
R589 VDPWR.t174 VDPWR.t118 84.2747
R590 VDPWR.t178 VDPWR.t124 84.2747
R591 VDPWR.t245 VDPWR.t216 84.2747
R592 VDPWR.t86 VDPWR.t223 84.2747
R593 VDPWR.t368 VDPWR.t396 84.2747
R594 VDPWR.t79 VDPWR.t251 83.3974
R595 VDPWR.t324 VDPWR.t317 83.3974
R596 VDPWR.n88 VDPWR.t103 78.8005
R597 VDPWR.n88 VDPWR.t261 78.8005
R598 VDPWR.n91 VDPWR.t35 78.8005
R599 VDPWR.n91 VDPWR.t18 78.8005
R600 VDPWR.n96 VDPWR.t115 78.8005
R601 VDPWR.n96 VDPWR.t57 78.8005
R602 VDPWR.n99 VDPWR.t210 78.8005
R603 VDPWR.n99 VDPWR.t90 78.8005
R604 VDPWR.n116 VDPWR.t78 78.8005
R605 VDPWR.n116 VDPWR.t96 78.8005
R606 VDPWR.n124 VDPWR.t88 78.8005
R607 VDPWR.n124 VDPWR.t71 78.8005
R608 VDPWR.n135 VDPWR.t202 78.8005
R609 VDPWR.n135 VDPWR.t62 78.8005
R610 VDPWR.n190 VDPWR.t418 78.8005
R611 VDPWR.n190 VDPWR.t375 78.8005
R612 VDPWR.n28 VDPWR.t257 78.8005
R613 VDPWR.n28 VDPWR.t385 78.8005
R614 VDPWR.n31 VDPWR.t154 78.8005
R615 VDPWR.n31 VDPWR.t395 78.8005
R616 VDPWR.n37 VDPWR.t11 78.8005
R617 VDPWR.n37 VDPWR.t163 78.8005
R618 VDPWR.n40 VDPWR.t76 78.8005
R619 VDPWR.n40 VDPWR.t424 78.8005
R620 VDPWR.n6 VDPWR.t85 78.8005
R621 VDPWR.n6 VDPWR.t52 78.8005
R622 VDPWR.n10 VDPWR.t83 78.8005
R623 VDPWR.n10 VDPWR.t194 78.8005
R624 VDPWR.n15 VDPWR.t212 78.8005
R625 VDPWR.n15 VDPWR.t263 78.8005
R626 VDPWR.t292 VDPWR.t247 76.1455
R627 VDPWR.t365 VDPWR.t19 76.1455
R628 VDPWR.n673 VDPWR.n672 75.7203
R629 VDPWR.n172 VDPWR.n170 74.7688
R630 VDPWR.n167 VDPWR.n160 74.7688
R631 VDPWR.n672 VDPWR.n624 70.4005
R632 VDPWR.n643 VDPWR.n620 70.4005
R633 VDPWR.n648 VDPWR.n620 70.4005
R634 VDPWR.n672 VDPWR.n671 70.4005
R635 VDPWR.n937 VDPWR.n364 69.8479
R636 VDPWR.n937 VDPWR.n363 69.8479
R637 VDPWR.n937 VDPWR.n366 69.8479
R638 VDPWR.n937 VDPWR.n365 69.8479
R639 VDPWR.n938 VDPWR.n362 69.8479
R640 VDPWR.n938 VDPWR.n361 69.8479
R641 VDPWR.n939 VDPWR.n358 69.8479
R642 VDPWR.n939 VDPWR.n357 69.8479
R643 VDPWR.n939 VDPWR.n360 69.8479
R644 VDPWR.n939 VDPWR.n359 69.8479
R645 VDPWR.n936 VDPWR.n935 69.8479
R646 VDPWR.n936 VDPWR.n367 69.8479
R647 VDPWR.n879 VDPWR.n878 69.8479
R648 VDPWR.n878 VDPWR.n877 69.8479
R649 VDPWR.n859 VDPWR.n858 69.8479
R650 VDPWR.n859 VDPWR.n850 69.8479
R651 VDPWR.n872 VDPWR.n871 69.8479
R652 VDPWR.n872 VDPWR.n860 69.8479
R653 VDPWR.n665 VDPWR.n652 69.8479
R654 VDPWR.n665 VDPWR.n653 69.8479
R655 VDPWR.n641 VDPWR.n628 69.8479
R656 VDPWR.n641 VDPWR.n627 69.8479
R657 VDPWR.t247 VDPWR.n641 68.8936
R658 VDPWR.t19 VDPWR.t149 68.8936
R659 VDPWR.n940 VDPWR.n356 65.8183
R660 VDPWR.n940 VDPWR.n355 65.8183
R661 VDPWR.n941 VDPWR.n354 65.8183
R662 VDPWR.n941 VDPWR.n353 65.8183
R663 VDPWR.n942 VDPWR.n352 65.8183
R664 VDPWR.n942 VDPWR.n351 65.8183
R665 VDPWR.n943 VDPWR.n350 65.8183
R666 VDPWR.n943 VDPWR.n349 65.8183
R667 VDPWR.n944 VDPWR.n348 65.8183
R668 VDPWR.n944 VDPWR.n347 65.8183
R669 VDPWR.n945 VDPWR.n346 65.8183
R670 VDPWR.n945 VDPWR.n345 65.8183
R671 VDPWR.n946 VDPWR.n342 65.8183
R672 VDPWR.n946 VDPWR.n341 65.8183
R673 VDPWR.n946 VDPWR.n344 65.8183
R674 VDPWR.n946 VDPWR.n343 65.8183
R675 VDPWR.n947 VDPWR.n333 65.8183
R676 VDPWR.n947 VDPWR.n322 65.8183
R677 VDPWR.n947 VDPWR.n340 65.8183
R678 VDPWR.n948 VDPWR.n947 65.8183
R679 VDPWR.n321 VDPWR.n311 65.8183
R680 VDPWR.n321 VDPWR.n303 65.8183
R681 VDPWR.n321 VDPWR.n320 65.8183
R682 VDPWR.n321 VDPWR.n312 65.8183
R683 VDPWR.n751 VDPWR.n750 65.8183
R684 VDPWR.n751 VDPWR.n716 65.8183
R685 VDPWR.n751 VDPWR.n715 65.8183
R686 VDPWR.n762 VDPWR.n761 65.8183
R687 VDPWR.n763 VDPWR.n762 65.8183
R688 VDPWR.n762 VDPWR.n711 65.8183
R689 VDPWR.n153 VDPWR.n142 65.8183
R690 VDPWR.n147 VDPWR.n142 65.8183
R691 VDPWR.n171 VDPWR.n156 65.8183
R692 VDPWR.n177 VDPWR.n156 65.8183
R693 VDPWR.n169 VDPWR.n168 65.8183
R694 VDPWR.n169 VDPWR.n158 65.8183
R695 VDPWR.n315 VDPWR.n292 64.4576
R696 VDPWR.n310 VDPWR.n292 64.4576
R697 VDPWR.n442 VDPWR.n441 64.4576
R698 VDPWR.n442 VDPWR.n434 64.4576
R699 VDPWR.n454 VDPWR.n453 64.4576
R700 VDPWR.n462 VDPWR.n461 64.4576
R701 VDPWR.n497 VDPWR.n496 63.6449
R702 VDPWR.n497 VDPWR.n489 63.6449
R703 VDPWR.n510 VDPWR.n509 63.6449
R704 VDPWR.n531 VDPWR.n530 63.6449
R705 VDPWR.n531 VDPWR.n523 63.6449
R706 VDPWR.n930 VDPWR.n929 63.6449
R707 VDPWR.t251 VDPWR.t45 61.6417
R708 VDPWR.t317 VDPWR.t47 61.6417
R709 VDPWR.n951 VDPWR.n298 60.8005
R710 VDPWR.n951 VDPWR.n950 60.8005
R711 VDPWR.n299 VDPWR.n298 60.8005
R712 VDPWR.n950 VDPWR.n299 60.8005
R713 VDPWR.n21 VDPWR.n2 60.8005
R714 VDPWR.n254 VDPWR.n253 60.8005
R715 VDPWR.n250 VDPWR.n249 60.8005
R716 VDPWR.n105 VDPWR.n94 60.8005
R717 VDPWR.n208 VDPWR.n207 60.8005
R718 VDPWR.n204 VDPWR.n203 60.8005
R719 VDPWR.n542 VDPWR.t429 58.8
R720 VDPWR.n541 VDPWR.t430 58.8
R721 VDPWR.n476 VDPWR.n386 58.0576
R722 VDPWR.n469 VDPWR.n402 58.0576
R723 VDPWR.n468 VDPWR.n409 58.0576
R724 VDPWR.n475 VDPWR.n393 58.0576
R725 VDPWR.n679 VDPWR.n620 54.4005
R726 VDPWR.n316 VDPWR.n312 53.3664
R727 VDPWR.n306 VDPWR.n303 53.3664
R728 VDPWR.n948 VDPWR.n302 53.3664
R729 VDPWR.n328 VDPWR.n322 53.3664
R730 VDPWR.n436 VDPWR.n343 53.3664
R731 VDPWR.n430 VDPWR.n341 53.3664
R732 VDPWR.n448 VDPWR.n345 53.3664
R733 VDPWR.n457 VDPWR.n347 53.3664
R734 VDPWR.n397 VDPWR.n349 53.3664
R735 VDPWR.n405 VDPWR.n351 53.3664
R736 VDPWR.n381 VDPWR.n353 53.3664
R737 VDPWR.n389 VDPWR.n355 53.3664
R738 VDPWR.n388 VDPWR.n356 53.3664
R739 VDPWR.n382 VDPWR.n354 53.3664
R740 VDPWR.n404 VDPWR.n352 53.3664
R741 VDPWR.n398 VDPWR.n350 53.3664
R742 VDPWR.n456 VDPWR.n348 53.3664
R743 VDPWR.n449 VDPWR.n346 53.3664
R744 VDPWR.n429 VDPWR.n342 53.3664
R745 VDPWR.n437 VDPWR.n344 53.3664
R746 VDPWR.n333 VDPWR.n323 53.3664
R747 VDPWR.n340 VDPWR.n334 53.3664
R748 VDPWR.n311 VDPWR.n304 53.3664
R749 VDPWR.n320 VDPWR.n313 53.3664
R750 VDPWR.n740 VDPWR.n715 53.3664
R751 VDPWR.n745 VDPWR.n716 53.3664
R752 VDPWR.n750 VDPWR.n717 53.3664
R753 VDPWR.n739 VDPWR.n716 53.3664
R754 VDPWR.n764 VDPWR.n763 53.3664
R755 VDPWR.n761 VDPWR.n752 53.3664
R756 VDPWR.n763 VDPWR.n714 53.3664
R757 VDPWR.n765 VDPWR.n711 53.3664
R758 VDPWR.n161 VDPWR.n158 53.3664
R759 VDPWR.n177 VDPWR.n176 53.3664
R760 VDPWR.n147 VDPWR.n145 53.3664
R761 VDPWR.n153 VDPWR.n152 53.3664
R762 VDPWR.n171 VDPWR.n157 53.3664
R763 VDPWR.n168 VDPWR.n159 53.3664
R764 VDPWR.n646 VDPWR.t160 50.7639
R765 VDPWR.n623 VDPWR.t306 49.2505
R766 VDPWR.n623 VDPWR.t113 49.2505
R767 VDPWR.n625 VDPWR.t240 49.2505
R768 VDPWR.n625 VDPWR.t198 49.2505
R769 VDPWR.n619 VDPWR.t20 49.2505
R770 VDPWR.n619 VDPWR.t176 49.2505
R771 VDPWR.n647 VDPWR.t137 49.2505
R772 VDPWR.n647 VDPWR.t318 49.2505
R773 VDPWR.n642 VDPWR.t298 49.2505
R774 VDPWR.n642 VDPWR.t92 49.2505
R775 VDPWR.n626 VDPWR.t9 49.2505
R776 VDPWR.n626 VDPWR.t289 49.2505
R777 VDPWR.n541 VDPWR.t428 49.164
R778 VDPWR.n543 VDPWR.t434 48.5159
R779 VDPWR.n670 VDPWR.n669 46.218
R780 VDPWR.n491 VDPWR.n359 45.3071
R781 VDPWR.n485 VDPWR.n357 45.3071
R782 VDPWR.n504 VDPWR.n361 45.3071
R783 VDPWR.n525 VDPWR.n365 45.3071
R784 VDPWR.n519 VDPWR.n363 45.3071
R785 VDPWR.n518 VDPWR.n364 45.3071
R786 VDPWR.n526 VDPWR.n366 45.3071
R787 VDPWR.n505 VDPWR.n362 45.3071
R788 VDPWR.n484 VDPWR.n358 45.3071
R789 VDPWR.n492 VDPWR.n360 45.3071
R790 VDPWR.n935 VDPWR.n368 45.3071
R791 VDPWR.n931 VDPWR.n367 45.3071
R792 VDPWR.n853 VDPWR.n850 45.3071
R793 VDPWR.n877 VDPWR.n876 45.3071
R794 VDPWR.n879 VDPWR.n849 45.3071
R795 VDPWR.n858 VDPWR.n851 45.3071
R796 VDPWR.n871 VDPWR.n870 45.3071
R797 VDPWR.n861 VDPWR.n860 45.3071
R798 VDPWR.n658 VDPWR.n653 45.3071
R799 VDPWR.n659 VDPWR.n652 45.3071
R800 VDPWR.n654 VDPWR.n653 45.3071
R801 VDPWR.n634 VDPWR.n628 45.3071
R802 VDPWR.n629 VDPWR.n628 45.3071
R803 VDPWR.n633 VDPWR.n627 45.3071
R804 VDPWR.t145 VDPWR.t249 39.886
R805 VDPWR.n706 VDPWR.n705 39.4993
R806 VDPWR.n673 VDPWR.n621 39.4988
R807 VDPWR.n568 VDPWR.t401 39.4005
R808 VDPWR.n568 VDPWR.t181 39.4005
R809 VDPWR.n566 VDPWR.t157 39.4005
R810 VDPWR.n566 VDPWR.t358 39.4005
R811 VDPWR.n564 VDPWR.t356 39.4005
R812 VDPWR.n564 VDPWR.t364 39.4005
R813 VDPWR.n562 VDPWR.t44 39.4005
R814 VDPWR.n562 VDPWR.t230 39.4005
R815 VDPWR.n560 VDPWR.t28 39.4005
R816 VDPWR.n560 VDPWR.t40 39.4005
R817 VDPWR.n558 VDPWR.t42 39.4005
R818 VDPWR.n558 VDPWR.t192 39.4005
R819 VDPWR.n556 VDPWR.t204 39.4005
R820 VDPWR.n556 VDPWR.t159 39.4005
R821 VDPWR.n554 VDPWR.t371 39.4005
R822 VDPWR.n554 VDPWR.t105 39.4005
R823 VDPWR.n550 VDPWR.t222 39.4005
R824 VDPWR.n550 VDPWR.t200 39.4005
R825 VDPWR.n593 VDPWR.t389 39.4005
R826 VDPWR.n593 VDPWR.t407 39.4005
R827 VDPWR.n591 VDPWR.t226 39.4005
R828 VDPWR.n591 VDPWR.t5 39.4005
R829 VDPWR.n589 VDPWR.t3 39.4005
R830 VDPWR.n589 VDPWR.t50 39.4005
R831 VDPWR.n587 VDPWR.t399 39.4005
R832 VDPWR.n587 VDPWR.t387 39.4005
R833 VDPWR.n585 VDPWR.t152 39.4005
R834 VDPWR.n585 VDPWR.t206 39.4005
R835 VDPWR.n583 VDPWR.t109 39.4005
R836 VDPWR.n583 VDPWR.t379 39.4005
R837 VDPWR.n581 VDPWR.t415 39.4005
R838 VDPWR.n581 VDPWR.t409 39.4005
R839 VDPWR.n579 VDPWR.t228 39.4005
R840 VDPWR.n579 VDPWR.t107 39.4005
R841 VDPWR.n546 VDPWR.t411 39.4005
R842 VDPWR.n546 VDPWR.t130 39.4005
R843 VDPWR.n800 VDPWR.t349 39.4005
R844 VDPWR.n800 VDPWR.t167 39.4005
R845 VDPWR.n798 VDPWR.t143 39.4005
R846 VDPWR.n798 VDPWR.t169 39.4005
R847 VDPWR.n796 VDPWR.t165 39.4005
R848 VDPWR.n796 VDPWR.t220 39.4005
R849 VDPWR.n794 VDPWR.t347 39.4005
R850 VDPWR.n794 VDPWR.t267 39.4005
R851 VDPWR.n789 VDPWR.t139 39.4005
R852 VDPWR.n789 VDPWR.t171 39.4005
R853 VDPWR.n817 VDPWR.t218 39.4005
R854 VDPWR.n817 VDPWR.t244 39.4005
R855 VDPWR.n815 VDPWR.t345 39.4005
R856 VDPWR.n815 VDPWR.t255 39.4005
R857 VDPWR.n813 VDPWR.t265 39.4005
R858 VDPWR.n813 VDPWR.t242 39.4005
R859 VDPWR.n811 VDPWR.t253 39.4005
R860 VDPWR.n811 VDPWR.t427 39.4005
R861 VDPWR.n784 VDPWR.t354 39.4005
R862 VDPWR.n784 VDPWR.t173 39.4005
R863 VDPWR.n651 VDPWR.t324 36.26
R864 VDPWR.t45 VDPWR.t81 32.6341
R865 VDPWR.t47 VDPWR.t136 32.6341
R866 VDPWR.n905 VDPWR.n842 32.2291
R867 VDPWR.n511 VDPWR.n374 32.0005
R868 VDPWR.n516 VDPWR.n374 32.0005
R869 VDPWR.n532 VDPWR.n372 32.0005
R870 VDPWR.n536 VDPWR.n372 32.0005
R871 VDPWR.n537 VDPWR.n536 32.0005
R872 VDPWR.n538 VDPWR.n537 32.0005
R873 VDPWR.n538 VDPWR.n370 32.0005
R874 VDPWR.n959 VDPWR.n292 32.0005
R875 VDPWR.n959 VDPWR.n958 32.0005
R876 VDPWR.n958 VDPWR.n957 32.0005
R877 VDPWR.n957 VDPWR.n294 32.0005
R878 VDPWR.n953 VDPWR.n294 32.0005
R879 VDPWR.n953 VDPWR.n952 32.0005
R880 VDPWR.n952 VDPWR.n951 32.0005
R881 VDPWR.n416 VDPWR.n299 32.0005
R882 VDPWR.n421 VDPWR.n416 32.0005
R883 VDPWR.n422 VDPWR.n421 32.0005
R884 VDPWR.n423 VDPWR.n422 32.0005
R885 VDPWR.n423 VDPWR.n414 32.0005
R886 VDPWR.n427 VDPWR.n414 32.0005
R887 VDPWR.n442 VDPWR.n427 32.0005
R888 VDPWR.n443 VDPWR.n412 32.0005
R889 VDPWR.n462 VDPWR.n454 32.0005
R890 VDPWR.n467 VDPWR.n466 32.0005
R891 VDPWR.n470 VDPWR.n394 32.0005
R892 VDPWR.n474 VDPWR.n394 32.0005
R893 VDPWR.n478 VDPWR.n477 32.0005
R894 VDPWR.n478 VDPWR.n378 32.0005
R895 VDPWR.n482 VDPWR.n378 32.0005
R896 VDPWR.n497 VDPWR.n482 32.0005
R897 VDPWR.n498 VDPWR.n376 32.0005
R898 VDPWR.n502 VDPWR.n376 32.0005
R899 VDPWR.n890 VDPWR.n846 32.0005
R900 VDPWR.n886 VDPWR.n846 32.0005
R901 VDPWR.n886 VDPWR.n885 32.0005
R902 VDPWR.n898 VDPWR.n844 32.0005
R903 VDPWR.n894 VDPWR.n844 32.0005
R904 VDPWR.n894 VDPWR.n893 32.0005
R905 VDPWR.n901 VDPWR.n841 32.0005
R906 VDPWR.n907 VDPWR.n906 32.0005
R907 VDPWR.n913 VDPWR.n835 32.0005
R908 VDPWR.n913 VDPWR.n912 32.0005
R909 VDPWR.n912 VDPWR.n911 32.0005
R910 VDPWR.n919 VDPWR.n832 32.0005
R911 VDPWR.n919 VDPWR.n918 32.0005
R912 VDPWR.n705 VDPWR.n607 32.0005
R913 VDPWR.n700 VDPWR.n607 32.0005
R914 VDPWR.n700 VDPWR.n699 32.0005
R915 VDPWR.n699 VDPWR.n698 32.0005
R916 VDPWR.n698 VDPWR.n610 32.0005
R917 VDPWR.n693 VDPWR.n610 32.0005
R918 VDPWR.n693 VDPWR.n692 32.0005
R919 VDPWR.n692 VDPWR.n691 32.0005
R920 VDPWR.n691 VDPWR.n613 32.0005
R921 VDPWR.n686 VDPWR.n613 32.0005
R922 VDPWR.n686 VDPWR.n685 32.0005
R923 VDPWR.n685 VDPWR.n684 32.0005
R924 VDPWR.n684 VDPWR.n616 32.0005
R925 VDPWR.n679 VDPWR.n616 32.0005
R926 VDPWR.n678 VDPWR.n677 32.0005
R927 VDPWR.n677 VDPWR.n621 32.0005
R928 VDPWR.n245 VDPWR.n23 32.0005
R929 VDPWR.n245 VDPWR.n244 32.0005
R930 VDPWR.n242 VDPWR.n89 32.0005
R931 VDPWR.n238 VDPWR.n89 32.0005
R932 VDPWR.n236 VDPWR.n92 32.0005
R933 VDPWR.n232 VDPWR.n92 32.0005
R934 VDPWR.n232 VDPWR.n231 32.0005
R935 VDPWR.n231 VDPWR.n230 32.0005
R936 VDPWR.n226 VDPWR.n225 32.0005
R937 VDPWR.n225 VDPWR.n224 32.0005
R938 VDPWR.n221 VDPWR.n220 32.0005
R939 VDPWR.n220 VDPWR.n219 32.0005
R940 VDPWR.n215 VDPWR.n214 32.0005
R941 VDPWR.n214 VDPWR.n213 32.0005
R942 VDPWR.n213 VDPWR.n102 32.0005
R943 VDPWR.n209 VDPWR.n102 32.0005
R944 VDPWR.n115 VDPWR.n104 32.0005
R945 VDPWR.n118 VDPWR.n115 32.0005
R946 VDPWR.n122 VDPWR.n112 32.0005
R947 VDPWR.n123 VDPWR.n122 32.0005
R948 VDPWR.n129 VDPWR.n110 32.0005
R949 VDPWR.n130 VDPWR.n129 32.0005
R950 VDPWR.n131 VDPWR.n130 32.0005
R951 VDPWR.n131 VDPWR.n107 32.0005
R952 VDPWR.n199 VDPWR.n108 32.0005
R953 VDPWR.n199 VDPWR.n198 32.0005
R954 VDPWR.n196 VDPWR.n136 32.0005
R955 VDPWR.n192 VDPWR.n136 32.0005
R956 VDPWR.n186 VDPWR.n185 32.0005
R957 VDPWR.n185 VDPWR.n184 32.0005
R958 VDPWR.n184 VDPWR.n139 32.0005
R959 VDPWR.n180 VDPWR.n139 32.0005
R960 VDPWR.n78 VDPWR.n26 32.0005
R961 VDPWR.n82 VDPWR.n26 32.0005
R962 VDPWR.n83 VDPWR.n82 32.0005
R963 VDPWR.n84 VDPWR.n83 32.0005
R964 VDPWR.n84 VDPWR.n24 32.0005
R965 VDPWR.n71 VDPWR.n29 32.0005
R966 VDPWR.n75 VDPWR.n29 32.0005
R967 VDPWR.n76 VDPWR.n75 32.0005
R968 VDPWR.n64 VDPWR.n63 32.0005
R969 VDPWR.n64 VDPWR.n32 32.0005
R970 VDPWR.n68 VDPWR.n32 32.0005
R971 VDPWR.n69 VDPWR.n68 32.0005
R972 VDPWR.n61 VDPWR.n34 32.0005
R973 VDPWR.n57 VDPWR.n55 32.0005
R974 VDPWR.n49 VDPWR.n48 32.0005
R975 VDPWR.n49 VDPWR.n38 32.0005
R976 VDPWR.n53 VDPWR.n38 32.0005
R977 VDPWR.n289 VDPWR.n288 32.0005
R978 VDPWR.n288 VDPWR.n287 32.0005
R979 VDPWR.n287 VDPWR.n4 32.0005
R980 VDPWR.n283 VDPWR.n282 32.0005
R981 VDPWR.n282 VDPWR.n281 32.0005
R982 VDPWR.n281 VDPWR.n8 32.0005
R983 VDPWR.n277 VDPWR.n8 32.0005
R984 VDPWR.n277 VDPWR.n276 32.0005
R985 VDPWR.n276 VDPWR.n275 32.0005
R986 VDPWR.n272 VDPWR.n271 32.0005
R987 VDPWR.n271 VDPWR.n270 32.0005
R988 VDPWR.n270 VDPWR.n13 32.0005
R989 VDPWR.n266 VDPWR.n13 32.0005
R990 VDPWR.n264 VDPWR.n16 32.0005
R991 VDPWR.n260 VDPWR.n16 32.0005
R992 VDPWR.n260 VDPWR.n259 32.0005
R993 VDPWR.n259 VDPWR.n258 32.0005
R994 VDPWR.n258 VDPWR.n18 32.0005
R995 VDPWR.n254 VDPWR.n18 32.0005
R996 VDPWR.n42 VDPWR.n20 32.0005
R997 VDPWR.n42 VDPWR.n41 32.0005
R998 VDPWR.n46 VDPWR.n41 32.0005
R999 VDPWR.n148 VDPWR.n140 30.2632
R1000 VDPWR.n667 VDPWR.n666 30.1875
R1001 VDPWR.n650 VDPWR.n649 30.1875
R1002 VDPWR.n645 VDPWR.n644 30.1875
R1003 VDPWR.n510 VDPWR.n502 28.8005
R1004 VDPWR.n907 VDPWR.n839 28.8005
R1005 VDPWR.n918 VDPWR.n917 28.8005
R1006 VDPWR.n925 VDPWR.n924 28.8005
R1007 VDPWR.n249 VDPWR.n23 28.8005
R1008 VDPWR.n237 VDPWR.n236 28.8005
R1009 VDPWR.n226 VDPWR.n94 28.8005
R1010 VDPWR.n215 VDPWR.n100 28.8005
R1011 VDPWR.n208 VDPWR.n104 28.8005
R1012 VDPWR.n125 VDPWR.n110 28.8005
R1013 VDPWR.n203 VDPWR.n108 28.8005
R1014 VDPWR.n55 VDPWR.n54 28.8005
R1015 VDPWR.n266 VDPWR.n265 28.8005
R1016 VDPWR.n531 VDPWR.n516 25.6005
R1017 VDPWR.n532 VDPWR.n531 25.6005
R1018 VDPWR.n475 VDPWR.n474 25.6005
R1019 VDPWR.t296 VDPWR.t402 25.3822
R1020 VDPWR.t149 VDPWR.t91 25.3822
R1021 VDPWR.n179 VDPWR.n178 24.991
R1022 VDPWR.n162 VDPWR.n137 24.991
R1023 VDPWR.n883 VDPWR.t196 24.6255
R1024 VDPWR.n883 VDPWR.t329 24.6255
R1025 VDPWR.n891 VDPWR.t7 24.6255
R1026 VDPWR.n891 VDPWR.t24 24.6255
R1027 VDPWR.n899 VDPWR.t283 24.6255
R1028 VDPWR.n899 VDPWR.t360 24.6255
R1029 VDPWR.n838 VDPWR.t1 24.6255
R1030 VDPWR.n838 VDPWR.t342 24.6255
R1031 VDPWR.n836 VDPWR.t362 24.6255
R1032 VDPWR.n836 VDPWR.t238 24.6255
R1033 VDPWR.n833 VDPWR.t302 24.6255
R1034 VDPWR.n833 VDPWR.t413 24.6255
R1035 VDPWR.n882 VDPWR.n881 24.361
R1036 VDPWR.n189 VDPWR.n188 24.1894
R1037 VDPWR.n736 VDPWR.n735 22.8576
R1038 VDPWR.n769 VDPWR.n768 22.8576
R1039 VDPWR.n511 VDPWR.n510 22.4005
R1040 VDPWR.n905 VDPWR.n841 22.4005
R1041 VDPWR.n901 VDPWR.n900 22.4005
R1042 VDPWR.n923 VDPWR.n832 22.4005
R1043 VDPWR.n238 VDPWR.n237 22.4005
R1044 VDPWR.n230 VDPWR.n94 22.4005
R1045 VDPWR.n219 VDPWR.n100 22.4005
R1046 VDPWR.n209 VDPWR.n208 22.4005
R1047 VDPWR.n125 VDPWR.n123 22.4005
R1048 VDPWR.n203 VDPWR.n107 22.4005
R1049 VDPWR.n192 VDPWR.n191 22.4005
R1050 VDPWR.n186 VDPWR.n137 22.4005
R1051 VDPWR.n180 VDPWR.n179 22.4005
R1052 VDPWR.n249 VDPWR.n24 22.4005
R1053 VDPWR.n54 VDPWR.n53 22.4005
R1054 VDPWR.n265 VDPWR.n264 22.4005
R1055 VDPWR.n639 VDPWR.n638 22.0449
R1056 VDPWR.n662 VDPWR.t326 19.7005
R1057 VDPWR.n637 VDPWR.t293 19.7005
R1058 VDPWR.n608 VDPWR.t294 19.7005
R1059 VDPWR.n608 VDPWR.t46 19.7005
R1060 VDPWR.n611 VDPWR.t80 19.7005
R1061 VDPWR.n611 VDPWR.t146 19.7005
R1062 VDPWR.n614 VDPWR.t161 19.7005
R1063 VDPWR.n614 VDPWR.t403 19.7005
R1064 VDPWR.n617 VDPWR.t150 19.7005
R1065 VDPWR.n617 VDPWR.t366 19.7005
R1066 VDPWR.n622 VDPWR.t48 19.7005
R1067 VDPWR.n622 VDPWR.t325 19.7005
R1068 VDPWR.n929 VDPWR.n370 19.2005
R1069 VDPWR.n951 VDPWR.n297 19.2005
R1070 VDPWR.n299 VDPWR.n297 19.2005
R1071 VDPWR.n443 VDPWR.n442 19.2005
R1072 VDPWR.n454 VDPWR.n412 19.2005
R1073 VDPWR.n463 VDPWR.n462 19.2005
R1074 VDPWR.n498 VDPWR.n497 19.2005
R1075 VDPWR.n679 VDPWR.n678 19.2005
R1076 VDPWR.n254 VDPWR.n20 19.2005
R1077 VDPWR.t250 VDPWR.t292 18.1303
R1078 VDPWR.t175 VDPWR.t365 18.1303
R1079 VDPWR.n925 VDPWR.n831 17.6005
R1080 VDPWR.n291 VDPWR.n2 17.0989
R1081 VDPWR.n545 VDPWR.t135 17.0848
R1082 VDPWR.n468 VDPWR.n467 16.0005
R1083 VDPWR.n885 VDPWR.n884 16.0005
R1084 VDPWR.n900 VDPWR.n898 16.0005
R1085 VDPWR.n906 VDPWR.n905 16.0005
R1086 VDPWR.n924 VDPWR.n923 16.0005
R1087 VDPWR.n243 VDPWR.n242 16.0005
R1088 VDPWR.n221 VDPWR.n97 16.0005
R1089 VDPWR.n117 VDPWR.n112 16.0005
R1090 VDPWR.n197 VDPWR.n196 16.0005
R1091 VDPWR.n71 VDPWR.n70 16.0005
R1092 VDPWR.n77 VDPWR.n76 16.0005
R1093 VDPWR.n7 VDPWR.n4 16.0005
R1094 VDPWR.n707 VDPWR.n706 15.647
R1095 VDPWR.n857 VDPWR.n831 15.6449
R1096 VDPWR.n881 VDPWR.n880 15.6449
R1097 VDPWR.n927 VDPWR.n926 15.5625
R1098 VDPWR.n962 VDPWR.n291 13.3726
R1099 VDPWR.n733 VDPWR.t190 13.1338
R1100 VDPWR.n733 VDPWR.t232 13.1338
R1101 VDPWR.n731 VDPWR.t187 13.1338
R1102 VDPWR.n731 VDPWR.t37 13.1338
R1103 VDPWR.n729 VDPWR.t381 13.1338
R1104 VDPWR.n729 VDPWR.t383 13.1338
R1105 VDPWR.n727 VDPWR.t64 13.1338
R1106 VDPWR.n727 VDPWR.t30 13.1338
R1107 VDPWR.n725 VDPWR.t184 13.1338
R1108 VDPWR.n725 VDPWR.t420 13.1338
R1109 VDPWR.n723 VDPWR.t422 13.1338
R1110 VDPWR.n723 VDPWR.t214 13.1338
R1111 VDPWR.n721 VDPWR.t133 13.1338
R1112 VDPWR.n721 VDPWR.t14 13.1338
R1113 VDPWR.n708 VDPWR.t16 13.1338
R1114 VDPWR.n708 VDPWR.t54 13.1338
R1115 VDPWR.n466 VDPWR.n410 12.8005
R1116 VDPWR.n470 VDPWR.n469 12.8005
R1117 VDPWR.n56 VDPWR.n34 12.8005
R1118 VDPWR.n62 VDPWR.n61 12.8005
R1119 VDPWR.n272 VDPWR.n11 12.8005
R1120 VDPWR.n962 VDPWR.n961 11.8717
R1121 VDPWR.t396 VDPWR.n944 11.4924
R1122 VDPWR.n943 VDPWR.t392 11.4924
R1123 VDPWR.t127 VDPWR.n942 11.4924
R1124 VDPWR.n941 VDPWR.t207 11.4924
R1125 VDPWR.t140 VDPWR.n940 11.4924
R1126 VDPWR.n735 VDPWR.n734 11.0565
R1127 VDPWR.t177 VDPWR.t79 10.8784
R1128 VDPWR.n770 VDPWR.n769 10.8682
R1129 VDPWR.n638 VDPWR.n606 9.613
R1130 VDPWR.n917 VDPWR.n835 9.6005
R1131 VDPWR.n911 VDPWR.n839 9.6005
R1132 VDPWR.n666 VDPWR.n624 9.6005
R1133 VDPWR.n649 VDPWR.n648 9.6005
R1134 VDPWR.n644 VDPWR.n643 9.6005
R1135 VDPWR.n671 VDPWR.n670 9.6005
R1136 VDPWR.n48 VDPWR.n47 9.6005
R1137 VDPWR.n289 VDPWR.n2 9.6005
R1138 VDPWR.n47 VDPWR.n46 9.6005
R1139 VDPWR.n576 VDPWR.n552 9.50883
R1140 VDPWR.n602 VDPWR.n548 9.50883
R1141 VDPWR.n768 VDPWR.n767 9.50883
R1142 VDPWR.n760 VDPWR.n759 9.50883
R1143 VDPWR.n738 VDPWR.n736 9.50883
R1144 VDPWR.n749 VDPWR.n748 9.50883
R1145 VDPWR.n780 VDPWR.n772 9.50883
R1146 VDPWR.n576 VDPWR.n575 9.3005
R1147 VDPWR.n602 VDPWR.n601 9.3005
R1148 VDPWR.n741 VDPWR.n738 9.3005
R1149 VDPWR.n737 VDPWR.n720 9.3005
R1150 VDPWR.n746 VDPWR.n719 9.3005
R1151 VDPWR.n748 VDPWR.n747 9.3005
R1152 VDPWR.n767 VDPWR.n766 9.3005
R1153 VDPWR.n713 VDPWR.n712 9.3005
R1154 VDPWR.n757 VDPWR.n754 9.3005
R1155 VDPWR.n759 VDPWR.n758 9.3005
R1156 VDPWR.n780 VDPWR.n779 9.3005
R1157 VDPWR.n923 VDPWR.n922 9.3005
R1158 VDPWR.n905 VDPWR.n904 9.3005
R1159 VDPWR.n900 VDPWR.n843 9.3005
R1160 VDPWR.n885 VDPWR.n847 9.3005
R1161 VDPWR.n887 VDPWR.n886 9.3005
R1162 VDPWR.n888 VDPWR.n846 9.3005
R1163 VDPWR.n890 VDPWR.n889 9.3005
R1164 VDPWR.n893 VDPWR.n845 9.3005
R1165 VDPWR.n895 VDPWR.n894 9.3005
R1166 VDPWR.n896 VDPWR.n844 9.3005
R1167 VDPWR.n898 VDPWR.n897 9.3005
R1168 VDPWR.n902 VDPWR.n901 9.3005
R1169 VDPWR.n903 VDPWR.n841 9.3005
R1170 VDPWR.n906 VDPWR.n840 9.3005
R1171 VDPWR.n908 VDPWR.n907 9.3005
R1172 VDPWR.n909 VDPWR.n839 9.3005
R1173 VDPWR.n911 VDPWR.n910 9.3005
R1174 VDPWR.n912 VDPWR.n837 9.3005
R1175 VDPWR.n914 VDPWR.n913 9.3005
R1176 VDPWR.n915 VDPWR.n835 9.3005
R1177 VDPWR.n917 VDPWR.n916 9.3005
R1178 VDPWR.n918 VDPWR.n834 9.3005
R1179 VDPWR.n920 VDPWR.n919 9.3005
R1180 VDPWR.n921 VDPWR.n832 9.3005
R1181 VDPWR.n924 VDPWR.n830 9.3005
R1182 VDPWR.n675 VDPWR.n621 9.3005
R1183 VDPWR.n677 VDPWR.n676 9.3005
R1184 VDPWR.n678 VDPWR.n618 9.3005
R1185 VDPWR.n680 VDPWR.n679 9.3005
R1186 VDPWR.n682 VDPWR.n616 9.3005
R1187 VDPWR.n684 VDPWR.n683 9.3005
R1188 VDPWR.n685 VDPWR.n615 9.3005
R1189 VDPWR.n687 VDPWR.n686 9.3005
R1190 VDPWR.n689 VDPWR.n613 9.3005
R1191 VDPWR.n691 VDPWR.n690 9.3005
R1192 VDPWR.n692 VDPWR.n612 9.3005
R1193 VDPWR.n694 VDPWR.n693 9.3005
R1194 VDPWR.n696 VDPWR.n610 9.3005
R1195 VDPWR.n698 VDPWR.n697 9.3005
R1196 VDPWR.n699 VDPWR.n609 9.3005
R1197 VDPWR.n701 VDPWR.n700 9.3005
R1198 VDPWR.n703 VDPWR.n607 9.3005
R1199 VDPWR.n705 VDPWR.n704 9.3005
R1200 VDPWR.n417 VDPWR.n297 9.3005
R1201 VDPWR.n540 VDPWR.n370 9.3005
R1202 VDPWR.n539 VDPWR.n538 9.3005
R1203 VDPWR.n537 VDPWR.n371 9.3005
R1204 VDPWR.n536 VDPWR.n535 9.3005
R1205 VDPWR.n534 VDPWR.n372 9.3005
R1206 VDPWR.n533 VDPWR.n532 9.3005
R1207 VDPWR.n531 VDPWR.n373 9.3005
R1208 VDPWR.n516 VDPWR.n515 9.3005
R1209 VDPWR.n514 VDPWR.n374 9.3005
R1210 VDPWR.n512 VDPWR.n511 9.3005
R1211 VDPWR.n510 VDPWR.n375 9.3005
R1212 VDPWR.n502 VDPWR.n501 9.3005
R1213 VDPWR.n500 VDPWR.n376 9.3005
R1214 VDPWR.n499 VDPWR.n498 9.3005
R1215 VDPWR.n497 VDPWR.n377 9.3005
R1216 VDPWR.n482 VDPWR.n481 9.3005
R1217 VDPWR.n480 VDPWR.n378 9.3005
R1218 VDPWR.n479 VDPWR.n478 9.3005
R1219 VDPWR.n477 VDPWR.n379 9.3005
R1220 VDPWR.n474 VDPWR.n473 9.3005
R1221 VDPWR.n472 VDPWR.n394 9.3005
R1222 VDPWR.n471 VDPWR.n470 9.3005
R1223 VDPWR.n467 VDPWR.n395 9.3005
R1224 VDPWR.n466 VDPWR.n465 9.3005
R1225 VDPWR.n464 VDPWR.n463 9.3005
R1226 VDPWR.n462 VDPWR.n411 9.3005
R1227 VDPWR.n454 VDPWR.n446 9.3005
R1228 VDPWR.n445 VDPWR.n412 9.3005
R1229 VDPWR.n444 VDPWR.n443 9.3005
R1230 VDPWR.n442 VDPWR.n413 9.3005
R1231 VDPWR.n427 VDPWR.n426 9.3005
R1232 VDPWR.n425 VDPWR.n414 9.3005
R1233 VDPWR.n424 VDPWR.n423 9.3005
R1234 VDPWR.n422 VDPWR.n415 9.3005
R1235 VDPWR.n421 VDPWR.n420 9.3005
R1236 VDPWR.n419 VDPWR.n416 9.3005
R1237 VDPWR.n418 VDPWR.n299 9.3005
R1238 VDPWR.n951 VDPWR.n296 9.3005
R1239 VDPWR.n952 VDPWR.n295 9.3005
R1240 VDPWR.n954 VDPWR.n953 9.3005
R1241 VDPWR.n955 VDPWR.n294 9.3005
R1242 VDPWR.n957 VDPWR.n956 9.3005
R1243 VDPWR.n958 VDPWR.n293 9.3005
R1244 VDPWR.n960 VDPWR.n959 9.3005
R1245 VDPWR.n181 VDPWR.n180 9.3005
R1246 VDPWR.n182 VDPWR.n139 9.3005
R1247 VDPWR.n184 VDPWR.n183 9.3005
R1248 VDPWR.n185 VDPWR.n138 9.3005
R1249 VDPWR.n187 VDPWR.n186 9.3005
R1250 VDPWR.n193 VDPWR.n192 9.3005
R1251 VDPWR.n194 VDPWR.n136 9.3005
R1252 VDPWR.n196 VDPWR.n195 9.3005
R1253 VDPWR.n198 VDPWR.n134 9.3005
R1254 VDPWR.n200 VDPWR.n199 9.3005
R1255 VDPWR.n201 VDPWR.n108 9.3005
R1256 VDPWR.n203 VDPWR.n202 9.3005
R1257 VDPWR.n133 VDPWR.n107 9.3005
R1258 VDPWR.n132 VDPWR.n131 9.3005
R1259 VDPWR.n130 VDPWR.n109 9.3005
R1260 VDPWR.n129 VDPWR.n128 9.3005
R1261 VDPWR.n127 VDPWR.n110 9.3005
R1262 VDPWR.n126 VDPWR.n125 9.3005
R1263 VDPWR.n123 VDPWR.n111 9.3005
R1264 VDPWR.n122 VDPWR.n121 9.3005
R1265 VDPWR.n120 VDPWR.n112 9.3005
R1266 VDPWR.n119 VDPWR.n118 9.3005
R1267 VDPWR.n115 VDPWR.n114 9.3005
R1268 VDPWR.n113 VDPWR.n104 9.3005
R1269 VDPWR.n208 VDPWR.n103 9.3005
R1270 VDPWR.n210 VDPWR.n209 9.3005
R1271 VDPWR.n211 VDPWR.n102 9.3005
R1272 VDPWR.n213 VDPWR.n212 9.3005
R1273 VDPWR.n214 VDPWR.n101 9.3005
R1274 VDPWR.n216 VDPWR.n215 9.3005
R1275 VDPWR.n217 VDPWR.n100 9.3005
R1276 VDPWR.n219 VDPWR.n218 9.3005
R1277 VDPWR.n220 VDPWR.n98 9.3005
R1278 VDPWR.n222 VDPWR.n221 9.3005
R1279 VDPWR.n224 VDPWR.n223 9.3005
R1280 VDPWR.n225 VDPWR.n95 9.3005
R1281 VDPWR.n227 VDPWR.n226 9.3005
R1282 VDPWR.n228 VDPWR.n94 9.3005
R1283 VDPWR.n230 VDPWR.n229 9.3005
R1284 VDPWR.n231 VDPWR.n93 9.3005
R1285 VDPWR.n233 VDPWR.n232 9.3005
R1286 VDPWR.n234 VDPWR.n92 9.3005
R1287 VDPWR.n236 VDPWR.n235 9.3005
R1288 VDPWR.n237 VDPWR.n90 9.3005
R1289 VDPWR.n239 VDPWR.n238 9.3005
R1290 VDPWR.n240 VDPWR.n89 9.3005
R1291 VDPWR.n242 VDPWR.n241 9.3005
R1292 VDPWR.n244 VDPWR.n87 9.3005
R1293 VDPWR.n246 VDPWR.n245 9.3005
R1294 VDPWR.n247 VDPWR.n23 9.3005
R1295 VDPWR.n249 VDPWR.n248 9.3005
R1296 VDPWR.n86 VDPWR.n24 9.3005
R1297 VDPWR.n85 VDPWR.n84 9.3005
R1298 VDPWR.n83 VDPWR.n25 9.3005
R1299 VDPWR.n82 VDPWR.n81 9.3005
R1300 VDPWR.n80 VDPWR.n26 9.3005
R1301 VDPWR.n79 VDPWR.n78 9.3005
R1302 VDPWR.n76 VDPWR.n27 9.3005
R1303 VDPWR.n75 VDPWR.n74 9.3005
R1304 VDPWR.n73 VDPWR.n29 9.3005
R1305 VDPWR.n72 VDPWR.n71 9.3005
R1306 VDPWR.n69 VDPWR.n30 9.3005
R1307 VDPWR.n68 VDPWR.n67 9.3005
R1308 VDPWR.n66 VDPWR.n32 9.3005
R1309 VDPWR.n65 VDPWR.n64 9.3005
R1310 VDPWR.n63 VDPWR.n33 9.3005
R1311 VDPWR.n61 VDPWR.n60 9.3005
R1312 VDPWR.n59 VDPWR.n34 9.3005
R1313 VDPWR.n58 VDPWR.n57 9.3005
R1314 VDPWR.n55 VDPWR.n35 9.3005
R1315 VDPWR.n54 VDPWR.n36 9.3005
R1316 VDPWR.n53 VDPWR.n52 9.3005
R1317 VDPWR.n51 VDPWR.n38 9.3005
R1318 VDPWR.n50 VDPWR.n49 9.3005
R1319 VDPWR.n48 VDPWR.n39 9.3005
R1320 VDPWR.n46 VDPWR.n45 9.3005
R1321 VDPWR.n44 VDPWR.n41 9.3005
R1322 VDPWR.n43 VDPWR.n42 9.3005
R1323 VDPWR.n20 VDPWR.n19 9.3005
R1324 VDPWR.n255 VDPWR.n254 9.3005
R1325 VDPWR.n256 VDPWR.n18 9.3005
R1326 VDPWR.n258 VDPWR.n257 9.3005
R1327 VDPWR.n259 VDPWR.n17 9.3005
R1328 VDPWR.n261 VDPWR.n260 9.3005
R1329 VDPWR.n262 VDPWR.n16 9.3005
R1330 VDPWR.n264 VDPWR.n263 9.3005
R1331 VDPWR.n265 VDPWR.n14 9.3005
R1332 VDPWR.n267 VDPWR.n266 9.3005
R1333 VDPWR.n268 VDPWR.n13 9.3005
R1334 VDPWR.n270 VDPWR.n269 9.3005
R1335 VDPWR.n271 VDPWR.n12 9.3005
R1336 VDPWR.n273 VDPWR.n272 9.3005
R1337 VDPWR.n275 VDPWR.n274 9.3005
R1338 VDPWR.n276 VDPWR.n9 9.3005
R1339 VDPWR.n278 VDPWR.n277 9.3005
R1340 VDPWR.n279 VDPWR.n8 9.3005
R1341 VDPWR.n281 VDPWR.n280 9.3005
R1342 VDPWR.n282 VDPWR.n5 9.3005
R1343 VDPWR.n284 VDPWR.n283 9.3005
R1344 VDPWR.n285 VDPWR.n4 9.3005
R1345 VDPWR.n287 VDPWR.n286 9.3005
R1346 VDPWR.n288 VDPWR.n3 9.3005
R1347 VDPWR.n290 VDPWR.n289 9.3005
R1348 VDPWR.n383 VDPWR.n380 9.14336
R1349 VDPWR.n399 VDPWR.n396 9.14336
R1350 VDPWR.n406 VDPWR.n403 9.14336
R1351 VDPWR.n390 VDPWR.n387 9.14336
R1352 VDPWR.n317 VDPWR.n314 9.14336
R1353 VDPWR.n307 VDPWR.n305 9.14336
R1354 VDPWR.n438 VDPWR.n435 9.14336
R1355 VDPWR.n431 VDPWR.n428 9.14336
R1356 VDPWR.n450 VDPWR.n447 9.14336
R1357 VDPWR.n458 VDPWR.n455 9.14336
R1358 VDPWR.n741 VDPWR.n720 9.14336
R1359 VDPWR.n746 VDPWR.n720 9.14336
R1360 VDPWR.n747 VDPWR.n746 9.14336
R1361 VDPWR.n766 VDPWR.n713 9.14336
R1362 VDPWR.n757 VDPWR.n713 9.14336
R1363 VDPWR.n758 VDPWR.n757 9.14336
R1364 VDPWR.n175 VDPWR.n174 9.14336
R1365 VDPWR.n165 VDPWR.n164 9.14336
R1366 VDPWR.n928 VDPWR.n927 8.93298
R1367 VDPWR.t234 VDPWR.t368 7.66179
R1368 VDPWR.n929 VDPWR.n928 7.49891
R1369 VDPWR.n191 VDPWR.n189 7.37605
R1370 VDPWR.n668 VDPWR.n665 7.25241
R1371 VDPWR.n493 VDPWR.n490 7.11161
R1372 VDPWR.n486 VDPWR.n483 7.11161
R1373 VDPWR.n506 VDPWR.n503 7.11161
R1374 VDPWR.n527 VDPWR.n524 7.11161
R1375 VDPWR.n520 VDPWR.n517 7.11161
R1376 VDPWR.n932 VDPWR.n369 7.11161
R1377 VDPWR.n854 VDPWR.n852 7.11161
R1378 VDPWR.n875 VDPWR.n874 7.11161
R1379 VDPWR.n657 VDPWR.n655 7.11161
R1380 VDPWR.n661 VDPWR.n660 7.11161
R1381 VDPWR.n635 VDPWR.n632 7.11161
R1382 VDPWR.n639 VDPWR.n630 7.11161
R1383 VDPWR.n829 VDPWR.n828 7.098
R1384 VDPWR.n188 VDPWR.n137 7.05969
R1385 VDPWR.n179 VDPWR.n140 7.05957
R1386 VDPWR.n961 VDPWR.n292 6.87881
R1387 VDPWR.n884 VDPWR.n882 6.54033
R1388 VDPWR.n463 VDPWR.n410 6.4005
R1389 VDPWR.n63 VDPWR.n62 6.4005
R1390 VDPWR.n57 VDPWR.n56 6.4005
R1391 VDPWR.n275 VDPWR.n11 6.4005
R1392 VDPWR.n926 VDPWR.n925 5.98166
R1393 VDPWR.n337 VDPWR.n336 5.81868
R1394 VDPWR.n330 VDPWR.n329 5.81868
R1395 VDPWR.n151 VDPWR.n150 5.81868
R1396 VDPWR.n386 VDPWR.n385 5.33286
R1397 VDPWR.n402 VDPWR.n401 5.33286
R1398 VDPWR.n409 VDPWR.n408 5.33286
R1399 VDPWR.n393 VDPWR.n392 5.33286
R1400 VDPWR.n318 VDPWR.n315 5.33286
R1401 VDPWR.n310 VDPWR.n309 5.33286
R1402 VDPWR.n441 VDPWR.n440 5.33286
R1403 VDPWR.n434 VDPWR.n433 5.33286
R1404 VDPWR.n453 VDPWR.n452 5.33286
R1405 VDPWR.n461 VDPWR.n460 5.33286
R1406 VDPWR.n742 VDPWR.n736 5.33286
R1407 VDPWR.n749 VDPWR.n718 5.33286
R1408 VDPWR.n768 VDPWR.n710 5.33286
R1409 VDPWR.n760 VDPWR.n753 5.33286
R1410 VDPWR.n167 VDPWR.n166 5.33286
R1411 VDPWR.n178 VDPWR.n141 5.33286
R1412 VDPWR.n173 VDPWR.n172 5.33286
R1413 VDPWR.n163 VDPWR.n162 5.33286
R1414 VDPWR.n802 VDPWR.n801 4.84425
R1415 VDPWR.n971 VDPWR.n962 4.80604
R1416 VDPWR.n804 VDPWR.n803 4.73979
R1417 VDPWR.n808 VDPWR.n791 4.73979
R1418 VDPWR.n822 VDPWR.n821 4.73979
R1419 VDPWR.n826 VDPWR.n786 4.73979
R1420 VDPWR.n803 VDPWR.n792 4.6505
R1421 VDPWR.n808 VDPWR.n807 4.6505
R1422 VDPWR.n821 VDPWR.n787 4.6505
R1423 VDPWR.n826 VDPWR.n825 4.6505
R1424 VDPWR.n869 VDPWR.n862 4.57193
R1425 VDPWR.n804 VDPWR.n793 4.54311
R1426 VDPWR.n793 VDPWR.n792 4.54311
R1427 VDPWR.n822 VDPWR.n788 4.54311
R1428 VDPWR.n788 VDPWR.n787 4.54311
R1429 VDPWR.n828 VDPWR.n827 4.5005
R1430 VDPWR.n820 VDPWR.n819 4.5005
R1431 VDPWR.n810 VDPWR.n809 4.5005
R1432 VDPWR.n575 VDPWR.n574 4.48641
R1433 VDPWR.n574 VDPWR.n552 4.48641
R1434 VDPWR.n601 VDPWR.n600 4.48641
R1435 VDPWR.n600 VDPWR.n548 4.48641
R1436 VDPWR.n779 VDPWR.n778 4.48641
R1437 VDPWR.n778 VDPWR.n772 4.48641
R1438 VDPWR.n807 VDPWR.n806 4.48641
R1439 VDPWR.n806 VDPWR.n791 4.48641
R1440 VDPWR.n825 VDPWR.n824 4.48641
R1441 VDPWR.n824 VDPWR.n786 4.48641
R1442 VDPWR.n496 VDPWR.n495 4.0479
R1443 VDPWR.n489 VDPWR.n488 4.0479
R1444 VDPWR.n509 VDPWR.n508 4.0479
R1445 VDPWR.n530 VDPWR.n529 4.0479
R1446 VDPWR.n523 VDPWR.n522 4.0479
R1447 VDPWR.n933 VDPWR.n930 4.0479
R1448 VDPWR.n857 VDPWR.n856 4.0479
R1449 VDPWR.n880 VDPWR.n848 4.0479
R1450 VDPWR VDPWR.n972 4.02487
R1451 VDPWR.n384 VDPWR.n383 3.75335
R1452 VDPWR.n385 VDPWR.n380 3.75335
R1453 VDPWR.n400 VDPWR.n399 3.75335
R1454 VDPWR.n401 VDPWR.n396 3.75335
R1455 VDPWR.n408 VDPWR.n403 3.75335
R1456 VDPWR.n407 VDPWR.n406 3.75335
R1457 VDPWR.n392 VDPWR.n387 3.75335
R1458 VDPWR.n391 VDPWR.n390 3.75335
R1459 VDPWR.n319 VDPWR.n314 3.75335
R1460 VDPWR.n318 VDPWR.n317 3.75335
R1461 VDPWR.n309 VDPWR.n305 3.75335
R1462 VDPWR.n308 VDPWR.n307 3.75335
R1463 VDPWR.n439 VDPWR.n438 3.75335
R1464 VDPWR.n440 VDPWR.n435 3.75335
R1465 VDPWR.n433 VDPWR.n428 3.75335
R1466 VDPWR.n432 VDPWR.n431 3.75335
R1467 VDPWR.n451 VDPWR.n450 3.75335
R1468 VDPWR.n452 VDPWR.n447 3.75335
R1469 VDPWR.n460 VDPWR.n455 3.75335
R1470 VDPWR.n459 VDPWR.n458 3.75335
R1471 VDPWR.n747 VDPWR.n718 3.75335
R1472 VDPWR.n742 VDPWR.n741 3.75335
R1473 VDPWR.n758 VDPWR.n753 3.75335
R1474 VDPWR.n766 VDPWR.n710 3.75335
R1475 VDPWR.n174 VDPWR.n173 3.75335
R1476 VDPWR.n175 VDPWR.n141 3.75335
R1477 VDPWR.n166 VDPWR.n165 3.75335
R1478 VDPWR.n164 VDPWR.n163 3.75335
R1479 VDPWR.n657 VDPWR.n656 3.53508
R1480 VDPWR.n660 VDPWR.n656 3.53508
R1481 VDPWR.n663 VDPWR.n655 3.53508
R1482 VDPWR.n636 VDPWR.n635 3.53508
R1483 VDPWR.n636 VDPWR.n630 3.53508
R1484 VDPWR.n632 VDPWR.n631 3.53508
R1485 VDPWR.n775 VDPWR.n774 3.46433
R1486 VDPWR.n571 VDPWR.n570 3.41464
R1487 VDPWR.n597 VDPWR.n596 3.41464
R1488 VDPWR.n967 VDPWR.n964 3.4105
R1489 VDPWR.n969 VDPWR.n964 3.4105
R1490 VDPWR.n971 VDPWR.n964 3.4105
R1491 VDPWR.n970 VDPWR.n969 3.4105
R1492 VDPWR.n971 VDPWR.n970 3.4105
R1493 VDPWR.n969 VDPWR.n963 3.4105
R1494 VDPWR.n971 VDPWR.n963 3.4105
R1495 VDPWR.n972 VDPWR.n971 3.4105
R1496 VDPWR.n949 VDPWR.n301 3.40194
R1497 VDPWR.n339 VDPWR.n335 3.40194
R1498 VDPWR.n327 VDPWR.n326 3.40194
R1499 VDPWR.n332 VDPWR.n324 3.40194
R1500 VDPWR.n149 VDPWR.n148 3.40194
R1501 VDPWR.n154 VDPWR.n143 3.40194
R1502 VDPWR.n469 VDPWR.n468 3.2005
R1503 VDPWR.n476 VDPWR.n475 3.2005
R1504 VDPWR.n477 VDPWR.n476 3.2005
R1505 VDPWR.n892 VDPWR.n890 3.2005
R1506 VDPWR.n893 VDPWR.n892 3.2005
R1507 VDPWR.n244 VDPWR.n243 3.2005
R1508 VDPWR.n224 VDPWR.n97 3.2005
R1509 VDPWR.n118 VDPWR.n117 3.2005
R1510 VDPWR.n198 VDPWR.n197 3.2005
R1511 VDPWR.n78 VDPWR.n77 3.2005
R1512 VDPWR.n70 VDPWR.n69 3.2005
R1513 VDPWR.n283 VDPWR.n7 3.2005
R1514 VDPWR.n571 VDPWR.n553 3.11118
R1515 VDPWR.n598 VDPWR.n597 3.11118
R1516 VDPWR.n572 VDPWR.n571 3.04304
R1517 VDPWR.n597 VDPWR.n549 3.04304
R1518 VDPWR.n494 VDPWR.n493 3.02841
R1519 VDPWR.n495 VDPWR.n490 3.02841
R1520 VDPWR.n488 VDPWR.n483 3.02841
R1521 VDPWR.n487 VDPWR.n486 3.02841
R1522 VDPWR.n507 VDPWR.n506 3.02841
R1523 VDPWR.n508 VDPWR.n503 3.02841
R1524 VDPWR.n528 VDPWR.n527 3.02841
R1525 VDPWR.n529 VDPWR.n524 3.02841
R1526 VDPWR.n522 VDPWR.n517 3.02841
R1527 VDPWR.n521 VDPWR.n520 3.02841
R1528 VDPWR.n934 VDPWR.n369 3.02841
R1529 VDPWR.n933 VDPWR.n932 3.02841
R1530 VDPWR.n856 VDPWR.n852 3.02841
R1531 VDPWR.n855 VDPWR.n854 3.02841
R1532 VDPWR.n874 VDPWR.n848 3.02841
R1533 VDPWR.n875 VDPWR.n873 3.02841
R1534 VDPWR.n776 VDPWR.n775 2.96855
R1535 VDPWR.n775 VDPWR.n773 2.90353
R1536 VDPWR.n866 VDPWR.n865 2.6074
R1537 VDPWR.n863 VDPWR.n842 2.6074
R1538 VDPWR.n605 VDPWR.n545 2.47421
R1539 VDPWR.n337 VDPWR.n335 2.39444
R1540 VDPWR.n336 VDPWR.n301 2.39444
R1541 VDPWR.n330 VDPWR.n324 2.39444
R1542 VDPWR.n329 VDPWR.n327 2.39444
R1543 VDPWR.n151 VDPWR.n143 2.39444
R1544 VDPWR.n150 VDPWR.n149 2.39444
R1545 VDPWR.n783 VDPWR.n782 2.36621
R1546 VDPWR.n605 VDPWR.n604 2.35058
R1547 VDPWR.n950 VDPWR.n949 2.32777
R1548 VDPWR.n332 VDPWR.n298 2.32777
R1549 VDPWR.n782 VDPWR.n781 2.00667
R1550 VDPWR.n869 VDPWR.n863 1.9508
R1551 VDPWR.n865 VDPWR.n862 1.9508
R1552 VDPWR.n774 VDPWR.n771 1.94319
R1553 VDPWR.n570 VDPWR.n569 1.90331
R1554 VDPWR.n604 VDPWR.n603 1.82095
R1555 VDPWR.n578 VDPWR.n577 1.77831
R1556 VDPWR.n596 VDPWR.n595 1.77831
R1557 VDPWR.n966 VDPWR.n965 1.70307
R1558 VDPWR.n968 VDPWR.n967 1.70307
R1559 VDPWR.n972 VDPWR.n1 1.70307
R1560 VDPWR.n965 VDPWR.n0 1.70307
R1561 VDPWR.n545 VDPWR.n543 1.05389
R1562 VDPWR.n819 VDPWR.n810 0.90675
R1563 VDPWR.n542 VDPWR.n541 0.75233
R1564 VDPWR.n882 VDPWR.n847 0.703395
R1565 VDPWR.n543 VDPWR.n542 0.648391
R1566 VDPWR.n783 VDPWR.n707 0.480239
R1567 VDPWR.n927 VDPWR.n829 0.4094
R1568 VDPWR.n801 VDPWR.n799 0.34425
R1569 VDPWR.n799 VDPWR.n797 0.34425
R1570 VDPWR.n797 VDPWR.n795 0.34425
R1571 VDPWR.n795 VDPWR.n790 0.34425
R1572 VDPWR.n810 VDPWR.n790 0.34425
R1573 VDPWR.n819 VDPWR.n818 0.34425
R1574 VDPWR.n818 VDPWR.n816 0.34425
R1575 VDPWR.n816 VDPWR.n814 0.34425
R1576 VDPWR.n814 VDPWR.n812 0.34425
R1577 VDPWR.n812 VDPWR.n785 0.34425
R1578 VDPWR.n828 VDPWR.n785 0.34425
R1579 VDPWR.n595 VDPWR.n578 0.333833
R1580 VDPWR.n771 VDPWR.n770 0.328625
R1581 VDPWR.n577 VDPWR.n576 0.2505
R1582 VDPWR.n603 VDPWR.n602 0.2505
R1583 VDPWR.n781 VDPWR.n780 0.2505
R1584 VDPWR.n829 VDPWR.n783 0.245239
R1585 VDPWR.n782 VDPWR.n771 0.229667
R1586 VDPWR.n926 VDPWR.n830 0.224356
R1587 VDPWR.n767 VDPWR.n712 0.208833
R1588 VDPWR.n754 VDPWR.n712 0.208833
R1589 VDPWR.n759 VDPWR.n754 0.208833
R1590 VDPWR.n738 VDPWR.n737 0.208833
R1591 VDPWR.n737 VDPWR.n719 0.208833
R1592 VDPWR.n748 VDPWR.n719 0.208833
R1593 VDPWR.n961 VDPWR.n960 0.206321
R1594 VDPWR.n181 VDPWR.n140 0.203053
R1595 VDPWR.n707 VDPWR.n605 0.202939
R1596 VDPWR.n188 VDPWR.n187 0.202927
R1597 VDPWR.n193 VDPWR.n189 0.196005
R1598 VDPWR.n928 VDPWR.n540 0.193961
R1599 VDPWR.n291 VDPWR.n290 0.193958
R1600 VDPWR.n734 VDPWR.n732 0.188
R1601 VDPWR.n732 VDPWR.n730 0.188
R1602 VDPWR.n730 VDPWR.n728 0.188
R1603 VDPWR.n728 VDPWR.n726 0.188
R1604 VDPWR.n726 VDPWR.n724 0.188
R1605 VDPWR.n724 VDPWR.n722 0.188
R1606 VDPWR.n722 VDPWR.n709 0.188
R1607 VDPWR.n770 VDPWR.n709 0.188
R1608 VDPWR.n809 VDPWR.n808 0.182048
R1609 VDPWR.n827 VDPWR.n826 0.182048
R1610 VDPWR.n803 VDPWR.n802 0.182048
R1611 VDPWR.n821 VDPWR.n820 0.182048
R1612 VDPWR.t117 VDPWR.t55 0.1603
R1613 VDPWR.t373 VDPWR.t117 0.1603
R1614 VDPWR.t116 VDPWR.t373 0.1603
R1615 VDPWR.t376 VDPWR.t116 0.1603
R1616 VDPWR.t65 VDPWR.t376 0.1603
R1617 VDPWR.t233 VDPWR.t65 0.1603
R1618 VDPWR.t38 VDPWR.t233 0.1603
R1619 VDPWR.t182 VDPWR.t38 0.1603
R1620 VDPWR.t121 VDPWR.t372 0.1603
R1621 VDPWR.t377 VDPWR.t121 0.1603
R1622 VDPWR.t188 VDPWR.t377 0.1603
R1623 VDPWR.t131 VDPWR.t188 0.1603
R1624 VDPWR.t215 VDPWR.t131 0.1603
R1625 VDPWR.t134 VDPWR.t215 0.1603
R1626 VDPWR.t31 VDPWR.t134 0.1603
R1627 VDPWR.t135 VDPWR.t31 0.1603
R1628 VDPWR.t120 VDPWR.n544 0.159278
R1629 VDPWR.n922 VDPWR.n830 0.15675
R1630 VDPWR.n922 VDPWR.n921 0.15675
R1631 VDPWR.n921 VDPWR.n920 0.15675
R1632 VDPWR.n920 VDPWR.n834 0.15675
R1633 VDPWR.n916 VDPWR.n834 0.15675
R1634 VDPWR.n916 VDPWR.n915 0.15675
R1635 VDPWR.n915 VDPWR.n914 0.15675
R1636 VDPWR.n914 VDPWR.n837 0.15675
R1637 VDPWR.n910 VDPWR.n837 0.15675
R1638 VDPWR.n910 VDPWR.n909 0.15675
R1639 VDPWR.n909 VDPWR.n908 0.15675
R1640 VDPWR.n908 VDPWR.n840 0.15675
R1641 VDPWR.n904 VDPWR.n840 0.15675
R1642 VDPWR.n904 VDPWR.n903 0.15675
R1643 VDPWR.n903 VDPWR.n902 0.15675
R1644 VDPWR.n902 VDPWR.n843 0.15675
R1645 VDPWR.n897 VDPWR.n843 0.15675
R1646 VDPWR.n897 VDPWR.n896 0.15675
R1647 VDPWR.n896 VDPWR.n895 0.15675
R1648 VDPWR.n895 VDPWR.n845 0.15675
R1649 VDPWR.n889 VDPWR.n845 0.15675
R1650 VDPWR.n889 VDPWR.n888 0.15675
R1651 VDPWR.n888 VDPWR.n887 0.15675
R1652 VDPWR.n887 VDPWR.n847 0.15675
R1653 VDPWR.n704 VDPWR.n703 0.15675
R1654 VDPWR.n701 VDPWR.n609 0.15675
R1655 VDPWR.n697 VDPWR.n609 0.15675
R1656 VDPWR.n697 VDPWR.n696 0.15675
R1657 VDPWR.n694 VDPWR.n612 0.15675
R1658 VDPWR.n690 VDPWR.n612 0.15675
R1659 VDPWR.n690 VDPWR.n689 0.15675
R1660 VDPWR.n687 VDPWR.n615 0.15675
R1661 VDPWR.n683 VDPWR.n615 0.15675
R1662 VDPWR.n683 VDPWR.n682 0.15675
R1663 VDPWR.n680 VDPWR.n618 0.15675
R1664 VDPWR.n676 VDPWR.n618 0.15675
R1665 VDPWR.n676 VDPWR.n675 0.15675
R1666 VDPWR.n960 VDPWR.n293 0.15675
R1667 VDPWR.n956 VDPWR.n293 0.15675
R1668 VDPWR.n956 VDPWR.n955 0.15675
R1669 VDPWR.n955 VDPWR.n954 0.15675
R1670 VDPWR.n954 VDPWR.n295 0.15675
R1671 VDPWR.n296 VDPWR.n295 0.15675
R1672 VDPWR.n417 VDPWR.n296 0.15675
R1673 VDPWR.n418 VDPWR.n417 0.15675
R1674 VDPWR.n419 VDPWR.n418 0.15675
R1675 VDPWR.n420 VDPWR.n419 0.15675
R1676 VDPWR.n420 VDPWR.n415 0.15675
R1677 VDPWR.n424 VDPWR.n415 0.15675
R1678 VDPWR.n425 VDPWR.n424 0.15675
R1679 VDPWR.n426 VDPWR.n425 0.15675
R1680 VDPWR.n426 VDPWR.n413 0.15675
R1681 VDPWR.n444 VDPWR.n413 0.15675
R1682 VDPWR.n445 VDPWR.n444 0.15675
R1683 VDPWR.n446 VDPWR.n445 0.15675
R1684 VDPWR.n446 VDPWR.n411 0.15675
R1685 VDPWR.n464 VDPWR.n411 0.15675
R1686 VDPWR.n465 VDPWR.n464 0.15675
R1687 VDPWR.n465 VDPWR.n395 0.15675
R1688 VDPWR.n471 VDPWR.n395 0.15675
R1689 VDPWR.n472 VDPWR.n471 0.15675
R1690 VDPWR.n473 VDPWR.n472 0.15675
R1691 VDPWR.n473 VDPWR.n379 0.15675
R1692 VDPWR.n479 VDPWR.n379 0.15675
R1693 VDPWR.n480 VDPWR.n479 0.15675
R1694 VDPWR.n481 VDPWR.n480 0.15675
R1695 VDPWR.n481 VDPWR.n377 0.15675
R1696 VDPWR.n499 VDPWR.n377 0.15675
R1697 VDPWR.n500 VDPWR.n499 0.15675
R1698 VDPWR.n501 VDPWR.n500 0.15675
R1699 VDPWR.n501 VDPWR.n375 0.15675
R1700 VDPWR.n512 VDPWR.n375 0.15675
R1701 VDPWR.n515 VDPWR.n514 0.15675
R1702 VDPWR.n515 VDPWR.n373 0.15675
R1703 VDPWR.n533 VDPWR.n373 0.15675
R1704 VDPWR.n534 VDPWR.n533 0.15675
R1705 VDPWR.n535 VDPWR.n534 0.15675
R1706 VDPWR.n535 VDPWR.n371 0.15675
R1707 VDPWR.n539 VDPWR.n371 0.15675
R1708 VDPWR.n540 VDPWR.n539 0.15675
R1709 VDPWR.n187 VDPWR.n138 0.15675
R1710 VDPWR.n183 VDPWR.n138 0.15675
R1711 VDPWR.n183 VDPWR.n182 0.15675
R1712 VDPWR.n182 VDPWR.n181 0.15675
R1713 VDPWR.n290 VDPWR.n3 0.15675
R1714 VDPWR.n286 VDPWR.n3 0.15675
R1715 VDPWR.n286 VDPWR.n285 0.15675
R1716 VDPWR.n285 VDPWR.n284 0.15675
R1717 VDPWR.n284 VDPWR.n5 0.15675
R1718 VDPWR.n280 VDPWR.n5 0.15675
R1719 VDPWR.n280 VDPWR.n279 0.15675
R1720 VDPWR.n279 VDPWR.n278 0.15675
R1721 VDPWR.n278 VDPWR.n9 0.15675
R1722 VDPWR.n274 VDPWR.n9 0.15675
R1723 VDPWR.n274 VDPWR.n273 0.15675
R1724 VDPWR.n273 VDPWR.n12 0.15675
R1725 VDPWR.n269 VDPWR.n12 0.15675
R1726 VDPWR.n269 VDPWR.n268 0.15675
R1727 VDPWR.n268 VDPWR.n267 0.15675
R1728 VDPWR.n267 VDPWR.n14 0.15675
R1729 VDPWR.n263 VDPWR.n14 0.15675
R1730 VDPWR.n263 VDPWR.n262 0.15675
R1731 VDPWR.n262 VDPWR.n261 0.15675
R1732 VDPWR.n261 VDPWR.n17 0.15675
R1733 VDPWR.n257 VDPWR.n17 0.15675
R1734 VDPWR.n257 VDPWR.n256 0.15675
R1735 VDPWR.n256 VDPWR.n255 0.15675
R1736 VDPWR.n255 VDPWR.n19 0.15675
R1737 VDPWR.n43 VDPWR.n19 0.15675
R1738 VDPWR.n44 VDPWR.n43 0.15675
R1739 VDPWR.n45 VDPWR.n44 0.15675
R1740 VDPWR.n45 VDPWR.n39 0.15675
R1741 VDPWR.n50 VDPWR.n39 0.15675
R1742 VDPWR.n51 VDPWR.n50 0.15675
R1743 VDPWR.n52 VDPWR.n51 0.15675
R1744 VDPWR.n52 VDPWR.n36 0.15675
R1745 VDPWR.n36 VDPWR.n35 0.15675
R1746 VDPWR.n58 VDPWR.n35 0.15675
R1747 VDPWR.n59 VDPWR.n58 0.15675
R1748 VDPWR.n60 VDPWR.n59 0.15675
R1749 VDPWR.n60 VDPWR.n33 0.15675
R1750 VDPWR.n65 VDPWR.n33 0.15675
R1751 VDPWR.n66 VDPWR.n65 0.15675
R1752 VDPWR.n67 VDPWR.n66 0.15675
R1753 VDPWR.n67 VDPWR.n30 0.15675
R1754 VDPWR.n72 VDPWR.n30 0.15675
R1755 VDPWR.n73 VDPWR.n72 0.15675
R1756 VDPWR.n74 VDPWR.n73 0.15675
R1757 VDPWR.n74 VDPWR.n27 0.15675
R1758 VDPWR.n79 VDPWR.n27 0.15675
R1759 VDPWR.n80 VDPWR.n79 0.15675
R1760 VDPWR.n81 VDPWR.n80 0.15675
R1761 VDPWR.n81 VDPWR.n25 0.15675
R1762 VDPWR.n85 VDPWR.n25 0.15675
R1763 VDPWR.n86 VDPWR.n85 0.15675
R1764 VDPWR.n248 VDPWR.n86 0.15675
R1765 VDPWR.n248 VDPWR.n247 0.15675
R1766 VDPWR.n247 VDPWR.n246 0.15675
R1767 VDPWR.n246 VDPWR.n87 0.15675
R1768 VDPWR.n241 VDPWR.n87 0.15675
R1769 VDPWR.n241 VDPWR.n240 0.15675
R1770 VDPWR.n240 VDPWR.n239 0.15675
R1771 VDPWR.n239 VDPWR.n90 0.15675
R1772 VDPWR.n235 VDPWR.n90 0.15675
R1773 VDPWR.n235 VDPWR.n234 0.15675
R1774 VDPWR.n234 VDPWR.n233 0.15675
R1775 VDPWR.n233 VDPWR.n93 0.15675
R1776 VDPWR.n229 VDPWR.n93 0.15675
R1777 VDPWR.n229 VDPWR.n228 0.15675
R1778 VDPWR.n228 VDPWR.n227 0.15675
R1779 VDPWR.n227 VDPWR.n95 0.15675
R1780 VDPWR.n223 VDPWR.n95 0.15675
R1781 VDPWR.n223 VDPWR.n222 0.15675
R1782 VDPWR.n222 VDPWR.n98 0.15675
R1783 VDPWR.n218 VDPWR.n98 0.15675
R1784 VDPWR.n218 VDPWR.n217 0.15675
R1785 VDPWR.n217 VDPWR.n216 0.15675
R1786 VDPWR.n216 VDPWR.n101 0.15675
R1787 VDPWR.n212 VDPWR.n101 0.15675
R1788 VDPWR.n212 VDPWR.n211 0.15675
R1789 VDPWR.n211 VDPWR.n210 0.15675
R1790 VDPWR.n210 VDPWR.n103 0.15675
R1791 VDPWR.n113 VDPWR.n103 0.15675
R1792 VDPWR.n114 VDPWR.n113 0.15675
R1793 VDPWR.n119 VDPWR.n114 0.15675
R1794 VDPWR.n120 VDPWR.n119 0.15675
R1795 VDPWR.n121 VDPWR.n120 0.15675
R1796 VDPWR.n121 VDPWR.n111 0.15675
R1797 VDPWR.n126 VDPWR.n111 0.15675
R1798 VDPWR.n127 VDPWR.n126 0.15675
R1799 VDPWR.n128 VDPWR.n127 0.15675
R1800 VDPWR.n128 VDPWR.n109 0.15675
R1801 VDPWR.n132 VDPWR.n109 0.15675
R1802 VDPWR.n133 VDPWR.n132 0.15675
R1803 VDPWR.n202 VDPWR.n133 0.15675
R1804 VDPWR.n202 VDPWR.n201 0.15675
R1805 VDPWR.n201 VDPWR.n200 0.15675
R1806 VDPWR.n200 VDPWR.n134 0.15675
R1807 VDPWR.n195 VDPWR.n134 0.15675
R1808 VDPWR.n195 VDPWR.n194 0.15675
R1809 VDPWR.n194 VDPWR.n193 0.15675
R1810 VDPWR.t372 VDPWR.t120 0.137822
R1811 VDPWR.n544 VDPWR.t182 0.1368
R1812 VDPWR.n706 VDPWR.n606 0.131176
R1813 VDPWR.n569 VDPWR.n567 0.1255
R1814 VDPWR.n567 VDPWR.n565 0.1255
R1815 VDPWR.n565 VDPWR.n563 0.1255
R1816 VDPWR.n563 VDPWR.n561 0.1255
R1817 VDPWR.n561 VDPWR.n559 0.1255
R1818 VDPWR.n559 VDPWR.n557 0.1255
R1819 VDPWR.n557 VDPWR.n555 0.1255
R1820 VDPWR.n555 VDPWR.n551 0.1255
R1821 VDPWR.n578 VDPWR.n551 0.1255
R1822 VDPWR.n595 VDPWR.n594 0.1255
R1823 VDPWR.n594 VDPWR.n592 0.1255
R1824 VDPWR.n592 VDPWR.n590 0.1255
R1825 VDPWR.n590 VDPWR.n588 0.1255
R1826 VDPWR.n588 VDPWR.n586 0.1255
R1827 VDPWR.n586 VDPWR.n584 0.1255
R1828 VDPWR.n584 VDPWR.n582 0.1255
R1829 VDPWR.n582 VDPWR.n580 0.1255
R1830 VDPWR.n580 VDPWR.n547 0.1255
R1831 VDPWR.n604 VDPWR.n547 0.1255
R1832 VDPWR.n674 VDPWR.n673 0.100307
R1833 VDPWR.n703 VDPWR.n702 0.09425
R1834 VDPWR.n696 VDPWR.n695 0.09425
R1835 VDPWR.n689 VDPWR.n688 0.09425
R1836 VDPWR.n682 VDPWR.n681 0.09425
R1837 VDPWR.n675 VDPWR.n674 0.09425
R1838 VDPWR.n513 VDPWR.n512 0.078625
R1839 VDPWR.n514 VDPWR.n513 0.078625
R1840 VDPWR.n704 VDPWR.n606 0.063
R1841 VDPWR.n702 VDPWR.n701 0.063
R1842 VDPWR.n695 VDPWR.n694 0.063
R1843 VDPWR.n688 VDPWR.n687 0.063
R1844 VDPWR.n681 VDPWR.n680 0.063
R1845 VDPWR.n971 VDPWR.n965 0.01225
R1846 VDPWR.n969 VDPWR.n965 0.01225
R1847 VDPWR.n967 VDPWR.n1 0.0068649
R1848 VDPWR.n970 VDPWR.n966 0.0068649
R1849 VDPWR.n968 VDPWR.n963 0.0068649
R1850 VDPWR.n972 VDPWR.n0 0.0068649
R1851 VDPWR.n966 VDPWR.n964 0.0068649
R1852 VDPWR.n970 VDPWR.n968 0.0068649
R1853 VDPWR.n963 VDPWR.n0 0.0068649
R1854 VDPWR.n969 VDPWR.n1 0.0068649
R1855 VDPWR.n544 VDPWR.t185 0.00152174
R1856 a_19190_29050.n4 a_19190_29050.t30 363.909
R1857 a_19190_29050.n4 a_19190_29050.t36 351.974
R1858 a_19190_29050.n12 a_19190_29050.n4 299.252
R1859 a_19190_29050.n4 a_19190_29050.n5 299.25
R1860 a_19190_29050.n4 a_19190_29050.n7 299.25
R1861 a_19190_29050.n3 a_19190_29050.t6 242.968
R1862 a_19190_29050.n10 a_19190_29050.n8 200.477
R1863 a_19190_29050.n10 a_19190_29050.n9 199.727
R1864 a_19190_29050.n6 a_19190_29050.t17 194.809
R1865 a_19190_29050.n6 a_19190_29050.t13 194.809
R1866 a_19190_29050.n11 a_19190_29050.t11 194.809
R1867 a_19190_29050.n11 a_19190_29050.t34 194.809
R1868 a_19190_29050.n4 a_19190_29050.n6 163.097
R1869 a_19190_29050.n3 a_19190_29050.n11 161.653
R1870 a_19190_29050.n8 a_19190_29050.t3 48.0005
R1871 a_19190_29050.n8 a_19190_29050.t1 48.0005
R1872 a_19190_29050.n9 a_19190_29050.t7 48.0005
R1873 a_19190_29050.n9 a_19190_29050.t2 48.0005
R1874 a_19190_29050.n5 a_19190_29050.t9 39.4005
R1875 a_19190_29050.n5 a_19190_29050.t4 39.4005
R1876 a_19190_29050.n7 a_19190_29050.t10 39.4005
R1877 a_19190_29050.n7 a_19190_29050.t5 39.4005
R1878 a_19190_29050.n12 a_19190_29050.t8 39.4005
R1879 a_19190_29050.t0 a_19190_29050.n12 39.4005
R1880 a_19190_29050.n3 a_19190_29050.n10 5.2505
R1881 a_19190_29050.n0 a_19190_29050.t18 4.8248
R1882 a_19190_29050.n1 a_19190_29050.t12 4.5005
R1883 a_19190_29050.n1 a_19190_29050.t21 4.5005
R1884 a_19190_29050.n0 a_19190_29050.t27 4.5005
R1885 a_19190_29050.n0 a_19190_29050.t22 4.5005
R1886 a_19190_29050.n0 a_19190_29050.t29 4.5005
R1887 a_19190_29050.n0 a_19190_29050.t33 4.5005
R1888 a_19190_29050.n0 a_19190_29050.t15 4.5005
R1889 a_19190_29050.n0 a_19190_29050.t35 4.5005
R1890 a_19190_29050.n1 a_19190_29050.t25 4.5005
R1891 a_19190_29050.n1 a_19190_29050.t19 4.5005
R1892 a_19190_29050.n1 a_19190_29050.t20 4.5005
R1893 a_19190_29050.n1 a_19190_29050.t26 4.5005
R1894 a_19190_29050.n1 a_19190_29050.t31 4.5005
R1895 a_19190_29050.n2 a_19190_29050.t28 4.5005
R1896 a_19190_29050.n2 a_19190_29050.t32 4.5005
R1897 a_19190_29050.n2 a_19190_29050.t14 4.5005
R1898 a_19190_29050.n2 a_19190_29050.t23 4.5005
R1899 a_19190_29050.n2 a_19190_29050.t16 4.5005
R1900 a_19190_29050.n2 a_19190_29050.t24 4.5005
R1901 a_19190_29050.n4 a_19190_29050.n2 11.6632
R1902 a_19190_29050.n2 a_19190_29050.n1 3.5678
R1903 a_19190_29050.n4 a_19190_29050.n3 2.7106
R1904 a_19190_29050.n1 a_19190_29050.n0 2.3035
R1905 a_14348_27710.n2 a_14348_27710.t27 355.784
R1906 a_14348_27710.n8 a_14348_27710.t42 355.502
R1907 a_14348_27710.n10 a_14348_27710.t48 354.75
R1908 a_14348_27710.n0 a_14348_27710.t37 351.002
R1909 a_14348_27710.n2 a_14348_27710.t28 310.401
R1910 a_14348_27710.n3 a_14348_27710.t15 310.401
R1911 a_14348_27710.n4 a_14348_27710.t16 310.401
R1912 a_14348_27710.n5 a_14348_27710.t18 310.401
R1913 a_14348_27710.n6 a_14348_27710.t19 310.401
R1914 a_14348_27710.n7 a_14348_27710.t20 310.401
R1915 a_14348_27710.n14 a_14348_27710.t39 310.401
R1916 a_14348_27710.n13 a_14348_27710.t40 310.401
R1917 a_14348_27710.n12 a_14348_27710.t33 310.401
R1918 a_14348_27710.n11 a_14348_27710.t46 310.401
R1919 a_14348_27710.n10 a_14348_27710.t47 310.401
R1920 a_14348_27710.n27 a_14348_27710.n26 306.808
R1921 a_14348_27710.n1 a_14348_27710.t38 305.901
R1922 a_14348_27710.n20 a_14348_27710.n19 301.933
R1923 a_14348_27710.n22 a_14348_27710.n21 301.933
R1924 a_14348_27710.n24 a_14348_27710.n23 301.933
R1925 a_14348_27710.n29 a_14348_27710.n28 297.433
R1926 a_14348_27710.n27 a_14348_27710.n25 297.433
R1927 a_14348_27710.t0 a_14348_27710.n50 149.127
R1928 a_14348_27710.n18 a_14348_27710.t9 98.9207
R1929 a_14348_27710.n28 a_14348_27710.t5 39.4005
R1930 a_14348_27710.n28 a_14348_27710.t11 39.4005
R1931 a_14348_27710.n26 a_14348_27710.t12 39.4005
R1932 a_14348_27710.n26 a_14348_27710.t1 39.4005
R1933 a_14348_27710.n25 a_14348_27710.t2 39.4005
R1934 a_14348_27710.n25 a_14348_27710.t10 39.4005
R1935 a_14348_27710.n19 a_14348_27710.t13 39.4005
R1936 a_14348_27710.n19 a_14348_27710.t3 39.4005
R1937 a_14348_27710.n21 a_14348_27710.t6 39.4005
R1938 a_14348_27710.n21 a_14348_27710.t7 39.4005
R1939 a_14348_27710.n23 a_14348_27710.t8 39.4005
R1940 a_14348_27710.n23 a_14348_27710.t4 39.4005
R1941 a_14348_27710.n50 a_14348_27710.n30 13.563
R1942 a_14348_27710.n50 a_14348_27710.n49 12.3446
R1943 a_14348_27710.n20 a_14348_27710.n18 4.90675
R1944 a_14348_27710.n31 a_14348_27710.t23 4.8248
R1945 a_14348_27710.n38 a_14348_27710.t44 4.5005
R1946 a_14348_27710.n37 a_14348_27710.t25 4.5005
R1947 a_14348_27710.n36 a_14348_27710.t31 4.5005
R1948 a_14348_27710.n35 a_14348_27710.t26 4.5005
R1949 a_14348_27710.n34 a_14348_27710.t32 4.5005
R1950 a_14348_27710.n33 a_14348_27710.t41 4.5005
R1951 a_14348_27710.n32 a_14348_27710.t22 4.5005
R1952 a_14348_27710.n31 a_14348_27710.t43 4.5005
R1953 a_14348_27710.n40 a_14348_27710.t14 4.5005
R1954 a_14348_27710.n39 a_14348_27710.t24 4.5005
R1955 a_14348_27710.n41 a_14348_27710.t36 4.5005
R1956 a_14348_27710.n42 a_14348_27710.t17 4.5005
R1957 a_14348_27710.n43 a_14348_27710.t29 4.5005
R1958 a_14348_27710.n44 a_14348_27710.t21 4.5005
R1959 a_14348_27710.n45 a_14348_27710.t30 4.5005
R1960 a_14348_27710.n46 a_14348_27710.t34 4.5005
R1961 a_14348_27710.n47 a_14348_27710.t45 4.5005
R1962 a_14348_27710.n48 a_14348_27710.t35 4.5005
R1963 a_14348_27710.n49 a_14348_27710.t49 4.5005
R1964 a_14348_27710.n15 a_14348_27710.n1 4.5005
R1965 a_14348_27710.n9 a_14348_27710.n0 4.5005
R1966 a_14348_27710.n17 a_14348_27710.n16 4.5005
R1967 a_14348_27710.n30 a_14348_27710.n29 4.5005
R1968 a_14348_27710.n29 a_14348_27710.n27 1.59425
R1969 a_14348_27710.n18 a_14348_27710.n17 1.28175
R1970 a_14348_27710.n22 a_14348_27710.n20 1.1255
R1971 a_14348_27710.n24 a_14348_27710.n22 1.1255
R1972 a_14348_27710.n30 a_14348_27710.n24 1.1255
R1973 a_14348_27710.n32 a_14348_27710.n31 0.3295
R1974 a_14348_27710.n33 a_14348_27710.n32 0.3295
R1975 a_14348_27710.n34 a_14348_27710.n33 0.3295
R1976 a_14348_27710.n35 a_14348_27710.n34 0.3295
R1977 a_14348_27710.n36 a_14348_27710.n35 0.3295
R1978 a_14348_27710.n37 a_14348_27710.n36 0.3295
R1979 a_14348_27710.n38 a_14348_27710.n37 0.3295
R1980 a_14348_27710.n40 a_14348_27710.n39 0.3295
R1981 a_14348_27710.n48 a_14348_27710.n47 0.3295
R1982 a_14348_27710.n47 a_14348_27710.n46 0.3295
R1983 a_14348_27710.n46 a_14348_27710.n45 0.3295
R1984 a_14348_27710.n45 a_14348_27710.n44 0.3295
R1985 a_14348_27710.n44 a_14348_27710.n43 0.3295
R1986 a_14348_27710.n43 a_14348_27710.n42 0.3295
R1987 a_14348_27710.n42 a_14348_27710.n41 0.3295
R1988 a_14348_27710.n49 a_14348_27710.n48 0.3248
R1989 a_14348_27710.n39 a_14348_27710.n38 0.306
R1990 a_14348_27710.n41 a_14348_27710.n40 0.306
R1991 a_14348_27710.n3 a_14348_27710.n2 0.28175
R1992 a_14348_27710.n4 a_14348_27710.n3 0.28175
R1993 a_14348_27710.n5 a_14348_27710.n4 0.28175
R1994 a_14348_27710.n6 a_14348_27710.n5 0.28175
R1995 a_14348_27710.n7 a_14348_27710.n6 0.28175
R1996 a_14348_27710.n8 a_14348_27710.n7 0.28175
R1997 a_14348_27710.n9 a_14348_27710.n8 0.28175
R1998 a_14348_27710.n15 a_14348_27710.n14 0.28175
R1999 a_14348_27710.n14 a_14348_27710.n13 0.28175
R2000 a_14348_27710.n13 a_14348_27710.n12 0.28175
R2001 a_14348_27710.n12 a_14348_27710.n11 0.28175
R2002 a_14348_27710.n11 a_14348_27710.n10 0.28175
R2003 a_14348_27710.n16 a_14348_27710.n9 0.141125
R2004 a_14348_27710.n16 a_14348_27710.n15 0.141125
R2005 a_14348_27710.n17 a_14348_27710.n0 0.078625
R2006 a_14348_27710.n17 a_14348_27710.n1 0.078625
R2007 a_19190_31610.n15 a_19190_31610.t20 310.488
R2008 a_19190_31610.n1 a_19190_31610.t21 310.488
R2009 a_19190_31610.n6 a_19190_31610.t17 310.488
R2010 a_19190_31610.n4 a_19190_31610.n0 297.433
R2011 a_19190_31610.n9 a_19190_31610.n5 297.433
R2012 a_19190_31610.n19 a_19190_31610.n18 297.433
R2013 a_19190_31610.n13 a_19190_31610.t16 248.133
R2014 a_19190_31610.n13 a_19190_31610.n12 199.383
R2015 a_19190_31610.n14 a_19190_31610.n11 194.883
R2016 a_19190_31610.n17 a_19190_31610.t11 184.097
R2017 a_19190_31610.n3 a_19190_31610.t7 184.097
R2018 a_19190_31610.n8 a_19190_31610.t3 184.097
R2019 a_19190_31610.n16 a_19190_31610.n15 167.094
R2020 a_19190_31610.n2 a_19190_31610.n1 167.094
R2021 a_19190_31610.n7 a_19190_31610.n6 167.094
R2022 a_19190_31610.n18 a_19190_31610.n17 161.3
R2023 a_19190_31610.n4 a_19190_31610.n3 161.3
R2024 a_19190_31610.n9 a_19190_31610.n8 161.3
R2025 a_19190_31610.n16 a_19190_31610.t13 120.501
R2026 a_19190_31610.n15 a_19190_31610.t19 120.501
R2027 a_19190_31610.n2 a_19190_31610.t9 120.501
R2028 a_19190_31610.n1 a_19190_31610.t22 120.501
R2029 a_19190_31610.n7 a_19190_31610.t5 120.501
R2030 a_19190_31610.n6 a_19190_31610.t18 120.501
R2031 a_19190_31610.n12 a_19190_31610.t15 48.0005
R2032 a_19190_31610.n12 a_19190_31610.t0 48.0005
R2033 a_19190_31610.n11 a_19190_31610.t2 48.0005
R2034 a_19190_31610.n11 a_19190_31610.t1 48.0005
R2035 a_19190_31610.n17 a_19190_31610.n16 40.7027
R2036 a_19190_31610.n3 a_19190_31610.n2 40.7027
R2037 a_19190_31610.n8 a_19190_31610.n7 40.7027
R2038 a_19190_31610.n0 a_19190_31610.t8 39.4005
R2039 a_19190_31610.n0 a_19190_31610.t10 39.4005
R2040 a_19190_31610.n5 a_19190_31610.t4 39.4005
R2041 a_19190_31610.n5 a_19190_31610.t6 39.4005
R2042 a_19190_31610.n19 a_19190_31610.t12 39.4005
R2043 a_19190_31610.t14 a_19190_31610.n19 39.4005
R2044 a_19190_31610.n10 a_19190_31610.n4 6.6255
R2045 a_19190_31610.n10 a_19190_31610.n9 6.6255
R2046 a_19190_31610.n14 a_19190_31610.n13 5.2505
R2047 a_19190_31610.n18 a_19190_31610.n10 4.5005
R2048 a_19190_31610.n18 a_19190_31610.n14 0.78175
R2049 a_19190_31850.n9 a_19190_31850.t25 362.342
R2050 a_19190_31850.n23 a_19190_31850.t32 355.094
R2051 a_19190_31850.n11 a_19190_31850.n10 302.183
R2052 a_19190_31850.n20 a_19190_31850.n19 302.183
R2053 a_19190_31850.n24 a_19190_31850.n23 302.183
R2054 a_19190_31850.n16 a_19190_31850.t1 242.968
R2055 a_19190_31850.n15 a_19190_31850.n13 200.477
R2056 a_19190_31850.n15 a_19190_31850.n14 199.727
R2057 a_19190_31850.n12 a_19190_31850.t19 194.809
R2058 a_19190_31850.n12 a_19190_31850.t17 194.809
R2059 a_19190_31850.n21 a_19190_31850.t12 194.809
R2060 a_19190_31850.n21 a_19190_31850.t11 194.809
R2061 a_19190_31850.n22 a_19190_31850.n21 166.03
R2062 a_19190_31850.n17 a_19190_31850.n12 161.53
R2063 a_19190_31850.n14 a_19190_31850.t2 48.0005
R2064 a_19190_31850.n14 a_19190_31850.t0 48.0005
R2065 a_19190_31850.n13 a_19190_31850.t3 48.0005
R2066 a_19190_31850.n13 a_19190_31850.t4 48.0005
R2067 a_19190_31850.n9 a_19190_31850.n8 40.0791
R2068 a_19190_31850.n10 a_19190_31850.t5 39.4005
R2069 a_19190_31850.n10 a_19190_31850.t6 39.4005
R2070 a_19190_31850.n19 a_19190_31850.t8 39.4005
R2071 a_19190_31850.n19 a_19190_31850.t7 39.4005
R2072 a_19190_31850.n24 a_19190_31850.t9 39.4005
R2073 a_19190_31850.t10 a_19190_31850.n24 39.4005
R2074 a_19190_31850.n16 a_19190_31850.n15 5.2505
R2075 a_19190_31850.n0 a_19190_31850.t23 4.8248
R2076 a_19190_31850.n3 a_19190_31850.t18 4.5005
R2077 a_19190_31850.n3 a_19190_31850.t27 4.5005
R2078 a_19190_31850.n2 a_19190_31850.t34 4.5005
R2079 a_19190_31850.n2 a_19190_31850.t28 4.5005
R2080 a_19190_31850.n1 a_19190_31850.t36 4.5005
R2081 a_19190_31850.n1 a_19190_31850.t15 4.5005
R2082 a_19190_31850.n0 a_19190_31850.t21 4.5005
R2083 a_19190_31850.n0 a_19190_31850.t16 4.5005
R2084 a_19190_31850.n7 a_19190_31850.t31 4.5005
R2085 a_19190_31850.n3 a_19190_31850.t24 4.5005
R2086 a_19190_31850.n7 a_19190_31850.t26 4.5005
R2087 a_19190_31850.n6 a_19190_31850.t33 4.5005
R2088 a_19190_31850.n6 a_19190_31850.t13 4.5005
R2089 a_19190_31850.n4 a_19190_31850.t35 4.5005
R2090 a_19190_31850.n4 a_19190_31850.t14 4.5005
R2091 a_19190_31850.n5 a_19190_31850.t20 4.5005
R2092 a_19190_31850.n5 a_19190_31850.t29 4.5005
R2093 a_19190_31850.n8 a_19190_31850.t22 4.5005
R2094 a_19190_31850.n8 a_19190_31850.t30 4.5005
R2095 a_19190_31850.n18 a_19190_31850.n17 4.5005
R2096 a_19190_31850.n11 a_19190_31850.n9 2.93757
R2097 a_19190_31850.n1 a_19190_31850.n0 0.9875
R2098 a_19190_31850.n8 a_19190_31850.n5 0.9828
R2099 a_19190_31850.n20 a_19190_31850.n18 0.7505
R2100 a_19190_31850.n23 a_19190_31850.n22 0.7505
R2101 a_19190_31850.n4 a_19190_31850.n6 0.6585
R2102 a_19190_31850.n5 a_19190_31850.n4 0.6585
R2103 a_19190_31850.n3 a_19190_31850.n2 0.6585
R2104 a_19190_31850.n2 a_19190_31850.n1 0.6585
R2105 a_19190_31850.n6 a_19190_31850.n7 0.635
R2106 a_19190_31850.n7 a_19190_31850.n3 0.635
R2107 a_19190_31850.n17 a_19190_31850.n16 0.422375
R2108 a_19190_31850.n18 a_19190_31850.n11 0.3755
R2109 a_19190_31850.n22 a_19190_31850.n20 0.3755
R2110 a_26300_25010.n5 a_26300_25010.t0 758.734
R2111 a_26300_25010.n4 a_26300_25010.t2 758.734
R2112 a_26300_25010.n0 a_26300_25010.t5 538.234
R2113 a_26300_25010.n3 a_26300_25010.n2 342.757
R2114 a_26300_25010.t1 a_26300_25010.n5 260.733
R2115 a_26300_25010.n3 a_26300_25010.t7 190.123
R2116 a_26300_25010.n4 a_26300_25010.n3 180.8
R2117 a_26300_25010.n0 a_26300_25010.t6 136.567
R2118 a_26300_25010.n1 a_26300_25010.t4 136.567
R2119 a_26300_25010.n2 a_26300_25010.t3 136.567
R2120 a_26300_25010.n1 a_26300_25010.n0 128.534
R2121 a_26300_25010.n2 a_26300_25010.n1 128.534
R2122 a_26300_25010.n5 a_26300_25010.n4 57.6005
R2123 a_26300_25670.n2 a_26300_25670.t0 755.889
R2124 a_26300_25670.n1 a_26300_25670.t4 343.034
R2125 a_26300_25670.t1 a_26300_25670.n2 270.334
R2126 a_26300_25670.n1 a_26300_25670.n0 212.733
R2127 a_26300_25670.n0 a_26300_25670.t2 48.0005
R2128 a_26300_25670.n0 a_26300_25670.t3 48.0005
R2129 a_26300_25670.n2 a_26300_25670.n1 35.2005
R2130 w_13193_29093.n2697 w_13193_29093.n2696 1.86032e+06
R2131 w_13193_29093.n2535 w_13193_29093.n2534 589600
R2132 w_13193_29093.n2696 w_13193_29093.n65 533500
R2133 w_13193_29093.n2534 w_13193_29093.n65 478500
R2134 w_13193_29093.n2442 w_13193_29093.n2441 312538
R2135 w_13193_29093.n2698 w_13193_29093.n65 286825
R2136 w_13193_29093.n2223 w_13193_29093.n61 263120
R2137 w_13193_29093.n2704 w_13193_29093.n2703 206882
R2138 w_13193_29093.n2439 w_13193_29093.n2223 132880
R2139 w_13193_29093.n2440 w_13193_29093.n0 112733
R2140 w_13193_29093.n2388 w_13193_29093.n61 88572
R2141 w_13193_29093.n2704 w_13193_29093.n60 74541.2
R2142 w_13193_29093.n2698 w_13193_29093.n2697 39524.8
R2143 w_13193_29093.t245 w_13193_29093.n2698 27530.6
R2144 w_13193_29093.n2445 w_13193_29093.n2442 24406.2
R2145 w_13193_29093.n2702 w_13193_29093.n2701 19915.8
R2146 w_13193_29093.n2443 w_13193_29093.n60 11768.9
R2147 w_13193_29093.n2441 w_13193_29093.n60 11350.7
R2148 w_13193_29093.n2441 w_13193_29093.n2440 7867.26
R2149 w_13193_29093.n2703 w_13193_29093.n2702 6049.26
R2150 w_13193_29093.n2699 w_13193_29093.n64 5433.26
R2151 w_13193_29093.n2702 w_13193_29093.n63 5222.9
R2152 w_13193_29093.n2442 w_13193_29093.n2221 4738.46
R2153 w_13193_29093.n2216 w_13193_29093.n62 4546.97
R2154 w_13193_29093.n2443 w_13193_29093.n62 4456.9
R2155 w_13193_29093.n2444 w_13193_29093.n2443 4150.65
R2156 w_13193_29093.n60 w_13193_29093.n0 3685.42
R2157 w_13193_29093.t31 w_13193_29093.n64 3396.4
R2158 w_13193_29093.n2444 w_13193_29093.n2216 3257.69
R2159 w_13193_29093.t53 w_13193_29093.t214 2857.38
R2160 w_13193_29093.n2703 w_13193_29093.n62 2550.86
R2161 w_13193_29093.n2764 w_13193_29093.n2763 2401.67
R2162 w_13193_29093.n2765 w_13193_29093.t5 2346.67
R2163 w_13193_29093.n2703 w_13193_29093.n61 1998.47
R2164 w_13193_29093.n2701 w_13193_29093.n2700 1910.53
R2165 w_13193_29093.t233 w_13193_29093.t208 1751.46
R2166 w_13193_29093.n2440 w_13193_29093.n2222 1452.43
R2167 w_13193_29093.n2699 w_13193_29093.t245 1444.58
R2168 w_13193_29093.n2445 w_13193_29093.n2444 1337.98
R2169 w_13193_29093.n1920 w_13193_29093.n321 1214.72
R2170 w_13193_29093.n326 w_13193_29093.n321 1214.72
R2171 w_13193_29093.n1913 w_13193_29093.n326 1214.72
R2172 w_13193_29093.n1913 w_13193_29093.n1912 1214.72
R2173 w_13193_29093.n1912 w_13193_29093.n1 1214.72
R2174 w_13193_29093.n364 w_13193_29093.n2 1214.72
R2175 w_13193_29093.n379 w_13193_29093.n364 1214.72
R2176 w_13193_29093.n379 w_13193_29093.n355 1214.72
R2177 w_13193_29093.n1842 w_13193_29093.n355 1214.72
R2178 w_13193_29093.n1842 w_13193_29093.n3 1214.72
R2179 w_13193_29093.n1386 w_13193_29093.n612 1214.72
R2180 w_13193_29093.n1465 w_13193_29093.n612 1214.72
R2181 w_13193_29093.n1465 w_13193_29093.n607 1214.72
R2182 w_13193_29093.n1474 w_13193_29093.n607 1214.72
R2183 w_13193_29093.n1474 w_13193_29093.n4 1214.72
R2184 w_13193_29093.n594 w_13193_29093.n5 1214.72
R2185 w_13193_29093.n1489 w_13193_29093.n594 1214.72
R2186 w_13193_29093.n1489 w_13193_29093.n589 1214.72
R2187 w_13193_29093.n1496 w_13193_29093.n589 1214.72
R2188 w_13193_29093.n1496 w_13193_29093.n6 1214.72
R2189 w_13193_29093.n1655 w_13193_29093.n489 1214.72
R2190 w_13193_29093.n1662 w_13193_29093.n489 1214.72
R2191 w_13193_29093.n1662 w_13193_29093.n473 1214.72
R2192 w_13193_29093.n1675 w_13193_29093.n473 1214.72
R2193 w_13193_29093.n1675 w_13193_29093.n7 1214.72
R2194 w_13193_29093.n468 w_13193_29093.n8 1214.72
R2195 w_13193_29093.n1684 w_13193_29093.n468 1214.72
R2196 w_13193_29093.n1684 w_13193_29093.n457 1214.72
R2197 w_13193_29093.n1717 w_13193_29093.n457 1214.72
R2198 w_13193_29093.n1717 w_13193_29093.n9 1214.72
R2199 w_13193_29093.n1589 w_13193_29093.n492 1214.72
R2200 w_13193_29093.n1583 w_13193_29093.n492 1214.72
R2201 w_13193_29093.n1583 w_13193_29093.n1582 1214.72
R2202 w_13193_29093.n1582 w_13193_29093.n1581 1214.72
R2203 w_13193_29093.n1581 w_13193_29093.n10 1214.72
R2204 w_13193_29093.n1574 w_13193_29093.n11 1214.72
R2205 w_13193_29093.n1574 w_13193_29093.n1573 1214.72
R2206 w_13193_29093.n1573 w_13193_29093.n449 1214.72
R2207 w_13193_29093.n1748 w_13193_29093.n449 1214.72
R2208 w_13193_29093.n1748 w_13193_29093.n12 1214.72
R2209 w_13193_29093.n2637 w_13193_29093.n159 1210.53
R2210 w_13193_29093.n2533 w_13193_29093.n171 1210.53
R2211 w_13193_29093.n2531 w_13193_29093.n183 1210.53
R2212 w_13193_29093.t4 w_13193_29093.n2708 1186
R2213 w_13193_29093.t4 w_13193_29093.n2716 1186
R2214 w_13193_29093.n2717 w_13193_29093.t4 1186
R2215 w_13193_29093.n2722 w_13193_29093.n2721 1186
R2216 w_13193_29093.n2693 w_13193_29093.n2692 1182.8
R2217 w_13193_29093.n2376 w_13193_29093.n147 1182.8
R2218 w_13193_29093.n2548 w_13193_29093.n2547 1173.78
R2219 w_13193_29093.n2551 w_13193_29093.n2550 1173.78
R2220 w_13193_29093.n2542 w_13193_29093.n2541 1173.78
R2221 w_13193_29093.n201 w_13193_29093.n64 1170
R2222 w_13193_29093.n2223 w_13193_29093.n2221 1110.68
R2223 w_13193_29093.t193 w_13193_29093.t150 974.047
R2224 w_13193_29093.t53 w_13193_29093.t5 932.106
R2225 w_13193_29093.n2278 w_13193_29093.t128 833.01
R2226 w_13193_29093.n2279 w_13193_29093.t50 833.01
R2227 w_13193_29093.t261 w_13193_29093.t176 808.649
R2228 w_13193_29093.n2439 w_13193_29093.n2438 807.577
R2229 w_13193_29093.n2461 w_13193_29093.t146 789.313
R2230 w_13193_29093.t39 w_13193_29093.t33 784.865
R2231 w_13193_29093.n2547 w_13193_29093.t313 728.524
R2232 w_13193_29093.n2550 w_13193_29093.t317 728.524
R2233 w_13193_29093.n2541 w_13193_29093.t314 728.524
R2234 w_13193_29093.t53 w_13193_29093.n30 704.505
R2235 w_13193_29093.n2537 w_13193_29093.n2536 686.717
R2236 w_13193_29093.n2543 w_13193_29093.n197 686.717
R2237 w_13193_29093.n2553 w_13193_29093.n2552 686.717
R2238 w_13193_29093.n761 w_13193_29093.n760 686.717
R2239 w_13193_29093.n769 w_13193_29093.n768 686.717
R2240 w_13193_29093.n248 w_13193_29093.n247 686.717
R2241 w_13193_29093.n257 w_13193_29093.n256 686.717
R2242 w_13193_29093.n261 w_13193_29093.n259 686.717
R2243 w_13193_29093.n262 w_13193_29093.n261 686.717
R2244 w_13193_29093.n2552 w_13193_29093.n203 686.717
R2245 w_13193_29093.n2545 w_13193_29093.n2543 686.717
R2246 w_13193_29093.n2539 w_13193_29093.n2536 686.717
R2247 w_13193_29093.n2386 w_13193_29093.n2385 673.669
R2248 w_13193_29093.n2529 w_13193_29093.n2528 673.669
R2249 w_13193_29093.t168 w_13193_29093.n2216 671.756
R2250 w_13193_29093.n227 w_13193_29093.n226 669.307
R2251 w_13193_29093.n2499 w_13193_29093.n206 669.307
R2252 w_13193_29093.n748 w_13193_29093.n745 669.307
R2253 w_13193_29093.n1081 w_13193_29093.n1080 669.307
R2254 w_13193_29093.n2524 w_13193_29093.n207 669.307
R2255 w_13193_29093.n2506 w_13193_29093.n205 669.307
R2256 w_13193_29093.n233 w_13193_29093.n232 669.307
R2257 w_13193_29093.n2381 w_13193_29093.n2377 669.307
R2258 w_13193_29093.n2204 w_13193_29093.n2203 654.972
R2259 w_13193_29093.t53 w_13193_29093.n2 634.356
R2260 w_13193_29093.t53 w_13193_29093.n5 634.356
R2261 w_13193_29093.t53 w_13193_29093.n8 634.356
R2262 w_13193_29093.t53 w_13193_29093.n11 634.356
R2263 w_13193_29093.n2446 w_13193_29093.n2445 621.375
R2264 w_13193_29093.t230 w_13193_29093.t308 616.66
R2265 w_13193_29093.n2277 w_13193_29093.n2276 598.058
R2266 w_13193_29093.n2709 w_13193_29093.n32 589.889
R2267 w_13193_29093.n2762 w_13193_29093.n2761 589.889
R2268 w_13193_29093.n2260 w_13193_29093.n2259 585.003
R2269 w_13193_29093.n2436 w_13193_29093.n2225 585.003
R2270 w_13193_29093.n2390 w_13193_29093.n2389 585.001
R2271 w_13193_29093.n2375 w_13193_29093.n2371 585.001
R2272 w_13193_29093.n2366 w_13193_29093.n68 585.001
R2273 w_13193_29093.n2694 w_13193_29093.n67 585.001
R2274 w_13193_29093.n2695 w_13193_29093.n66 585.001
R2275 w_13193_29093.n2434 w_13193_29093.n2433 585.001
R2276 w_13193_29093.n2435 w_13193_29093.n2226 585.001
R2277 w_13193_29093.n2437 w_13193_29093.n2224 585.001
R2278 w_13193_29093.n2462 w_13193_29093.n2461 585.001
R2279 w_13193_29093.n2460 w_13193_29093.n2459 585.001
R2280 w_13193_29093.n2447 w_13193_29093.n2446 585.001
R2281 w_13193_29093.n2280 w_13193_29093.n2279 585.001
R2282 w_13193_29093.n2278 w_13193_29093.n2273 585.001
R2283 w_13193_29093.n2277 w_13193_29093.n2270 585.001
R2284 w_13193_29093.n2276 w_13193_29093.n2266 585.001
R2285 w_13193_29093.n2252 w_13193_29093.n2222 585.001
R2286 w_13193_29093.n1388 w_13193_29093.n1387 585
R2287 w_13193_29093.n1387 w_13193_29093.n1386 585
R2288 w_13193_29093.n1389 w_13193_29093.n613 585
R2289 w_13193_29093.n613 w_13193_29093.n612 585
R2290 w_13193_29093.n1464 w_13193_29093.n1463 585
R2291 w_13193_29093.n1465 w_13193_29093.n1464 585
R2292 w_13193_29093.n615 w_13193_29093.n604 585
R2293 w_13193_29093.n607 w_13193_29093.n604 585
R2294 w_13193_29093.n1475 w_13193_29093.n606 585
R2295 w_13193_29093.n1475 w_13193_29093.n1474 585
R2296 w_13193_29093.n1476 w_13193_29093.n603 585
R2297 w_13193_29093.n1476 w_13193_29093.n4 585
R2298 w_13193_29093.n1478 w_13193_29093.n1477 585
R2299 w_13193_29093.n1477 w_13193_29093.n5 585
R2300 w_13193_29093.n600 w_13193_29093.n595 585
R2301 w_13193_29093.n595 w_13193_29093.n594 585
R2302 w_13193_29093.n1488 w_13193_29093.n1487 585
R2303 w_13193_29093.n1489 w_13193_29093.n1488 585
R2304 w_13193_29093.n597 w_13193_29093.n587 585
R2305 w_13193_29093.n589 w_13193_29093.n587 585
R2306 w_13193_29093.n1497 w_13193_29093.n588 585
R2307 w_13193_29093.n1497 w_13193_29093.n1496 585
R2308 w_13193_29093.n1498 w_13193_29093.n582 585
R2309 w_13193_29093.n1498 w_13193_29093.n6 585
R2310 w_13193_29093.n1493 w_13193_29093.n591 585
R2311 w_13193_29093.n591 w_13193_29093.n6 585
R2312 w_13193_29093.n1495 w_13193_29093.n1494 585
R2313 w_13193_29093.n1496 w_13193_29093.n1495 585
R2314 w_13193_29093.n1492 w_13193_29093.n590 585
R2315 w_13193_29093.n590 w_13193_29093.n589 585
R2316 w_13193_29093.n1491 w_13193_29093.n1490 585
R2317 w_13193_29093.n1490 w_13193_29093.n1489 585
R2318 w_13193_29093.n593 w_13193_29093.n592 585
R2319 w_13193_29093.n594 w_13193_29093.n593 585
R2320 w_13193_29093.n1470 w_13193_29093.n1469 585
R2321 w_13193_29093.n1469 w_13193_29093.n5 585
R2322 w_13193_29093.n1471 w_13193_29093.n609 585
R2323 w_13193_29093.n609 w_13193_29093.n4 585
R2324 w_13193_29093.n1473 w_13193_29093.n1472 585
R2325 w_13193_29093.n1474 w_13193_29093.n1473 585
R2326 w_13193_29093.n1468 w_13193_29093.n608 585
R2327 w_13193_29093.n608 w_13193_29093.n607 585
R2328 w_13193_29093.n1467 w_13193_29093.n1466 585
R2329 w_13193_29093.n1466 w_13193_29093.n1465 585
R2330 w_13193_29093.n611 w_13193_29093.n610 585
R2331 w_13193_29093.n612 w_13193_29093.n611 585
R2332 w_13193_29093.n1385 w_13193_29093.n1384 585
R2333 w_13193_29093.n1386 w_13193_29093.n1385 585
R2334 w_13193_29093.n1720 w_13193_29093.n1719 585
R2335 w_13193_29093.n1719 w_13193_29093.n9 585
R2336 w_13193_29093.n1718 w_13193_29093.n455 585
R2337 w_13193_29093.n1718 w_13193_29093.n1717 585
R2338 w_13193_29093.n1681 w_13193_29093.n456 585
R2339 w_13193_29093.n457 w_13193_29093.n456 585
R2340 w_13193_29093.n1683 w_13193_29093.n1682 585
R2341 w_13193_29093.n1684 w_13193_29093.n1683 585
R2342 w_13193_29093.n1680 w_13193_29093.n469 585
R2343 w_13193_29093.n469 w_13193_29093.n468 585
R2344 w_13193_29093.n1679 w_13193_29093.n1678 585
R2345 w_13193_29093.n1678 w_13193_29093.n8 585
R2346 w_13193_29093.n1677 w_13193_29093.n470 585
R2347 w_13193_29093.n1677 w_13193_29093.n7 585
R2348 w_13193_29093.n1676 w_13193_29093.n472 585
R2349 w_13193_29093.n1676 w_13193_29093.n1675 585
R2350 w_13193_29093.n1659 w_13193_29093.n471 585
R2351 w_13193_29093.n473 w_13193_29093.n471 585
R2352 w_13193_29093.n1661 w_13193_29093.n1660 585
R2353 w_13193_29093.n1662 w_13193_29093.n1661 585
R2354 w_13193_29093.n1658 w_13193_29093.n1657 585
R2355 w_13193_29093.n1657 w_13193_29093.n489 585
R2356 w_13193_29093.n1656 w_13193_29093.n384 585
R2357 w_13193_29093.n1656 w_13193_29093.n1655 585
R2358 w_13193_29093.n1750 w_13193_29093.n446 585
R2359 w_13193_29093.n1750 w_13193_29093.n12 585
R2360 w_13193_29093.n1749 w_13193_29093.n448 585
R2361 w_13193_29093.n1749 w_13193_29093.n1748 585
R2362 w_13193_29093.n503 w_13193_29093.n447 585
R2363 w_13193_29093.n449 w_13193_29093.n447 585
R2364 w_13193_29093.n505 w_13193_29093.n504 585
R2365 w_13193_29093.n1573 w_13193_29093.n505 585
R2366 w_13193_29093.n1575 w_13193_29093.n502 585
R2367 w_13193_29093.n1575 w_13193_29093.n1574 585
R2368 w_13193_29093.n1577 w_13193_29093.n1576 585
R2369 w_13193_29093.n1576 w_13193_29093.n11 585
R2370 w_13193_29093.n1578 w_13193_29093.n501 585
R2371 w_13193_29093.n501 w_13193_29093.n10 585
R2372 w_13193_29093.n1580 w_13193_29093.n1579 585
R2373 w_13193_29093.n1581 w_13193_29093.n1580 585
R2374 w_13193_29093.n497 w_13193_29093.n496 585
R2375 w_13193_29093.n1582 w_13193_29093.n497 585
R2376 w_13193_29093.n1585 w_13193_29093.n1584 585
R2377 w_13193_29093.n1584 w_13193_29093.n1583 585
R2378 w_13193_29093.n1586 w_13193_29093.n494 585
R2379 w_13193_29093.n494 w_13193_29093.n492 585
R2380 w_13193_29093.n1588 w_13193_29093.n1587 585
R2381 w_13193_29093.n1589 w_13193_29093.n1588 585
R2382 w_13193_29093.n1545 w_13193_29093.n491 585
R2383 w_13193_29093.n1589 w_13193_29093.n491 585
R2384 w_13193_29093.n1548 w_13193_29093.n1547 585
R2385 w_13193_29093.n1547 w_13193_29093.n492 585
R2386 w_13193_29093.n1549 w_13193_29093.n498 585
R2387 w_13193_29093.n1583 w_13193_29093.n498 585
R2388 w_13193_29093.n513 w_13193_29093.n499 585
R2389 w_13193_29093.n1582 w_13193_29093.n499 585
R2390 w_13193_29093.n1557 w_13193_29093.n500 585
R2391 w_13193_29093.n1581 w_13193_29093.n500 585
R2392 w_13193_29093.n1560 w_13193_29093.n1559 585
R2393 w_13193_29093.n1560 w_13193_29093.n10 585
R2394 w_13193_29093.n1562 w_13193_29093.n1561 585
R2395 w_13193_29093.n1561 w_13193_29093.n11 585
R2396 w_13193_29093.n510 w_13193_29093.n506 585
R2397 w_13193_29093.n1574 w_13193_29093.n506 585
R2398 w_13193_29093.n1572 w_13193_29093.n1571 585
R2399 w_13193_29093.n1573 w_13193_29093.n1572 585
R2400 w_13193_29093.n508 w_13193_29093.n450 585
R2401 w_13193_29093.n450 w_13193_29093.n449 585
R2402 w_13193_29093.n1747 w_13193_29093.n1746 585
R2403 w_13193_29093.n1748 w_13193_29093.n1747 585
R2404 w_13193_29093.n1744 w_13193_29093.n451 585
R2405 w_13193_29093.n451 w_13193_29093.n12 585
R2406 w_13193_29093.n1052 w_13193_29093.n493 585
R2407 w_13193_29093.n1050 w_13193_29093.n1049 585
R2408 w_13193_29093.n1057 w_13193_29093.n1047 585
R2409 w_13193_29093.n1058 w_13193_29093.n1045 585
R2410 w_13193_29093.n1059 w_13193_29093.n1044 585
R2411 w_13193_29093.n1042 w_13193_29093.n1039 585
R2412 w_13193_29093.n1064 w_13193_29093.n1038 585
R2413 w_13193_29093.n1065 w_13193_29093.n1036 585
R2414 w_13193_29093.n1066 w_13193_29093.n1035 585
R2415 w_13193_29093.n1033 w_13193_29093.n1029 585
R2416 w_13193_29093.n1032 w_13193_29093.n1028 585
R2417 w_13193_29093.n1073 w_13193_29093.n1027 585
R2418 w_13193_29093.n490 w_13193_29093.n383 585
R2419 w_13193_29093.n1521 w_13193_29093.n1520 585
R2420 w_13193_29093.n1527 w_13193_29093.n1518 585
R2421 w_13193_29093.n1528 w_13193_29093.n1516 585
R2422 w_13193_29093.n1529 w_13193_29093.n1515 585
R2423 w_13193_29093.n1513 w_13193_29093.n1510 585
R2424 w_13193_29093.n1534 w_13193_29093.n1509 585
R2425 w_13193_29093.n1535 w_13193_29093.n1507 585
R2426 w_13193_29093.n1536 w_13193_29093.n1506 585
R2427 w_13193_29093.n1504 w_13193_29093.n1500 585
R2428 w_13193_29093.n1503 w_13193_29093.n586 585
R2429 w_13193_29093.n1543 w_13193_29093.n585 585
R2430 w_13193_29093.n584 w_13193_29093.n583 585
R2431 w_13193_29093.n584 w_13193_29093.n16 585
R2432 w_13193_29093.n1053 w_13193_29093.n1052 585
R2433 w_13193_29093.n1055 w_13193_29093.n1050 585
R2434 w_13193_29093.n1057 w_13193_29093.n1056 585
R2435 w_13193_29093.n1058 w_13193_29093.n1041 585
R2436 w_13193_29093.n1060 w_13193_29093.n1059 585
R2437 w_13193_29093.n1062 w_13193_29093.n1039 585
R2438 w_13193_29093.n1064 w_13193_29093.n1063 585
R2439 w_13193_29093.n1065 w_13193_29093.n1030 585
R2440 w_13193_29093.n1067 w_13193_29093.n1066 585
R2441 w_13193_29093.n1069 w_13193_29093.n1029 585
R2442 w_13193_29093.n1070 w_13193_29093.n1028 585
R2443 w_13193_29093.n1073 w_13193_29093.n1072 585
R2444 w_13193_29093.n1523 w_13193_29093.n383 585
R2445 w_13193_29093.n1525 w_13193_29093.n1521 585
R2446 w_13193_29093.n1527 w_13193_29093.n1526 585
R2447 w_13193_29093.n1528 w_13193_29093.n1512 585
R2448 w_13193_29093.n1530 w_13193_29093.n1529 585
R2449 w_13193_29093.n1532 w_13193_29093.n1510 585
R2450 w_13193_29093.n1534 w_13193_29093.n1533 585
R2451 w_13193_29093.n1535 w_13193_29093.n1501 585
R2452 w_13193_29093.n1537 w_13193_29093.n1536 585
R2453 w_13193_29093.n1539 w_13193_29093.n1500 585
R2454 w_13193_29093.n1540 w_13193_29093.n586 585
R2455 w_13193_29093.n1543 w_13193_29093.n1542 585
R2456 w_13193_29093.n1499 w_13193_29093.n583 585
R2457 w_13193_29093.n1499 w_13193_29093.n14 585
R2458 w_13193_29093.n1213 w_13193_29093.n622 585
R2459 w_13193_29093.n1122 w_13193_29093.n624 585
R2460 w_13193_29093.n1127 w_13193_29093.n1123 585
R2461 w_13193_29093.n1128 w_13193_29093.n1119 585
R2462 w_13193_29093.n1129 w_13193_29093.n1118 585
R2463 w_13193_29093.n1116 w_13193_29093.n1113 585
R2464 w_13193_29093.n1134 w_13193_29093.n1112 585
R2465 w_13193_29093.n1135 w_13193_29093.n1110 585
R2466 w_13193_29093.n1136 w_13193_29093.n1109 585
R2467 w_13193_29093.n1107 w_13193_29093.n1104 585
R2468 w_13193_29093.n1141 w_13193_29093.n1103 585
R2469 w_13193_29093.n1142 w_13193_29093.n1101 585
R2470 w_13193_29093.n1213 w_13193_29093.n1212 585
R2471 w_13193_29093.n1125 w_13193_29093.n624 585
R2472 w_13193_29093.n1127 w_13193_29093.n1126 585
R2473 w_13193_29093.n1128 w_13193_29093.n1115 585
R2474 w_13193_29093.n1130 w_13193_29093.n1129 585
R2475 w_13193_29093.n1132 w_13193_29093.n1113 585
R2476 w_13193_29093.n1134 w_13193_29093.n1133 585
R2477 w_13193_29093.n1135 w_13193_29093.n1106 585
R2478 w_13193_29093.n1137 w_13193_29093.n1136 585
R2479 w_13193_29093.n1139 w_13193_29093.n1104 585
R2480 w_13193_29093.n1141 w_13193_29093.n1140 585
R2481 w_13193_29093.n1142 w_13193_29093.n739 585
R2482 w_13193_29093.n1782 w_13193_29093.n1781 585
R2483 w_13193_29093.n1784 w_13193_29093.n420 585
R2484 w_13193_29093.n1786 w_13193_29093.n1785 585
R2485 w_13193_29093.n1787 w_13193_29093.n419 585
R2486 w_13193_29093.n1789 w_13193_29093.n1788 585
R2487 w_13193_29093.n1791 w_13193_29093.n417 585
R2488 w_13193_29093.n1793 w_13193_29093.n1792 585
R2489 w_13193_29093.n1794 w_13193_29093.n416 585
R2490 w_13193_29093.n1796 w_13193_29093.n1795 585
R2491 w_13193_29093.n1798 w_13193_29093.n415 585
R2492 w_13193_29093.n1799 w_13193_29093.n414 585
R2493 w_13193_29093.n1802 w_13193_29093.n1801 585
R2494 w_13193_29093.n2181 w_13193_29093.n2180 585
R2495 w_13193_29093.n2179 w_13193_29093.n2178 585
R2496 w_13193_29093.n2177 w_13193_29093.n277 585
R2497 w_13193_29093.n2175 w_13193_29093.n2174 585
R2498 w_13193_29093.n2173 w_13193_29093.n278 585
R2499 w_13193_29093.n2172 w_13193_29093.n2171 585
R2500 w_13193_29093.n2169 w_13193_29093.n279 585
R2501 w_13193_29093.n2167 w_13193_29093.n2166 585
R2502 w_13193_29093.n2165 w_13193_29093.n280 585
R2503 w_13193_29093.n2164 w_13193_29093.n2163 585
R2504 w_13193_29093.n2161 w_13193_29093.n281 585
R2505 w_13193_29093.n2159 w_13193_29093.n2158 585
R2506 w_13193_29093.n1752 w_13193_29093.n1751 585
R2507 w_13193_29093.n1754 w_13193_29093.n1753 585
R2508 w_13193_29093.n1756 w_13193_29093.n1755 585
R2509 w_13193_29093.n1758 w_13193_29093.n1757 585
R2510 w_13193_29093.n1760 w_13193_29093.n1759 585
R2511 w_13193_29093.n1762 w_13193_29093.n1761 585
R2512 w_13193_29093.n1764 w_13193_29093.n1763 585
R2513 w_13193_29093.n1766 w_13193_29093.n1765 585
R2514 w_13193_29093.n1768 w_13193_29093.n1767 585
R2515 w_13193_29093.n1770 w_13193_29093.n1769 585
R2516 w_13193_29093.n1772 w_13193_29093.n1771 585
R2517 w_13193_29093.n1776 w_13193_29093.n1775 585
R2518 w_13193_29093.n1721 w_13193_29093.n431 585
R2519 w_13193_29093.n1776 w_13193_29093.n431 585
R2520 w_13193_29093.n1723 w_13193_29093.n1722 585
R2521 w_13193_29093.n1725 w_13193_29093.n1724 585
R2522 w_13193_29093.n1727 w_13193_29093.n1726 585
R2523 w_13193_29093.n1729 w_13193_29093.n1728 585
R2524 w_13193_29093.n1731 w_13193_29093.n1730 585
R2525 w_13193_29093.n1733 w_13193_29093.n1732 585
R2526 w_13193_29093.n1735 w_13193_29093.n1734 585
R2527 w_13193_29093.n1737 w_13193_29093.n1736 585
R2528 w_13193_29093.n1739 w_13193_29093.n1738 585
R2529 w_13193_29093.n1741 w_13193_29093.n1740 585
R2530 w_13193_29093.n1743 w_13193_29093.n454 585
R2531 w_13193_29093.n1743 w_13193_29093.n1742 585
R2532 w_13193_29093.n1780 w_13193_29093.n422 585
R2533 w_13193_29093.n1779 w_13193_29093.n1778 585
R2534 w_13193_29093.n424 w_13193_29093.n423 585
R2535 w_13193_29093.n1697 w_13193_29093.n1696 585
R2536 w_13193_29093.n1699 w_13193_29093.n1698 585
R2537 w_13193_29093.n1701 w_13193_29093.n1700 585
R2538 w_13193_29093.n1703 w_13193_29093.n1702 585
R2539 w_13193_29093.n1705 w_13193_29093.n1704 585
R2540 w_13193_29093.n1707 w_13193_29093.n1706 585
R2541 w_13193_29093.n1709 w_13193_29093.n1708 585
R2542 w_13193_29093.n1711 w_13193_29093.n1710 585
R2543 w_13193_29093.n255 w_13193_29093.n242 585
R2544 w_13193_29093.n254 w_13193_29093.n253 585
R2545 w_13193_29093.n254 w_13193_29093.t219 585
R2546 w_13193_29093.n249 w_13193_29093.n244 585
R2547 w_13193_29093.n1082 w_13193_29093.n780 585
R2548 w_13193_29093.n1078 w_13193_29093.n779 585
R2549 w_13193_29093.n1079 w_13193_29093.n1078 585
R2550 w_13193_29093.n1026 w_13193_29093.n901 585
R2551 w_13193_29093.n1026 w_13193_29093.n1025 585
R2552 w_13193_29093.n902 w_13193_29093.n900 585
R2553 w_13193_29093.n1024 w_13193_29093.n902 585
R2554 w_13193_29093.n1022 w_13193_29093.n1021 585
R2555 w_13193_29093.n1023 w_13193_29093.n1022 585
R2556 w_13193_29093.n905 w_13193_29093.n903 585
R2557 w_13193_29093.n987 w_13193_29093.n903 585
R2558 w_13193_29093.n996 w_13193_29093.n995 585
R2559 w_13193_29093.n997 w_13193_29093.n996 585
R2560 w_13193_29093.n992 w_13193_29093.n985 585
R2561 w_13193_29093.n998 w_13193_29093.n985 585
R2562 w_13193_29093.n1000 w_13193_29093.n986 585
R2563 w_13193_29093.n1000 w_13193_29093.n999 585
R2564 w_13193_29093.n1002 w_13193_29093.n1001 585
R2565 w_13193_29093.n1001 w_13193_29093.n29 585
R2566 w_13193_29093.n983 w_13193_29093.n982 585
R2567 w_13193_29093.n982 w_13193_29093.n981 585
R2568 w_13193_29093.n1009 w_13193_29093.n1008 585
R2569 w_13193_29093.n1010 w_13193_29093.n1009 585
R2570 w_13193_29093.n980 w_13193_29093.n926 585
R2571 w_13193_29093.n1011 w_13193_29093.n980 585
R2572 w_13193_29093.n1014 w_13193_29093.n1013 585
R2573 w_13193_29093.n1013 w_13193_29093.n1012 585
R2574 w_13193_29093.n445 w_13193_29093.n444 585
R2575 w_13193_29093.n444 w_13193_29093.n28 585
R2576 w_13193_29093.n1094 w_13193_29093.n746 585
R2577 w_13193_29093.n1096 w_13193_29093.n1095 585
R2578 w_13193_29093.n1097 w_13193_29093.n1096 585
R2579 w_13193_29093.n767 w_13193_29093.n766 585
R2580 w_13193_29093.n764 w_13193_29093.n756 585
R2581 w_13193_29093.n756 w_13193_29093.t21 585
R2582 w_13193_29093.n759 w_13193_29093.n757 585
R2583 w_13193_29093.n1144 w_13193_29093.n740 585
R2584 w_13193_29093.n740 w_13193_29093.n24 585
R2585 w_13193_29093.n1100 w_13193_29093.n1099 585
R2586 w_13193_29093.n1099 w_13193_29093.n1098 585
R2587 w_13193_29093.n813 w_13193_29093.n743 585
R2588 w_13193_29093.n744 w_13193_29093.n743 585
R2589 w_13193_29093.n873 w_13193_29093.n872 585
R2590 w_13193_29093.n874 w_13193_29093.n873 585
R2591 w_13193_29093.n868 w_13193_29093.n812 585
R2592 w_13193_29093.n875 w_13193_29093.n812 585
R2593 w_13193_29093.n878 w_13193_29093.n877 585
R2594 w_13193_29093.n877 w_13193_29093.n876 585
R2595 w_13193_29093.n810 w_13193_29093.n809 585
R2596 w_13193_29093.n809 w_13193_29093.n13 585
R2597 w_13193_29093.n885 w_13193_29093.n884 585
R2598 w_13193_29093.n886 w_13193_29093.n885 585
R2599 w_13193_29093.n807 w_13193_29093.n805 585
R2600 w_13193_29093.n887 w_13193_29093.n807 585
R2601 w_13193_29093.n891 w_13193_29093.n890 585
R2602 w_13193_29093.n890 w_13193_29093.n889 585
R2603 w_13193_29093.n808 w_13193_29093.n785 585
R2604 w_13193_29093.n888 w_13193_29093.n808 585
R2605 w_13193_29093.n898 w_13193_29093.n782 585
R2606 w_13193_29093.n782 w_13193_29093.n781 585
R2607 w_13193_29093.n1076 w_13193_29093.n1075 585
R2608 w_13193_29093.n1077 w_13193_29093.n1076 585
R2609 w_13193_29093.n901 w_13193_29093.n783 585
R2610 w_13193_29093.n783 w_13193_29093.n15 585
R2611 w_13193_29093.n1164 w_13193_29093.n1163 585
R2612 w_13193_29093.n1163 w_13193_29093.n20 585
R2613 w_13193_29093.n1162 w_13193_29093.n634 585
R2614 w_13193_29093.n1162 w_13193_29093.n1161 585
R2615 w_13193_29093.n660 w_13193_29093.n633 585
R2616 w_13193_29093.n1160 w_13193_29093.n633 585
R2617 w_13193_29093.n1158 w_13193_29093.n1157 585
R2618 w_13193_29093.n1159 w_13193_29093.n1158 585
R2619 w_13193_29093.n638 w_13193_29093.n636 585
R2620 w_13193_29093.n636 w_13193_29093.n635 585
R2621 w_13193_29093.n722 w_13193_29093.n721 585
R2622 w_13193_29093.n721 w_13193_29093.n21 585
R2623 w_13193_29093.n725 w_13193_29093.n719 585
R2624 w_13193_29093.n719 w_13193_29093.n718 585
R2625 w_13193_29093.n733 w_13193_29093.n732 585
R2626 w_13193_29093.n734 w_13193_29093.n733 585
R2627 w_13193_29093.n728 w_13193_29093.n717 585
R2628 w_13193_29093.n735 w_13193_29093.n717 585
R2629 w_13193_29093.n737 w_13193_29093.n659 585
R2630 w_13193_29093.n737 w_13193_29093.n736 585
R2631 w_13193_29093.n1150 w_13193_29093.n1149 585
R2632 w_13193_29093.n1149 w_13193_29093.n1148 585
R2633 w_13193_29093.n741 w_13193_29093.n738 585
R2634 w_13193_29093.n1147 w_13193_29093.n738 585
R2635 w_13193_29093.n1145 w_13193_29093.n1144 585
R2636 w_13193_29093.n1146 w_13193_29093.n1145 585
R2637 w_13193_29093.n1211 w_13193_29093.n623 585
R2638 w_13193_29093.n1209 w_13193_29093.n1208 585
R2639 w_13193_29093.n1207 w_13193_29093.n626 585
R2640 w_13193_29093.n1206 w_13193_29093.n1205 585
R2641 w_13193_29093.n1203 w_13193_29093.n627 585
R2642 w_13193_29093.n1201 w_13193_29093.n1200 585
R2643 w_13193_29093.n1199 w_13193_29093.n628 585
R2644 w_13193_29093.n1198 w_13193_29093.n1197 585
R2645 w_13193_29093.n1195 w_13193_29093.n629 585
R2646 w_13193_29093.n1193 w_13193_29093.n1192 585
R2647 w_13193_29093.n1191 w_13193_29093.n630 585
R2648 w_13193_29093.n1190 w_13193_29093.n1189 585
R2649 w_13193_29093.n1961 w_13193_29093.n1960 585
R2650 w_13193_29093.n1939 w_13193_29093.n1938 585
R2651 w_13193_29093.n2030 w_13193_29093.n2029 585
R2652 w_13193_29093.n2032 w_13193_29093.n1937 585
R2653 w_13193_29093.n2035 w_13193_29093.n2034 585
R2654 w_13193_29093.n1934 w_13193_29093.n1933 585
R2655 w_13193_29093.n2045 w_13193_29093.n2044 585
R2656 w_13193_29093.n2047 w_13193_29093.n1932 585
R2657 w_13193_29093.n2050 w_13193_29093.n2049 585
R2658 w_13193_29093.n1929 w_13193_29093.n1925 585
R2659 w_13193_29093.n2061 w_13193_29093.n2060 585
R2660 w_13193_29093.n2063 w_13193_29093.n1924 585
R2661 w_13193_29093.n1187 w_13193_29093.n1186 585
R2662 w_13193_29093.n1185 w_13193_29093.n1184 585
R2663 w_13193_29093.n1183 w_13193_29093.n1182 585
R2664 w_13193_29093.n1181 w_13193_29093.n1180 585
R2665 w_13193_29093.n1179 w_13193_29093.n1178 585
R2666 w_13193_29093.n1177 w_13193_29093.n1176 585
R2667 w_13193_29093.n1175 w_13193_29093.n1174 585
R2668 w_13193_29093.n1173 w_13193_29093.n1172 585
R2669 w_13193_29093.n1171 w_13193_29093.n1170 585
R2670 w_13193_29093.n1169 w_13193_29093.n1168 585
R2671 w_13193_29093.n1167 w_13193_29093.n1166 585
R2672 w_13193_29093.n2153 w_13193_29093.n285 585
R2673 w_13193_29093.n2157 w_13193_29093.n282 585
R2674 w_13193_29093.n2156 w_13193_29093.n2155 585
R2675 w_13193_29093.n284 w_13193_29093.n283 585
R2676 w_13193_29093.n1943 w_13193_29093.n1942 585
R2677 w_13193_29093.n1945 w_13193_29093.n1944 585
R2678 w_13193_29093.n1947 w_13193_29093.n1946 585
R2679 w_13193_29093.n1949 w_13193_29093.n1948 585
R2680 w_13193_29093.n1951 w_13193_29093.n1950 585
R2681 w_13193_29093.n1953 w_13193_29093.n1952 585
R2682 w_13193_29093.n1955 w_13193_29093.n1954 585
R2683 w_13193_29093.n1957 w_13193_29093.n1956 585
R2684 w_13193_29093.n2153 w_13193_29093.n304 585
R2685 w_13193_29093.n2153 w_13193_29093.n2152 585
R2686 w_13193_29093.n2153 w_13193_29093.n292 585
R2687 w_13193_29093.n1233 w_13193_29093.n1232 585
R2688 w_13193_29093.n1229 w_13193_29093.n1228 585
R2689 w_13193_29093.n1302 w_13193_29093.n1301 585
R2690 w_13193_29093.n1304 w_13193_29093.n1227 585
R2691 w_13193_29093.n1307 w_13193_29093.n1306 585
R2692 w_13193_29093.n1224 w_13193_29093.n1223 585
R2693 w_13193_29093.n1317 w_13193_29093.n1316 585
R2694 w_13193_29093.n1319 w_13193_29093.n1222 585
R2695 w_13193_29093.n1322 w_13193_29093.n1321 585
R2696 w_13193_29093.n1219 w_13193_29093.n1215 585
R2697 w_13193_29093.n1333 w_13193_29093.n1332 585
R2698 w_13193_29093.n1335 w_13193_29093.n1214 585
R2699 w_13193_29093.n2131 w_13193_29093.n298 585
R2700 w_13193_29093.n2153 w_13193_29093.n298 585
R2701 w_13193_29093.n2133 w_13193_29093.n2132 585
R2702 w_13193_29093.n2135 w_13193_29093.n2134 585
R2703 w_13193_29093.n2137 w_13193_29093.n2136 585
R2704 w_13193_29093.n2139 w_13193_29093.n2138 585
R2705 w_13193_29093.n2141 w_13193_29093.n2140 585
R2706 w_13193_29093.n2143 w_13193_29093.n2142 585
R2707 w_13193_29093.n2145 w_13193_29093.n2144 585
R2708 w_13193_29093.n2147 w_13193_29093.n2146 585
R2709 w_13193_29093.n2149 w_13193_29093.n2148 585
R2710 w_13193_29093.n2151 w_13193_29093.n2150 585
R2711 w_13193_29093.n2110 w_13193_29093.n2109 585
R2712 w_13193_29093.n2112 w_13193_29093.n313 585
R2713 w_13193_29093.n2114 w_13193_29093.n2113 585
R2714 w_13193_29093.n2115 w_13193_29093.n312 585
R2715 w_13193_29093.n2117 w_13193_29093.n2116 585
R2716 w_13193_29093.n2119 w_13193_29093.n310 585
R2717 w_13193_29093.n2121 w_13193_29093.n2120 585
R2718 w_13193_29093.n2122 w_13193_29093.n309 585
R2719 w_13193_29093.n2124 w_13193_29093.n2123 585
R2720 w_13193_29093.n2126 w_13193_29093.n308 585
R2721 w_13193_29093.n2127 w_13193_29093.n307 585
R2722 w_13193_29093.n2130 w_13193_29093.n2129 585
R2723 w_13193_29093.n1839 w_13193_29093.n357 585
R2724 w_13193_29093.n357 w_13193_29093.n3 585
R2725 w_13193_29093.n1841 w_13193_29093.n1840 585
R2726 w_13193_29093.n1842 w_13193_29093.n1841 585
R2727 w_13193_29093.n382 w_13193_29093.n356 585
R2728 w_13193_29093.n356 w_13193_29093.n355 585
R2729 w_13193_29093.n381 w_13193_29093.n380 585
R2730 w_13193_29093.n380 w_13193_29093.n379 585
R2731 w_13193_29093.n363 w_13193_29093.n358 585
R2732 w_13193_29093.n364 w_13193_29093.n363 585
R2733 w_13193_29093.n362 w_13193_29093.n361 585
R2734 w_13193_29093.n362 w_13193_29093.n2 585
R2735 w_13193_29093.n360 w_13193_29093.n359 585
R2736 w_13193_29093.n359 w_13193_29093.n1 585
R2737 w_13193_29093.n325 w_13193_29093.n324 585
R2738 w_13193_29093.n1912 w_13193_29093.n325 585
R2739 w_13193_29093.n1915 w_13193_29093.n1914 585
R2740 w_13193_29093.n1914 w_13193_29093.n1913 585
R2741 w_13193_29093.n1916 w_13193_29093.n323 585
R2742 w_13193_29093.n326 w_13193_29093.n323 585
R2743 w_13193_29093.n1918 w_13193_29093.n1917 585
R2744 w_13193_29093.n1918 w_13193_29093.n321 585
R2745 w_13193_29093.n1919 w_13193_29093.n316 585
R2746 w_13193_29093.n1920 w_13193_29093.n1919 585
R2747 w_13193_29093.n322 w_13193_29093.n317 585
R2748 w_13193_29093.n1362 w_13193_29093.n1361 585
R2749 w_13193_29093.n1363 w_13193_29093.n1359 585
R2750 w_13193_29093.n1357 w_13193_29093.n1353 585
R2751 w_13193_29093.n1368 w_13193_29093.n1352 585
R2752 w_13193_29093.n1369 w_13193_29093.n1350 585
R2753 w_13193_29093.n1370 w_13193_29093.n1349 585
R2754 w_13193_29093.n1347 w_13193_29093.n1344 585
R2755 w_13193_29093.n1375 w_13193_29093.n1343 585
R2756 w_13193_29093.n1376 w_13193_29093.n1341 585
R2757 w_13193_29093.n1377 w_13193_29093.n1340 585
R2758 w_13193_29093.n1338 w_13193_29093.n1336 585
R2759 w_13193_29093.n1382 w_13193_29093.n621 585
R2760 w_13193_29093.n621 w_13193_29093.n25 585
R2761 w_13193_29093.n317 w_13193_29093.n315 585
R2762 w_13193_29093.n1362 w_13193_29093.n1356 585
R2763 w_13193_29093.n1364 w_13193_29093.n1363 585
R2764 w_13193_29093.n1366 w_13193_29093.n1353 585
R2765 w_13193_29093.n1368 w_13193_29093.n1367 585
R2766 w_13193_29093.n1369 w_13193_29093.n1346 585
R2767 w_13193_29093.n1371 w_13193_29093.n1370 585
R2768 w_13193_29093.n1373 w_13193_29093.n1344 585
R2769 w_13193_29093.n1375 w_13193_29093.n1374 585
R2770 w_13193_29093.n1376 w_13193_29093.n1337 585
R2771 w_13193_29093.n1378 w_13193_29093.n1377 585
R2772 w_13193_29093.n1380 w_13193_29093.n1336 585
R2773 w_13193_29093.n1382 w_13193_29093.n1381 585
R2774 w_13193_29093.n1381 w_13193_29093.n23 585
R2775 w_13193_29093.n2184 w_13193_29093.n2183 585
R2776 w_13193_29093.n2086 w_13193_29093.n273 585
R2777 w_13193_29093.n2088 w_13193_29093.n2087 585
R2778 w_13193_29093.n2084 w_13193_29093.n2081 585
R2779 w_13193_29093.n2093 w_13193_29093.n2080 585
R2780 w_13193_29093.n2094 w_13193_29093.n2078 585
R2781 w_13193_29093.n2095 w_13193_29093.n2077 585
R2782 w_13193_29093.n2075 w_13193_29093.n2072 585
R2783 w_13193_29093.n2100 w_13193_29093.n2071 585
R2784 w_13193_29093.n2101 w_13193_29093.n2069 585
R2785 w_13193_29093.n2102 w_13193_29093.n2068 585
R2786 w_13193_29093.n2066 w_13193_29093.n2064 585
R2787 w_13193_29093.n2107 w_13193_29093.n318 585
R2788 w_13193_29093.n318 w_13193_29093.n25 585
R2789 w_13193_29093.n2183 w_13193_29093.n2182 585
R2790 w_13193_29093.n2083 w_13193_29093.n273 585
R2791 w_13193_29093.n2089 w_13193_29093.n2088 585
R2792 w_13193_29093.n2091 w_13193_29093.n2081 585
R2793 w_13193_29093.n2093 w_13193_29093.n2092 585
R2794 w_13193_29093.n2094 w_13193_29093.n2074 585
R2795 w_13193_29093.n2096 w_13193_29093.n2095 585
R2796 w_13193_29093.n2098 w_13193_29093.n2072 585
R2797 w_13193_29093.n2100 w_13193_29093.n2099 585
R2798 w_13193_29093.n2101 w_13193_29093.n2065 585
R2799 w_13193_29093.n2103 w_13193_29093.n2102 585
R2800 w_13193_29093.n2105 w_13193_29093.n2064 585
R2801 w_13193_29093.n2107 w_13193_29093.n2106 585
R2802 w_13193_29093.n2106 w_13193_29093.n23 585
R2803 w_13193_29093.n1922 w_13193_29093.n1921 585
R2804 w_13193_29093.n1921 w_13193_29093.n1920 585
R2805 w_13193_29093.n1899 w_13193_29093.n320 585
R2806 w_13193_29093.n321 w_13193_29093.n320 585
R2807 w_13193_29093.n1901 w_13193_29093.n1900 585
R2808 w_13193_29093.n1900 w_13193_29093.n326 585
R2809 w_13193_29093.n332 w_13193_29093.n327 585
R2810 w_13193_29093.n1913 w_13193_29093.n327 585
R2811 w_13193_29093.n1911 w_13193_29093.n1910 585
R2812 w_13193_29093.n1912 w_13193_29093.n1911 585
R2813 w_13193_29093.n330 w_13193_29093.n328 585
R2814 w_13193_29093.n328 w_13193_29093.n1 585
R2815 w_13193_29093.n369 w_13193_29093.n368 585
R2816 w_13193_29093.n368 w_13193_29093.n2 585
R2817 w_13193_29093.n366 w_13193_29093.n365 585
R2818 w_13193_29093.n365 w_13193_29093.n364 585
R2819 w_13193_29093.n378 w_13193_29093.n377 585
R2820 w_13193_29093.n379 w_13193_29093.n378 585
R2821 w_13193_29093.n353 w_13193_29093.n351 585
R2822 w_13193_29093.n355 w_13193_29093.n353 585
R2823 w_13193_29093.n1844 w_13193_29093.n1843 585
R2824 w_13193_29093.n1843 w_13193_29093.n1842 585
R2825 w_13193_29093.n386 w_13193_29093.n354 585
R2826 w_13193_29093.n354 w_13193_29093.n3 585
R2827 w_13193_29093.n1654 w_13193_29093.n1653 585
R2828 w_13193_29093.n1655 w_13193_29093.n1654 585
R2829 w_13193_29093.n488 w_13193_29093.n487 585
R2830 w_13193_29093.n489 w_13193_29093.n488 585
R2831 w_13193_29093.n1664 w_13193_29093.n1663 585
R2832 w_13193_29093.n1663 w_13193_29093.n1662 585
R2833 w_13193_29093.n484 w_13193_29093.n474 585
R2834 w_13193_29093.n474 w_13193_29093.n473 585
R2835 w_13193_29093.n1674 w_13193_29093.n1673 585
R2836 w_13193_29093.n1675 w_13193_29093.n1674 585
R2837 w_13193_29093.n477 w_13193_29093.n475 585
R2838 w_13193_29093.n475 w_13193_29093.n7 585
R2839 w_13193_29093.n481 w_13193_29093.n480 585
R2840 w_13193_29093.n480 w_13193_29093.n8 585
R2841 w_13193_29093.n467 w_13193_29093.n466 585
R2842 w_13193_29093.n468 w_13193_29093.n467 585
R2843 w_13193_29093.n1686 w_13193_29093.n1685 585
R2844 w_13193_29093.n1685 w_13193_29093.n1684 585
R2845 w_13193_29093.n463 w_13193_29093.n458 585
R2846 w_13193_29093.n458 w_13193_29093.n457 585
R2847 w_13193_29093.n1716 w_13193_29093.n1715 585
R2848 w_13193_29093.n1717 w_13193_29093.n1716 585
R2849 w_13193_29093.n1713 w_13193_29093.n459 585
R2850 w_13193_29093.n459 w_13193_29093.n9 585
R2851 w_13193_29093.n1776 w_13193_29093.n437 585
R2852 w_13193_29093.n1816 w_13193_29093.n413 585
R2853 w_13193_29093.n1817 w_13193_29093.n411 585
R2854 w_13193_29093.n1818 w_13193_29093.n410 585
R2855 w_13193_29093.n408 w_13193_29093.n405 585
R2856 w_13193_29093.n1823 w_13193_29093.n404 585
R2857 w_13193_29093.n1824 w_13193_29093.n402 585
R2858 w_13193_29093.n1825 w_13193_29093.n401 585
R2859 w_13193_29093.n399 w_13193_29093.n396 585
R2860 w_13193_29093.n1830 w_13193_29093.n395 585
R2861 w_13193_29093.n1831 w_13193_29093.n393 585
R2862 w_13193_29093.n1832 w_13193_29093.n392 585
R2863 w_13193_29093.n390 w_13193_29093.n388 585
R2864 w_13193_29093.n1837 w_13193_29093.n385 585
R2865 w_13193_29093.n385 w_13193_29093.n16 585
R2866 w_13193_29093.n1816 w_13193_29093.n1815 585
R2867 w_13193_29093.n1817 w_13193_29093.n407 585
R2868 w_13193_29093.n1819 w_13193_29093.n1818 585
R2869 w_13193_29093.n1821 w_13193_29093.n405 585
R2870 w_13193_29093.n1823 w_13193_29093.n1822 585
R2871 w_13193_29093.n1824 w_13193_29093.n398 585
R2872 w_13193_29093.n1826 w_13193_29093.n1825 585
R2873 w_13193_29093.n1828 w_13193_29093.n396 585
R2874 w_13193_29093.n1830 w_13193_29093.n1829 585
R2875 w_13193_29093.n1831 w_13193_29093.n389 585
R2876 w_13193_29093.n1833 w_13193_29093.n1832 585
R2877 w_13193_29093.n1835 w_13193_29093.n388 585
R2878 w_13193_29093.n1837 w_13193_29093.n1836 585
R2879 w_13193_29093.n1836 w_13193_29093.n14 585
R2880 w_13193_29093.n1814 w_13193_29093.n1813 585
R2881 w_13193_29093.n1812 w_13193_29093.n1811 585
R2882 w_13193_29093.n1810 w_13193_29093.n1806 585
R2883 w_13193_29093.n1810 w_13193_29093.n31 585
R2884 w_13193_29093.n1809 w_13193_29093.n1807 585
R2885 w_13193_29093.n268 w_13193_29093.n267 585
R2886 w_13193_29093.n2197 w_13193_29093.n2196 585
R2887 w_13193_29093.n2194 w_13193_29093.n266 585
R2888 w_13193_29093.n2193 w_13193_29093.n269 585
R2889 w_13193_29093.n2191 w_13193_29093.n2190 585
R2890 w_13193_29093.n2189 w_13193_29093.n270 585
R2891 w_13193_29093.n2188 w_13193_29093.n2187 585
R2892 w_13193_29093.n2185 w_13193_29093.n271 585
R2893 w_13193_29093.n2185 w_13193_29093.n31 585
R2894 w_13193_29093.n2205 w_13193_29093.n2200 585
R2895 w_13193_29093.n2201 w_13193_29093.n2199 585
R2896 w_13193_29093.n2202 w_13193_29093.n2201 585
R2897 w_13193_29093.n209 w_13193_29093.n208 585
R2898 w_13193_29093.n2526 w_13193_29093.n2525 585
R2899 w_13193_29093.n2503 w_13193_29093.n2502 585
R2900 w_13193_29093.n2501 w_13193_29093.n2497 585
R2901 w_13193_29093.n229 w_13193_29093.n223 585
R2902 w_13193_29093.n231 w_13193_29093.n230 585
R2903 w_13193_29093.n2379 w_13193_29093.n2378 585
R2904 w_13193_29093.n2383 w_13193_29093.n2382 585
R2905 w_13193_29093.n2763 w_13193_29093.n32 585
R2906 w_13193_29093.n2711 w_13193_29093.n2710 585
R2907 w_13193_29093.n2712 w_13193_29093.n2711 585
R2908 w_13193_29093.n2763 w_13193_29093.n2762 585
R2909 w_13193_29093.n2760 w_13193_29093.n33 585
R2910 w_13193_29093.n2712 w_13193_29093.n33 585
R2911 w_13193_29093.t53 w_13193_29093.n1 580.369
R2912 w_13193_29093.t53 w_13193_29093.n4 580.369
R2913 w_13193_29093.t53 w_13193_29093.n7 580.369
R2914 w_13193_29093.t53 w_13193_29093.n10 580.369
R2915 w_13193_29093.t162 w_13193_29093.n2222 576.699
R2916 w_13193_29093.n2259 w_13193_29093.t200 576.699
R2917 w_13193_29093.n2259 w_13193_29093.t206 576.699
R2918 w_13193_29093.n2276 w_13193_29093.t143 576.699
R2919 w_13193_29093.t174 w_13193_29093.n2277 576.699
R2920 w_13193_29093.t50 w_13193_29093.n2278 576.699
R2921 w_13193_29093.n2279 w_13193_29093.t154 576.699
R2922 w_13193_29093.n2368 w_13193_29093.t316 566.966
R2923 w_13193_29093.t53 w_13193_29093.t2 541.827
R2924 w_13193_29093.t53 w_13193_29093.t37 541.827
R2925 w_13193_29093.t141 w_13193_29093.n2223 533.981
R2926 w_13193_29093.t4 w_13193_29093.n2712 525.878
R2927 w_13193_29093.t189 w_13193_29093.n2387 524.22
R2928 w_13193_29093.t148 w_13193_29093.t224 523.244
R2929 w_13193_29093.n2446 w_13193_29093.t168 520.611
R2930 w_13193_29093.t146 w_13193_29093.n2460 520.611
R2931 w_13193_29093.n2461 w_13193_29093.t193 520.611
R2932 w_13193_29093.n2375 w_13193_29093.t254 487.568
R2933 w_13193_29093.t208 w_13193_29093.t162 469.904
R2934 w_13193_29093.t200 w_13193_29093.t233 469.904
R2935 w_13193_29093.t206 w_13193_29093.t228 469.904
R2936 w_13193_29093.t143 w_13193_29093.t141 469.904
R2937 w_13193_29093.t128 w_13193_29093.t174 469.904
R2938 w_13193_29093.n2695 w_13193_29093.t231 463.784
R2939 w_13193_29093.t195 w_13193_29093.n2542 459.776
R2940 w_13193_29093.t129 w_13193_29093.n2548 459.776
R2941 w_13193_29093.t140 w_13193_29093.t134 454.832
R2942 w_13193_29093.t213 w_13193_29093.t281 449.502
R2943 w_13193_29093.n2445 w_13193_29093.t154 422.62
R2944 w_13193_29093.t281 w_13193_29093.n30 415.76
R2945 w_13193_29093.t191 w_13193_29093.n68 392.433
R2946 w_13193_29093.t287 w_13193_29093.t138 380.541
R2947 w_13193_29093.t71 w_13193_29093.t35 378.125
R2948 w_13193_29093.t4 w_13193_29093.n2704 352.193
R2949 w_13193_29093.n225 w_13193_29093.t100 336.329
R2950 w_13193_29093.n225 w_13193_29093.t54 336.329
R2951 w_13193_29093.n2498 w_13193_29093.t66 336.329
R2952 w_13193_29093.n2498 w_13193_29093.t70 336.329
R2953 w_13193_29093.t282 w_13193_29093.t11 332.974
R2954 w_13193_29093.n1920 w_13193_29093.t53 323.926
R2955 w_13193_29093.n1386 w_13193_29093.t53 323.926
R2956 w_13193_29093.n1655 w_13193_29093.t53 323.926
R2957 w_13193_29093.t53 w_13193_29093.n1589 323.926
R2958 w_13193_29093.t197 w_13193_29093.n2693 321.082
R2959 w_13193_29093.n2523 w_13193_29093.t78 320.7
R2960 w_13193_29093.n2380 w_13193_29093.t86 320.7
R2961 w_13193_29093.t284 w_13193_29093.t0 317.969
R2962 w_13193_29093.t122 w_13193_29093.t220 317.969
R2963 w_13193_29093.t120 w_13193_29093.t79 317.969
R2964 w_13193_29093.t116 w_13193_29093.n159 309.375
R2965 w_13193_29093.n2533 w_13193_29093.t67 309.375
R2966 w_13193_29093.t224 w_13193_29093.t118 309.19
R2967 w_13193_29093.n233 w_13193_29093.n221 305
R2968 w_13193_29093.n227 w_13193_29093.n224 305
R2969 w_13193_29093.n2506 w_13193_29093.n2496 305
R2970 w_13193_29093.n2500 w_13193_29093.n2499 305
R2971 w_13193_29093.n2707 w_13193_29093.t93 304.634
R2972 w_13193_29093.n2715 w_13193_29093.t63 304.634
R2973 w_13193_29093.n2718 w_13193_29093.t96 304.634
R2974 w_13193_29093.n2723 w_13193_29093.t82 304.634
R2975 w_13193_29093.n97 w_13193_29093.t283 302.334
R2976 w_13193_29093.n2684 w_13193_29093.t177 302.334
R2977 w_13193_29093.n2678 w_13193_29093.t255 302.334
R2978 w_13193_29093.n2535 w_13193_29093.t108 301.574
R2979 w_13193_29093.n2438 w_13193_29093.t306 293.161
R2980 w_13193_29093.n57 w_13193_29093.t90 292.584
R2981 w_13193_29093.n2759 w_13193_29093.t60 292.584
R2982 w_13193_29093.n2531 w_13193_29093.n2530 292.188
R2983 w_13193_29093.t53 w_13193_29093.n0 281.973
R2984 w_13193_29093.n2762 w_13193_29093.n33 275.8
R2985 w_13193_29093.n2711 w_13193_29093.n32 275.8
R2986 w_13193_29093.n2376 w_13193_29093.t199 273.514
R2987 w_13193_29093.t53 w_13193_29093.n3 269.94
R2988 w_13193_29093.t53 w_13193_29093.n6 269.94
R2989 w_13193_29093.t53 w_13193_29093.n9 269.94
R2990 w_13193_29093.t53 w_13193_29093.n12 269.94
R2991 w_13193_29093.n2203 w_13193_29093.n2202 267.704
R2992 w_13193_29093.t138 w_13193_29093.t282 261.623
R2993 w_13193_29093.t11 w_13193_29093.t45 261.623
R2994 w_13193_29093.t15 w_13193_29093.t43 261.623
R2995 w_13193_29093.t216 w_13193_29093.t172 261.623
R2996 w_13193_29093.t41 w_13193_29093.t180 261.623
R2997 w_13193_29093.n2389 w_13193_29093.n2376 261.623
R2998 w_13193_29093.t248 w_13193_29093.t237 261.623
R2999 w_13193_29093.n89 w_13193_29093.n88 260.199
R3000 w_13193_29093.n203 w_13193_29093.t256 260
R3001 w_13193_29093.n2553 w_13193_29093.t256 260
R3002 w_13193_29093.n262 w_13193_29093.t3 260
R3003 w_13193_29093.t3 w_13193_29093.n259 260
R3004 w_13193_29093.n2185 w_13193_29093.n2184 259.416
R3005 w_13193_29093.n2159 w_13193_29093.n282 259.416
R3006 w_13193_29093.n1801 w_13193_29093.n413 259.416
R3007 w_13193_29093.n1189 w_13193_29093.n1187 259.416
R3008 w_13193_29093.n1588 w_13193_29093.n493 259.416
R3009 w_13193_29093.n1656 w_13193_29093.n490 259.416
R3010 w_13193_29093.n1919 w_13193_29093.n322 259.416
R3011 w_13193_29093.n1385 w_13193_29093.n622 259.416
R3012 w_13193_29093.n2129 w_13193_29093.n298 259.416
R3013 w_13193_29093.n1618 w_13193_29093.n1617 258.334
R3014 w_13193_29093.n1865 w_13193_29093.n1864 258.334
R3015 w_13193_29093.n1991 w_13193_29093.n1990 258.334
R3016 w_13193_29093.n548 w_13193_29093.n547 258.334
R3017 w_13193_29093.n962 w_13193_29093.n961 258.334
R3018 w_13193_29093.n1425 w_13193_29093.n1424 258.334
R3019 w_13193_29093.n830 w_13193_29093.n829 258.334
R3020 w_13193_29093.n699 w_13193_29093.n698 258.334
R3021 w_13193_29093.n1263 w_13193_29093.n1262 258.334
R3022 w_13193_29093.n1048 w_13193_29093.n16 254.34
R3023 w_13193_29093.n1046 w_13193_29093.n16 254.34
R3024 w_13193_29093.n1043 w_13193_29093.n16 254.34
R3025 w_13193_29093.n1037 w_13193_29093.n16 254.34
R3026 w_13193_29093.n1034 w_13193_29093.n16 254.34
R3027 w_13193_29093.n1031 w_13193_29093.n16 254.34
R3028 w_13193_29093.n1519 w_13193_29093.n16 254.34
R3029 w_13193_29093.n1517 w_13193_29093.n16 254.34
R3030 w_13193_29093.n1514 w_13193_29093.n16 254.34
R3031 w_13193_29093.n1508 w_13193_29093.n16 254.34
R3032 w_13193_29093.n1505 w_13193_29093.n16 254.34
R3033 w_13193_29093.n1502 w_13193_29093.n16 254.34
R3034 w_13193_29093.n1054 w_13193_29093.n14 254.34
R3035 w_13193_29093.n1051 w_13193_29093.n14 254.34
R3036 w_13193_29093.n1061 w_13193_29093.n14 254.34
R3037 w_13193_29093.n1040 w_13193_29093.n14 254.34
R3038 w_13193_29093.n1068 w_13193_29093.n14 254.34
R3039 w_13193_29093.n1071 w_13193_29093.n14 254.34
R3040 w_13193_29093.n1524 w_13193_29093.n14 254.34
R3041 w_13193_29093.n1522 w_13193_29093.n14 254.34
R3042 w_13193_29093.n1531 w_13193_29093.n14 254.34
R3043 w_13193_29093.n1511 w_13193_29093.n14 254.34
R3044 w_13193_29093.n1538 w_13193_29093.n14 254.34
R3045 w_13193_29093.n1541 w_13193_29093.n14 254.34
R3046 w_13193_29093.n1121 w_13193_29093.n25 254.34
R3047 w_13193_29093.n1120 w_13193_29093.n25 254.34
R3048 w_13193_29093.n1117 w_13193_29093.n25 254.34
R3049 w_13193_29093.n1111 w_13193_29093.n25 254.34
R3050 w_13193_29093.n1108 w_13193_29093.n25 254.34
R3051 w_13193_29093.n1102 w_13193_29093.n25 254.34
R3052 w_13193_29093.n625 w_13193_29093.n23 254.34
R3053 w_13193_29093.n1124 w_13193_29093.n23 254.34
R3054 w_13193_29093.n1131 w_13193_29093.n23 254.34
R3055 w_13193_29093.n1114 w_13193_29093.n23 254.34
R3056 w_13193_29093.n1138 w_13193_29093.n23 254.34
R3057 w_13193_29093.n1105 w_13193_29093.n23 254.34
R3058 w_13193_29093.n1783 w_13193_29093.n31 254.34
R3059 w_13193_29093.n421 w_13193_29093.n31 254.34
R3060 w_13193_29093.n1790 w_13193_29093.n31 254.34
R3061 w_13193_29093.n418 w_13193_29093.n31 254.34
R3062 w_13193_29093.n1797 w_13193_29093.n31 254.34
R3063 w_13193_29093.n1800 w_13193_29093.n31 254.34
R3064 w_13193_29093.n276 w_13193_29093.n31 254.34
R3065 w_13193_29093.n2176 w_13193_29093.n31 254.34
R3066 w_13193_29093.n2170 w_13193_29093.n31 254.34
R3067 w_13193_29093.n2168 w_13193_29093.n31 254.34
R3068 w_13193_29093.n2162 w_13193_29093.n31 254.34
R3069 w_13193_29093.n2160 w_13193_29093.n31 254.34
R3070 w_13193_29093.n1776 w_13193_29093.n438 254.34
R3071 w_13193_29093.n1776 w_13193_29093.n439 254.34
R3072 w_13193_29093.n1776 w_13193_29093.n440 254.34
R3073 w_13193_29093.n1776 w_13193_29093.n441 254.34
R3074 w_13193_29093.n1776 w_13193_29093.n442 254.34
R3075 w_13193_29093.n1776 w_13193_29093.n443 254.34
R3076 w_13193_29093.n1774 w_13193_29093.n1773 254.34
R3077 w_13193_29093.n1776 w_13193_29093.n430 254.34
R3078 w_13193_29093.n1776 w_13193_29093.n429 254.34
R3079 w_13193_29093.n1776 w_13193_29093.n428 254.34
R3080 w_13193_29093.n1776 w_13193_29093.n427 254.34
R3081 w_13193_29093.n1776 w_13193_29093.n426 254.34
R3082 w_13193_29093.n1776 w_13193_29093.n425 254.34
R3083 w_13193_29093.n1777 w_13193_29093.n1776 254.34
R3084 w_13193_29093.n1776 w_13193_29093.n436 254.34
R3085 w_13193_29093.n1776 w_13193_29093.n435 254.34
R3086 w_13193_29093.n1776 w_13193_29093.n434 254.34
R3087 w_13193_29093.n1776 w_13193_29093.n433 254.34
R3088 w_13193_29093.n1210 w_13193_29093.n19 254.34
R3089 w_13193_29093.n1204 w_13193_29093.n19 254.34
R3090 w_13193_29093.n1202 w_13193_29093.n19 254.34
R3091 w_13193_29093.n1196 w_13193_29093.n19 254.34
R3092 w_13193_29093.n1194 w_13193_29093.n19 254.34
R3093 w_13193_29093.n1188 w_13193_29093.n19 254.34
R3094 w_13193_29093.n1959 w_13193_29093.n26 254.34
R3095 w_13193_29093.n2031 w_13193_29093.n26 254.34
R3096 w_13193_29093.n2033 w_13193_29093.n26 254.34
R3097 w_13193_29093.n2046 w_13193_29093.n26 254.34
R3098 w_13193_29093.n2048 w_13193_29093.n26 254.34
R3099 w_13193_29093.n2062 w_13193_29093.n26 254.34
R3100 w_13193_29093.n2153 w_13193_29093.n291 254.34
R3101 w_13193_29093.n2153 w_13193_29093.n290 254.34
R3102 w_13193_29093.n2153 w_13193_29093.n289 254.34
R3103 w_13193_29093.n2153 w_13193_29093.n288 254.34
R3104 w_13193_29093.n2153 w_13193_29093.n287 254.34
R3105 w_13193_29093.n2153 w_13193_29093.n286 254.34
R3106 w_13193_29093.n1165 w_13193_29093.n631 254.34
R3107 w_13193_29093.n2154 w_13193_29093.n2153 254.34
R3108 w_13193_29093.n2153 w_13193_29093.n299 254.34
R3109 w_13193_29093.n2153 w_13193_29093.n300 254.34
R3110 w_13193_29093.n2153 w_13193_29093.n301 254.34
R3111 w_13193_29093.n2153 w_13193_29093.n302 254.34
R3112 w_13193_29093.n2153 w_13193_29093.n303 254.34
R3113 w_13193_29093.n1958 w_13193_29093.n1941 254.34
R3114 w_13193_29093.n306 w_13193_29093.n305 254.34
R3115 w_13193_29093.n1231 w_13193_29093.n22 254.34
R3116 w_13193_29093.n1303 w_13193_29093.n22 254.34
R3117 w_13193_29093.n1305 w_13193_29093.n22 254.34
R3118 w_13193_29093.n1318 w_13193_29093.n22 254.34
R3119 w_13193_29093.n1320 w_13193_29093.n22 254.34
R3120 w_13193_29093.n1334 w_13193_29093.n22 254.34
R3121 w_13193_29093.n2153 w_13193_29093.n297 254.34
R3122 w_13193_29093.n2153 w_13193_29093.n296 254.34
R3123 w_13193_29093.n2153 w_13193_29093.n295 254.34
R3124 w_13193_29093.n2153 w_13193_29093.n294 254.34
R3125 w_13193_29093.n2153 w_13193_29093.n293 254.34
R3126 w_13193_29093.n2111 w_13193_29093.n18 254.34
R3127 w_13193_29093.n314 w_13193_29093.n18 254.34
R3128 w_13193_29093.n2118 w_13193_29093.n18 254.34
R3129 w_13193_29093.n311 w_13193_29093.n18 254.34
R3130 w_13193_29093.n2125 w_13193_29093.n18 254.34
R3131 w_13193_29093.n2128 w_13193_29093.n18 254.34
R3132 w_13193_29093.n1360 w_13193_29093.n25 254.34
R3133 w_13193_29093.n1358 w_13193_29093.n25 254.34
R3134 w_13193_29093.n1351 w_13193_29093.n25 254.34
R3135 w_13193_29093.n1348 w_13193_29093.n25 254.34
R3136 w_13193_29093.n1342 w_13193_29093.n25 254.34
R3137 w_13193_29093.n1339 w_13193_29093.n25 254.34
R3138 w_13193_29093.n1355 w_13193_29093.n23 254.34
R3139 w_13193_29093.n1365 w_13193_29093.n23 254.34
R3140 w_13193_29093.n1354 w_13193_29093.n23 254.34
R3141 w_13193_29093.n1372 w_13193_29093.n23 254.34
R3142 w_13193_29093.n1345 w_13193_29093.n23 254.34
R3143 w_13193_29093.n1379 w_13193_29093.n23 254.34
R3144 w_13193_29093.n272 w_13193_29093.n25 254.34
R3145 w_13193_29093.n2085 w_13193_29093.n25 254.34
R3146 w_13193_29093.n2079 w_13193_29093.n25 254.34
R3147 w_13193_29093.n2076 w_13193_29093.n25 254.34
R3148 w_13193_29093.n2070 w_13193_29093.n25 254.34
R3149 w_13193_29093.n2067 w_13193_29093.n25 254.34
R3150 w_13193_29093.n275 w_13193_29093.n23 254.34
R3151 w_13193_29093.n2090 w_13193_29093.n23 254.34
R3152 w_13193_29093.n2082 w_13193_29093.n23 254.34
R3153 w_13193_29093.n2097 w_13193_29093.n23 254.34
R3154 w_13193_29093.n2073 w_13193_29093.n23 254.34
R3155 w_13193_29093.n2104 w_13193_29093.n23 254.34
R3156 w_13193_29093.n1712 w_13193_29093.n1695 254.34
R3157 w_13193_29093.n1776 w_13193_29093.n432 254.34
R3158 w_13193_29093.n412 w_13193_29093.n16 254.34
R3159 w_13193_29093.n409 w_13193_29093.n16 254.34
R3160 w_13193_29093.n403 w_13193_29093.n16 254.34
R3161 w_13193_29093.n400 w_13193_29093.n16 254.34
R3162 w_13193_29093.n394 w_13193_29093.n16 254.34
R3163 w_13193_29093.n391 w_13193_29093.n16 254.34
R3164 w_13193_29093.n1804 w_13193_29093.n14 254.34
R3165 w_13193_29093.n1820 w_13193_29093.n14 254.34
R3166 w_13193_29093.n406 w_13193_29093.n14 254.34
R3167 w_13193_29093.n1827 w_13193_29093.n14 254.34
R3168 w_13193_29093.n397 w_13193_29093.n14 254.34
R3169 w_13193_29093.n1834 w_13193_29093.n14 254.34
R3170 w_13193_29093.n1805 w_13193_29093.n31 254.34
R3171 w_13193_29093.n1808 w_13193_29093.n31 254.34
R3172 w_13193_29093.n2195 w_13193_29093.n31 254.34
R3173 w_13193_29093.n2192 w_13193_29093.n31 254.34
R3174 w_13193_29093.n2186 w_13193_29093.n31 254.34
R3175 w_13193_29093.n87 w_13193_29093.n86 254.333
R3176 w_13193_29093.n82 w_13193_29093.n81 254.333
R3177 w_13193_29093.n106 w_13193_29093.n105 254.333
R3178 w_13193_29093.n114 w_13193_29093.n113 254.333
R3179 w_13193_29093.n126 w_13193_29093.n125 254.333
R3180 w_13193_29093.n73 w_13193_29093.n72 254.333
R3181 w_13193_29093.n142 w_13193_29093.n141 254.333
R3182 w_13193_29093.n2670 w_13193_29093.n144 254.333
R3183 w_13193_29093.n151 w_13193_29093.n150 254.333
R3184 w_13193_29093.n2650 w_13193_29093.n153 254.333
R3185 w_13193_29093.n157 w_13193_29093.n156 253.114
R3186 w_13193_29093.n1815 w_13193_29093.n1814 251.614
R3187 w_13193_29093.n2182 w_13193_29093.n2181 251.614
R3188 w_13193_29093.n1782 w_13193_29093.n422 251.614
R3189 w_13193_29093.n1212 w_13193_29093.n1211 251.614
R3190 w_13193_29093.n1751 w_13193_29093.n1750 251.614
R3191 w_13193_29093.n1719 w_13193_29093.n431 251.614
R3192 w_13193_29093.n1523 w_13193_29093.n357 251.614
R3193 w_13193_29093.n1053 w_13193_29093.n591 251.614
R3194 w_13193_29093.n2110 w_13193_29093.n315 251.614
R3195 w_13193_29093.n1080 w_13193_29093.n1079 250.349
R3196 w_13193_29093.n1097 w_13193_29093.n745 250.349
R3197 w_13193_29093.n2530 w_13193_29093.n2529 250.349
R3198 w_13193_29093.n2530 w_13193_29093.n207 250.349
R3199 w_13193_29093.n2532 w_13193_29093.n206 250.349
R3200 w_13193_29093.n2532 w_13193_29093.n205 250.349
R3201 w_13193_29093.n226 w_13193_29093.n204 250.349
R3202 w_13193_29093.n232 w_13193_29093.n204 250.349
R3203 w_13193_29093.n2387 w_13193_29093.n2386 250.349
R3204 w_13193_29093.n2387 w_13193_29093.n2377 250.349
R3205 w_13193_29093.n2434 w_13193_29093.t19 249.731
R3206 w_13193_29093.n759 w_13193_29093.n756 246.25
R3207 w_13193_29093.n767 w_13193_29093.n756 246.25
R3208 w_13193_29093.n254 w_13193_29093.n244 246.25
R3209 w_13193_29093.n255 w_13193_29093.n254 246.25
R3210 w_13193_29093.n2708 w_13193_29093.t95 245
R3211 w_13193_29093.n2716 w_13193_29093.t64 245
R3212 w_13193_29093.n2717 w_13193_29093.t97 245
R3213 w_13193_29093.n2722 w_13193_29093.t85 245
R3214 w_13193_29093.n261 w_13193_29093.n260 241.643
R3215 w_13193_29093.n256 w_13193_29093.t219 241.643
R3216 w_13193_29093.n247 w_13193_29093.t219 241.643
R3217 w_13193_29093.n768 w_13193_29093.t21 241.643
R3218 w_13193_29093.n760 w_13193_29093.t21 241.643
R3219 w_13193_29093.n2552 w_13193_29093.n2551 241.643
R3220 w_13193_29093.n2548 w_13193_29093.n2543 241.643
R3221 w_13193_29093.n2542 w_13193_29093.n2536 241.643
R3222 w_13193_29093.n2534 w_13193_29093.n204 240.625
R3223 w_13193_29093.n2693 w_13193_29093.n68 237.839
R3224 w_13193_29093.t180 w_13193_29093.t113 237.839
R3225 w_13193_29093.t296 w_13193_29093.t267 236.281
R3226 w_13193_29093.n2692 w_13193_29093.t198 233
R3227 w_13193_29093.n147 w_13193_29093.t249 233
R3228 w_13193_29093.n2546 w_13193_29093.t260 233
R3229 w_13193_29093.n2549 w_13193_29093.t262 233
R3230 w_13193_29093.n2540 w_13193_29093.t257 233
R3231 w_13193_29093.n2632 w_13193_29093.n162 225.534
R3232 w_13193_29093.n164 w_13193_29093.n163 225.534
R3233 w_13193_29093.n2620 w_13193_29093.n168 225.534
R3234 w_13193_29093.n2613 w_13193_29093.n173 225.534
R3235 w_13193_29093.n177 w_13193_29093.n176 225.534
R3236 w_13193_29093.n2601 w_13193_29093.n180 225.534
R3237 w_13193_29093.n2594 w_13193_29093.n185 225.534
R3238 w_13193_29093.n189 w_13193_29093.n188 225.534
R3239 w_13193_29093.n2582 w_13193_29093.n2581 225.534
R3240 w_13193_29093.t150 w_13193_29093.n61 218.321
R3241 w_13193_29093.n2765 w_13193_29093.n2764 217.106
R3242 w_13193_29093.t7 w_13193_29093.t156 214.054
R3243 w_13193_29093.t136 w_13193_29093.t287 214.054
R3244 w_13193_29093.t45 w_13193_29093.t311 214.054
R3245 w_13193_29093.t19 w_13193_29093.t302 214.054
R3246 w_13193_29093.n41 w_13193_29093.n40 210.601
R3247 w_13193_29093.n2706 w_13193_29093.n2705 210.601
R3248 w_13193_29093.n2714 w_13193_29093.n2713 210.601
R3249 w_13193_29093.n2231 w_13193_29093.t125 204.458
R3250 w_13193_29093.n2350 w_13193_29093.t292 204.458
R3251 w_13193_29093.n2336 w_13193_29093.t12 204.458
R3252 w_13193_29093.n2331 w_13193_29093.t288 204.458
R3253 w_13193_29093.n2323 w_13193_29093.t209 204.458
R3254 w_13193_29093.n2318 w_13193_29093.t234 204.458
R3255 w_13193_29093.n2305 w_13193_29093.t142 204.458
R3256 w_13193_29093.n2310 w_13193_29093.t229 204.458
R3257 w_13193_29093.n2725 w_13193_29093.n58 204.201
R3258 w_13193_29093.n2719 w_13193_29093.n59 204.201
R3259 w_13193_29093.n2724 w_13193_29093.n2720 204.201
R3260 w_13193_29093.t25 w_13193_29093.n2765 203.913
R3261 w_13193_29093.t205 w_13193_29093.n2694 202.162
R3262 w_13193_29093.n2382 w_13193_29093.n2378 197
R3263 w_13193_29093.n231 w_13193_29093.n223 197
R3264 w_13193_29093.n2502 w_13193_29093.n2501 197
R3265 w_13193_29093.n2525 w_13193_29093.n208 197
R3266 w_13193_29093.n1096 w_13193_29093.n746 197
R3267 w_13193_29093.n1078 w_13193_29093.n780 197
R3268 w_13193_29093.t199 w_13193_29093.t41 190.27
R3269 w_13193_29093.t293 w_13193_29093.t230 190.27
R3270 w_13193_29093.t308 w_13193_29093.t222 189.062
R3271 w_13193_29093.t222 w_13193_29093.t203 189.062
R3272 w_13193_29093.t132 w_13193_29093.t298 189.062
R3273 w_13193_29093.t272 w_13193_29093.t105 189.062
R3274 w_13193_29093.t276 w_13193_29093.t274 189.062
R3275 w_13193_29093.t271 w_13193_29093.t164 189.062
R3276 w_13193_29093.t250 w_13193_29093.t304 189.062
R3277 w_13193_29093.t29 w_13193_29093.t235 189.062
R3278 w_13193_29093.t145 w_13193_29093.t160 189.062
R3279 w_13193_29093.n229 w_13193_29093.n224 185
R3280 w_13193_29093.n230 w_13193_29093.n221 185
R3281 w_13193_29093.n2503 w_13193_29093.n2500 185
R3282 w_13193_29093.n2497 w_13193_29093.n2496 185
R3283 w_13193_29093.n1617 w_13193_29093.n1599 185
R3284 w_13193_29093.n1615 w_13193_29093.n1614 185
R3285 w_13193_29093.n1613 w_13193_29093.n1601 185
R3286 w_13193_29093.n1612 w_13193_29093.n1611 185
R3287 w_13193_29093.n1609 w_13193_29093.n1602 185
R3288 w_13193_29093.n1607 w_13193_29093.n1606 185
R3289 w_13193_29093.n1605 w_13193_29093.n1604 185
R3290 w_13193_29093.n462 w_13193_29093.n461 185
R3291 w_13193_29093.n1694 w_13193_29093.n1693 185
R3292 w_13193_29093.n1619 w_13193_29093.n1618 185
R3293 w_13193_29093.n1620 w_13193_29093.n1598 185
R3294 w_13193_29093.n1622 w_13193_29093.n1621 185
R3295 w_13193_29093.n1624 w_13193_29093.n1596 185
R3296 w_13193_29093.n1626 w_13193_29093.n1625 185
R3297 w_13193_29093.n1627 w_13193_29093.n1595 185
R3298 w_13193_29093.n1629 w_13193_29093.n1628 185
R3299 w_13193_29093.n1631 w_13193_29093.n1594 185
R3300 w_13193_29093.n1634 w_13193_29093.n1633 185
R3301 w_13193_29093.n1635 w_13193_29093.n1593 185
R3302 w_13193_29093.n1637 w_13193_29093.n1636 185
R3303 w_13193_29093.n1639 w_13193_29093.n1592 185
R3304 w_13193_29093.n1642 w_13193_29093.n1641 185
R3305 w_13193_29093.n1643 w_13193_29093.n1591 185
R3306 w_13193_29093.n1645 w_13193_29093.n1644 185
R3307 w_13193_29093.n1647 w_13193_29093.n1590 185
R3308 w_13193_29093.n1650 w_13193_29093.n1649 185
R3309 w_13193_29093.n1651 w_13193_29093.n486 185
R3310 w_13193_29093.n1864 w_13193_29093.n344 185
R3311 w_13193_29093.n1862 w_13193_29093.n1861 185
R3312 w_13193_29093.n1860 w_13193_29093.n346 185
R3313 w_13193_29093.n1859 w_13193_29093.n1858 185
R3314 w_13193_29093.n1856 w_13193_29093.n347 185
R3315 w_13193_29093.n1854 w_13193_29093.n1853 185
R3316 w_13193_29093.n1852 w_13193_29093.n348 185
R3317 w_13193_29093.n1851 w_13193_29093.n1850 185
R3318 w_13193_29093.n1848 w_13193_29093.n349 185
R3319 w_13193_29093.n1866 w_13193_29093.n1865 185
R3320 w_13193_29093.n1867 w_13193_29093.n343 185
R3321 w_13193_29093.n1869 w_13193_29093.n1868 185
R3322 w_13193_29093.n1871 w_13193_29093.n341 185
R3323 w_13193_29093.n1873 w_13193_29093.n1872 185
R3324 w_13193_29093.n1874 w_13193_29093.n340 185
R3325 w_13193_29093.n1876 w_13193_29093.n1875 185
R3326 w_13193_29093.n1878 w_13193_29093.n339 185
R3327 w_13193_29093.n1881 w_13193_29093.n1880 185
R3328 w_13193_29093.n1882 w_13193_29093.n338 185
R3329 w_13193_29093.n1884 w_13193_29093.n1883 185
R3330 w_13193_29093.n1886 w_13193_29093.n337 185
R3331 w_13193_29093.n1889 w_13193_29093.n1888 185
R3332 w_13193_29093.n1890 w_13193_29093.n336 185
R3333 w_13193_29093.n1892 w_13193_29093.n1891 185
R3334 w_13193_29093.n1894 w_13193_29093.n335 185
R3335 w_13193_29093.n1896 w_13193_29093.n1895 185
R3336 w_13193_29093.n1898 w_13193_29093.n1897 185
R3337 w_13193_29093.n769 w_13193_29093.n755 185
R3338 w_13193_29093.n762 w_13193_29093.n761 185
R3339 w_13193_29093.n246 w_13193_29093.n242 185
R3340 w_13193_29093.n248 w_13193_29093.n246 185
R3341 w_13193_29093.n1990 w_13193_29093.n1972 185
R3342 w_13193_29093.n1988 w_13193_29093.n1987 185
R3343 w_13193_29093.n1986 w_13193_29093.n1974 185
R3344 w_13193_29093.n1985 w_13193_29093.n1984 185
R3345 w_13193_29093.n1982 w_13193_29093.n1975 185
R3346 w_13193_29093.n1980 w_13193_29093.n1979 185
R3347 w_13193_29093.n1978 w_13193_29093.n1977 185
R3348 w_13193_29093.n1928 w_13193_29093.n1927 185
R3349 w_13193_29093.n2058 w_13193_29093.n2057 185
R3350 w_13193_29093.n1992 w_13193_29093.n1991 185
R3351 w_13193_29093.n1993 w_13193_29093.n1971 185
R3352 w_13193_29093.n1995 w_13193_29093.n1994 185
R3353 w_13193_29093.n1997 w_13193_29093.n1969 185
R3354 w_13193_29093.n1999 w_13193_29093.n1998 185
R3355 w_13193_29093.n2000 w_13193_29093.n1968 185
R3356 w_13193_29093.n2002 w_13193_29093.n2001 185
R3357 w_13193_29093.n2004 w_13193_29093.n1967 185
R3358 w_13193_29093.n2007 w_13193_29093.n2006 185
R3359 w_13193_29093.n2008 w_13193_29093.n1966 185
R3360 w_13193_29093.n2010 w_13193_29093.n2009 185
R3361 w_13193_29093.n2012 w_13193_29093.n1965 185
R3362 w_13193_29093.n2015 w_13193_29093.n2014 185
R3363 w_13193_29093.n2016 w_13193_29093.n1964 185
R3364 w_13193_29093.n2018 w_13193_29093.n2017 185
R3365 w_13193_29093.n2020 w_13193_29093.n1963 185
R3366 w_13193_29093.n2022 w_13193_29093.n2021 185
R3367 w_13193_29093.n2024 w_13193_29093.n2023 185
R3368 w_13193_29093.n2027 w_13193_29093.n2026 185
R3369 w_13193_29093.n2028 w_13193_29093.n1936 185
R3370 w_13193_29093.n2037 w_13193_29093.n2036 185
R3371 w_13193_29093.n2039 w_13193_29093.n1935 185
R3372 w_13193_29093.n2042 w_13193_29093.n2041 185
R3373 w_13193_29093.n2043 w_13193_29093.n1931 185
R3374 w_13193_29093.n2052 w_13193_29093.n2051 185
R3375 w_13193_29093.n2054 w_13193_29093.n1930 185
R3376 w_13193_29093.n2055 w_13193_29093.n1926 185
R3377 w_13193_29093.n547 w_13193_29093.n525 185
R3378 w_13193_29093.n545 w_13193_29093.n544 185
R3379 w_13193_29093.n543 w_13193_29093.n527 185
R3380 w_13193_29093.n542 w_13193_29093.n541 185
R3381 w_13193_29093.n539 w_13193_29093.n528 185
R3382 w_13193_29093.n537 w_13193_29093.n536 185
R3383 w_13193_29093.n535 w_13193_29093.n529 185
R3384 w_13193_29093.n534 w_13193_29093.n533 185
R3385 w_13193_29093.n531 w_13193_29093.n453 185
R3386 w_13193_29093.n549 w_13193_29093.n548 185
R3387 w_13193_29093.n550 w_13193_29093.n524 185
R3388 w_13193_29093.n552 w_13193_29093.n551 185
R3389 w_13193_29093.n554 w_13193_29093.n522 185
R3390 w_13193_29093.n556 w_13193_29093.n555 185
R3391 w_13193_29093.n557 w_13193_29093.n521 185
R3392 w_13193_29093.n559 w_13193_29093.n558 185
R3393 w_13193_29093.n561 w_13193_29093.n520 185
R3394 w_13193_29093.n564 w_13193_29093.n563 185
R3395 w_13193_29093.n565 w_13193_29093.n519 185
R3396 w_13193_29093.n567 w_13193_29093.n566 185
R3397 w_13193_29093.n569 w_13193_29093.n518 185
R3398 w_13193_29093.n572 w_13193_29093.n571 185
R3399 w_13193_29093.n573 w_13193_29093.n517 185
R3400 w_13193_29093.n575 w_13193_29093.n574 185
R3401 w_13193_29093.n577 w_13193_29093.n516 185
R3402 w_13193_29093.n580 w_13193_29093.n579 185
R3403 w_13193_29093.n581 w_13193_29093.n515 185
R3404 w_13193_29093.n963 w_13193_29093.n962 185
R3405 w_13193_29093.n965 w_13193_29093.n964 185
R3406 w_13193_29093.n967 w_13193_29093.n966 185
R3407 w_13193_29093.n969 w_13193_29093.n968 185
R3408 w_13193_29093.n971 w_13193_29093.n970 185
R3409 w_13193_29093.n973 w_13193_29093.n972 185
R3410 w_13193_29093.n975 w_13193_29093.n974 185
R3411 w_13193_29093.n977 w_13193_29093.n976 185
R3412 w_13193_29093.n978 w_13193_29093.n924 185
R3413 w_13193_29093.n961 w_13193_29093.n960 185
R3414 w_13193_29093.n959 w_13193_29093.n958 185
R3415 w_13193_29093.n957 w_13193_29093.n956 185
R3416 w_13193_29093.n955 w_13193_29093.n954 185
R3417 w_13193_29093.n953 w_13193_29093.n952 185
R3418 w_13193_29093.n951 w_13193_29093.n950 185
R3419 w_13193_29093.n949 w_13193_29093.n948 185
R3420 w_13193_29093.n947 w_13193_29093.n946 185
R3421 w_13193_29093.n945 w_13193_29093.n944 185
R3422 w_13193_29093.n943 w_13193_29093.n942 185
R3423 w_13193_29093.n941 w_13193_29093.n940 185
R3424 w_13193_29093.n939 w_13193_29093.n938 185
R3425 w_13193_29093.n937 w_13193_29093.n936 185
R3426 w_13193_29093.n935 w_13193_29093.n934 185
R3427 w_13193_29093.n933 w_13193_29093.n932 185
R3428 w_13193_29093.n931 w_13193_29093.n930 185
R3429 w_13193_29093.n929 w_13193_29093.n928 185
R3430 w_13193_29093.n927 w_13193_29093.n906 185
R3431 w_13193_29093.n1020 w_13193_29093.n1019 185
R3432 w_13193_29093.n988 w_13193_29093.n907 185
R3433 w_13193_29093.n994 w_13193_29093.n993 185
R3434 w_13193_29093.n991 w_13193_29093.n990 185
R3435 w_13193_29093.n989 w_13193_29093.n984 185
R3436 w_13193_29093.n1004 w_13193_29093.n1003 185
R3437 w_13193_29093.n1006 w_13193_29093.n1005 185
R3438 w_13193_29093.n1007 w_13193_29093.n925 185
R3439 w_13193_29093.n1016 w_13193_29093.n1015 185
R3440 w_13193_29093.n1424 w_13193_29093.n1400 185
R3441 w_13193_29093.n1422 w_13193_29093.n1421 185
R3442 w_13193_29093.n1420 w_13193_29093.n1402 185
R3443 w_13193_29093.n1419 w_13193_29093.n1418 185
R3444 w_13193_29093.n1416 w_13193_29093.n1403 185
R3445 w_13193_29093.n1414 w_13193_29093.n1413 185
R3446 w_13193_29093.n1412 w_13193_29093.n1404 185
R3447 w_13193_29093.n1411 w_13193_29093.n1410 185
R3448 w_13193_29093.n1408 w_13193_29093.n1406 185
R3449 w_13193_29093.n1426 w_13193_29093.n1425 185
R3450 w_13193_29093.n1427 w_13193_29093.n1399 185
R3451 w_13193_29093.n1429 w_13193_29093.n1428 185
R3452 w_13193_29093.n1431 w_13193_29093.n1397 185
R3453 w_13193_29093.n1433 w_13193_29093.n1432 185
R3454 w_13193_29093.n1434 w_13193_29093.n1396 185
R3455 w_13193_29093.n1436 w_13193_29093.n1435 185
R3456 w_13193_29093.n1438 w_13193_29093.n1395 185
R3457 w_13193_29093.n1441 w_13193_29093.n1440 185
R3458 w_13193_29093.n1442 w_13193_29093.n1394 185
R3459 w_13193_29093.n1444 w_13193_29093.n1443 185
R3460 w_13193_29093.n1446 w_13193_29093.n1393 185
R3461 w_13193_29093.n1449 w_13193_29093.n1448 185
R3462 w_13193_29093.n1450 w_13193_29093.n1392 185
R3463 w_13193_29093.n1452 w_13193_29093.n1451 185
R3464 w_13193_29093.n1454 w_13193_29093.n1391 185
R3465 w_13193_29093.n1456 w_13193_29093.n1455 185
R3466 w_13193_29093.n1458 w_13193_29093.n1457 185
R3467 w_13193_29093.n1459 w_13193_29093.n614 185
R3468 w_13193_29093.n1462 w_13193_29093.n1461 185
R3469 w_13193_29093.n618 w_13193_29093.n617 185
R3470 w_13193_29093.n605 w_13193_29093.n602 185
R3471 w_13193_29093.n1480 w_13193_29093.n1479 185
R3472 w_13193_29093.n1482 w_13193_29093.n601 185
R3473 w_13193_29093.n1483 w_13193_29093.n596 185
R3474 w_13193_29093.n1486 w_13193_29093.n1485 185
R3475 w_13193_29093.n599 w_13193_29093.n598 185
R3476 w_13193_29093.n829 w_13193_29093.n828 185
R3477 w_13193_29093.n827 w_13193_29093.n826 185
R3478 w_13193_29093.n825 w_13193_29093.n824 185
R3479 w_13193_29093.n823 w_13193_29093.n822 185
R3480 w_13193_29093.n821 w_13193_29093.n820 185
R3481 w_13193_29093.n819 w_13193_29093.n818 185
R3482 w_13193_29093.n817 w_13193_29093.n816 185
R3483 w_13193_29093.n815 w_13193_29093.n814 185
R3484 w_13193_29093.n787 w_13193_29093.n784 185
R3485 w_13193_29093.n831 w_13193_29093.n830 185
R3486 w_13193_29093.n833 w_13193_29093.n832 185
R3487 w_13193_29093.n835 w_13193_29093.n834 185
R3488 w_13193_29093.n837 w_13193_29093.n836 185
R3489 w_13193_29093.n839 w_13193_29093.n838 185
R3490 w_13193_29093.n841 w_13193_29093.n840 185
R3491 w_13193_29093.n843 w_13193_29093.n842 185
R3492 w_13193_29093.n845 w_13193_29093.n844 185
R3493 w_13193_29093.n847 w_13193_29093.n846 185
R3494 w_13193_29093.n849 w_13193_29093.n848 185
R3495 w_13193_29093.n851 w_13193_29093.n850 185
R3496 w_13193_29093.n853 w_13193_29093.n852 185
R3497 w_13193_29093.n855 w_13193_29093.n854 185
R3498 w_13193_29093.n857 w_13193_29093.n856 185
R3499 w_13193_29093.n859 w_13193_29093.n858 185
R3500 w_13193_29093.n861 w_13193_29093.n860 185
R3501 w_13193_29093.n863 w_13193_29093.n862 185
R3502 w_13193_29093.n865 w_13193_29093.n864 185
R3503 w_13193_29093.n700 w_13193_29093.n699 185
R3504 w_13193_29093.n702 w_13193_29093.n701 185
R3505 w_13193_29093.n704 w_13193_29093.n703 185
R3506 w_13193_29093.n706 w_13193_29093.n705 185
R3507 w_13193_29093.n708 w_13193_29093.n707 185
R3508 w_13193_29093.n710 w_13193_29093.n709 185
R3509 w_13193_29093.n712 w_13193_29093.n711 185
R3510 w_13193_29093.n714 w_13193_29093.n713 185
R3511 w_13193_29093.n715 w_13193_29093.n657 185
R3512 w_13193_29093.n698 w_13193_29093.n697 185
R3513 w_13193_29093.n696 w_13193_29093.n695 185
R3514 w_13193_29093.n694 w_13193_29093.n693 185
R3515 w_13193_29093.n692 w_13193_29093.n691 185
R3516 w_13193_29093.n690 w_13193_29093.n689 185
R3517 w_13193_29093.n688 w_13193_29093.n687 185
R3518 w_13193_29093.n686 w_13193_29093.n685 185
R3519 w_13193_29093.n684 w_13193_29093.n683 185
R3520 w_13193_29093.n682 w_13193_29093.n681 185
R3521 w_13193_29093.n680 w_13193_29093.n679 185
R3522 w_13193_29093.n678 w_13193_29093.n677 185
R3523 w_13193_29093.n676 w_13193_29093.n675 185
R3524 w_13193_29093.n674 w_13193_29093.n673 185
R3525 w_13193_29093.n672 w_13193_29093.n671 185
R3526 w_13193_29093.n670 w_13193_29093.n669 185
R3527 w_13193_29093.n668 w_13193_29093.n667 185
R3528 w_13193_29093.n666 w_13193_29093.n665 185
R3529 w_13193_29093.n664 w_13193_29093.n663 185
R3530 w_13193_29093.n662 w_13193_29093.n661 185
R3531 w_13193_29093.n639 w_13193_29093.n637 185
R3532 w_13193_29093.n1156 w_13193_29093.n1155 185
R3533 w_13193_29093.n720 w_13193_29093.n640 185
R3534 w_13193_29093.n724 w_13193_29093.n723 185
R3535 w_13193_29093.n729 w_13193_29093.n726 185
R3536 w_13193_29093.n731 w_13193_29093.n730 185
R3537 w_13193_29093.n727 w_13193_29093.n658 185
R3538 w_13193_29093.n1152 w_13193_29093.n1151 185
R3539 w_13193_29093.n867 w_13193_29093.n866 185
R3540 w_13193_29093.n871 w_13193_29093.n870 185
R3541 w_13193_29093.n869 w_13193_29093.n811 185
R3542 w_13193_29093.n880 w_13193_29093.n879 185
R3543 w_13193_29093.n882 w_13193_29093.n881 185
R3544 w_13193_29093.n883 w_13193_29093.n804 185
R3545 w_13193_29093.n893 w_13193_29093.n892 185
R3546 w_13193_29093.n806 w_13193_29093.n786 185
R3547 w_13193_29093.n897 w_13193_29093.n896 185
R3548 w_13193_29093.n1551 w_13193_29093.n1550 185
R3549 w_13193_29093.n1553 w_13193_29093.n514 185
R3550 w_13193_29093.n1556 w_13193_29093.n1555 185
R3551 w_13193_29093.n1558 w_13193_29093.n512 185
R3552 w_13193_29093.n1564 w_13193_29093.n1563 185
R3553 w_13193_29093.n1566 w_13193_29093.n511 185
R3554 w_13193_29093.n1567 w_13193_29093.n507 185
R3555 w_13193_29093.n1570 w_13193_29093.n1569 185
R3556 w_13193_29093.n509 w_13193_29093.n452 185
R3557 w_13193_29093.n1262 w_13193_29093.n1244 185
R3558 w_13193_29093.n1260 w_13193_29093.n1259 185
R3559 w_13193_29093.n1258 w_13193_29093.n1246 185
R3560 w_13193_29093.n1257 w_13193_29093.n1256 185
R3561 w_13193_29093.n1254 w_13193_29093.n1247 185
R3562 w_13193_29093.n1252 w_13193_29093.n1251 185
R3563 w_13193_29093.n1250 w_13193_29093.n1249 185
R3564 w_13193_29093.n1218 w_13193_29093.n1217 185
R3565 w_13193_29093.n1330 w_13193_29093.n1329 185
R3566 w_13193_29093.n1264 w_13193_29093.n1263 185
R3567 w_13193_29093.n1265 w_13193_29093.n1243 185
R3568 w_13193_29093.n1267 w_13193_29093.n1266 185
R3569 w_13193_29093.n1269 w_13193_29093.n1241 185
R3570 w_13193_29093.n1271 w_13193_29093.n1270 185
R3571 w_13193_29093.n1272 w_13193_29093.n1240 185
R3572 w_13193_29093.n1274 w_13193_29093.n1273 185
R3573 w_13193_29093.n1276 w_13193_29093.n1239 185
R3574 w_13193_29093.n1279 w_13193_29093.n1278 185
R3575 w_13193_29093.n1280 w_13193_29093.n1238 185
R3576 w_13193_29093.n1282 w_13193_29093.n1281 185
R3577 w_13193_29093.n1284 w_13193_29093.n1237 185
R3578 w_13193_29093.n1287 w_13193_29093.n1286 185
R3579 w_13193_29093.n1288 w_13193_29093.n1236 185
R3580 w_13193_29093.n1290 w_13193_29093.n1289 185
R3581 w_13193_29093.n1292 w_13193_29093.n1235 185
R3582 w_13193_29093.n1294 w_13193_29093.n1293 185
R3583 w_13193_29093.n1296 w_13193_29093.n1295 185
R3584 w_13193_29093.n1299 w_13193_29093.n1298 185
R3585 w_13193_29093.n1300 w_13193_29093.n1226 185
R3586 w_13193_29093.n1309 w_13193_29093.n1308 185
R3587 w_13193_29093.n1311 w_13193_29093.n1225 185
R3588 w_13193_29093.n1314 w_13193_29093.n1313 185
R3589 w_13193_29093.n1315 w_13193_29093.n1221 185
R3590 w_13193_29093.n1324 w_13193_29093.n1323 185
R3591 w_13193_29093.n1326 w_13193_29093.n1220 185
R3592 w_13193_29093.n1327 w_13193_29093.n1216 185
R3593 w_13193_29093.n1903 w_13193_29093.n1902 185
R3594 w_13193_29093.n1905 w_13193_29093.n333 185
R3595 w_13193_29093.n1906 w_13193_29093.n329 185
R3596 w_13193_29093.n1909 w_13193_29093.n1908 185
R3597 w_13193_29093.n367 w_13193_29093.n331 185
R3598 w_13193_29093.n372 w_13193_29093.n370 185
R3599 w_13193_29093.n375 w_13193_29093.n374 185
R3600 w_13193_29093.n376 w_13193_29093.n350 185
R3601 w_13193_29093.n1846 w_13193_29093.n1845 185
R3602 w_13193_29093.n1666 w_13193_29093.n1665 185
R3603 w_13193_29093.n1668 w_13193_29093.n485 185
R3604 w_13193_29093.n1669 w_13193_29093.n476 185
R3605 w_13193_29093.n1672 w_13193_29093.n1671 185
R3606 w_13193_29093.n483 w_13193_29093.n482 185
R3607 w_13193_29093.n479 w_13193_29093.n465 185
R3608 w_13193_29093.n1688 w_13193_29093.n1687 185
R3609 w_13193_29093.n1690 w_13193_29093.n464 185
R3610 w_13193_29093.n1691 w_13193_29093.n460 185
R3611 w_13193_29093.n2187 w_13193_29093.n2185 175.546
R3612 w_13193_29093.n2191 w_13193_29093.n270 175.546
R3613 w_13193_29093.n2194 w_13193_29093.n2193 175.546
R3614 w_13193_29093.n2196 w_13193_29093.n268 175.546
R3615 w_13193_29093.n1810 w_13193_29093.n1809 175.546
R3616 w_13193_29093.n1811 w_13193_29093.n1810 175.546
R3617 w_13193_29093.n1836 w_13193_29093.n1835 175.546
R3618 w_13193_29093.n1833 w_13193_29093.n389 175.546
R3619 w_13193_29093.n1829 w_13193_29093.n1828 175.546
R3620 w_13193_29093.n1826 w_13193_29093.n398 175.546
R3621 w_13193_29093.n1822 w_13193_29093.n1821 175.546
R3622 w_13193_29093.n1819 w_13193_29093.n407 175.546
R3623 w_13193_29093.n1921 w_13193_29093.n320 175.546
R3624 w_13193_29093.n1900 w_13193_29093.n320 175.546
R3625 w_13193_29093.n1900 w_13193_29093.n327 175.546
R3626 w_13193_29093.n1911 w_13193_29093.n327 175.546
R3627 w_13193_29093.n1911 w_13193_29093.n328 175.546
R3628 w_13193_29093.n368 w_13193_29093.n328 175.546
R3629 w_13193_29093.n368 w_13193_29093.n365 175.546
R3630 w_13193_29093.n378 w_13193_29093.n365 175.546
R3631 w_13193_29093.n378 w_13193_29093.n353 175.546
R3632 w_13193_29093.n1843 w_13193_29093.n353 175.546
R3633 w_13193_29093.n1843 w_13193_29093.n354 175.546
R3634 w_13193_29093.n2066 w_13193_29093.n318 175.546
R3635 w_13193_29093.n2069 w_13193_29093.n2068 175.546
R3636 w_13193_29093.n2075 w_13193_29093.n2071 175.546
R3637 w_13193_29093.n2078 w_13193_29093.n2077 175.546
R3638 w_13193_29093.n2084 w_13193_29093.n2080 175.546
R3639 w_13193_29093.n2087 w_13193_29093.n2086 175.546
R3640 w_13193_29093.n1956 w_13193_29093.n1955 175.546
R3641 w_13193_29093.n1952 w_13193_29093.n1951 175.546
R3642 w_13193_29093.n1948 w_13193_29093.n1947 175.546
R3643 w_13193_29093.n1944 w_13193_29093.n1943 175.546
R3644 w_13193_29093.n2155 w_13193_29093.n284 175.546
R3645 w_13193_29093.n2030 w_13193_29093.n1938 175.546
R3646 w_13193_29093.n2034 w_13193_29093.n2032 175.546
R3647 w_13193_29093.n2045 w_13193_29093.n1933 175.546
R3648 w_13193_29093.n2049 w_13193_29093.n2047 175.546
R3649 w_13193_29093.n2061 w_13193_29093.n1925 175.546
R3650 w_13193_29093.n2106 w_13193_29093.n2105 175.546
R3651 w_13193_29093.n2103 w_13193_29093.n2065 175.546
R3652 w_13193_29093.n2099 w_13193_29093.n2098 175.546
R3653 w_13193_29093.n2096 w_13193_29093.n2074 175.546
R3654 w_13193_29093.n2092 w_13193_29093.n2091 175.546
R3655 w_13193_29093.n2089 w_13193_29093.n2083 175.546
R3656 w_13193_29093.n2163 w_13193_29093.n2161 175.546
R3657 w_13193_29093.n2167 w_13193_29093.n280 175.546
R3658 w_13193_29093.n2171 w_13193_29093.n2169 175.546
R3659 w_13193_29093.n2175 w_13193_29093.n278 175.546
R3660 w_13193_29093.n2178 w_13193_29093.n2177 175.546
R3661 w_13193_29093.n390 w_13193_29093.n385 175.546
R3662 w_13193_29093.n393 w_13193_29093.n392 175.546
R3663 w_13193_29093.n399 w_13193_29093.n395 175.546
R3664 w_13193_29093.n402 w_13193_29093.n401 175.546
R3665 w_13193_29093.n408 w_13193_29093.n404 175.546
R3666 w_13193_29093.n411 w_13193_29093.n410 175.546
R3667 w_13193_29093.n1654 w_13193_29093.n488 175.546
R3668 w_13193_29093.n1663 w_13193_29093.n488 175.546
R3669 w_13193_29093.n1663 w_13193_29093.n474 175.546
R3670 w_13193_29093.n1674 w_13193_29093.n474 175.546
R3671 w_13193_29093.n1674 w_13193_29093.n475 175.546
R3672 w_13193_29093.n480 w_13193_29093.n475 175.546
R3673 w_13193_29093.n480 w_13193_29093.n467 175.546
R3674 w_13193_29093.n1685 w_13193_29093.n467 175.546
R3675 w_13193_29093.n1685 w_13193_29093.n458 175.546
R3676 w_13193_29093.n1716 w_13193_29093.n458 175.546
R3677 w_13193_29093.n1716 w_13193_29093.n459 175.546
R3678 w_13193_29093.n1710 w_13193_29093.n1709 175.546
R3679 w_13193_29093.n1706 w_13193_29093.n1705 175.546
R3680 w_13193_29093.n1702 w_13193_29093.n1701 175.546
R3681 w_13193_29093.n1698 w_13193_29093.n1697 175.546
R3682 w_13193_29093.n1778 w_13193_29093.n424 175.546
R3683 w_13193_29093.n1799 w_13193_29093.n1798 175.546
R3684 w_13193_29093.n1796 w_13193_29093.n416 175.546
R3685 w_13193_29093.n1792 w_13193_29093.n1791 175.546
R3686 w_13193_29093.n1789 w_13193_29093.n419 175.546
R3687 w_13193_29093.n1785 w_13193_29093.n1784 175.546
R3688 w_13193_29093.n1163 w_13193_29093.n1162 175.546
R3689 w_13193_29093.n1162 w_13193_29093.n633 175.546
R3690 w_13193_29093.n1158 w_13193_29093.n633 175.546
R3691 w_13193_29093.n1158 w_13193_29093.n636 175.546
R3692 w_13193_29093.n721 w_13193_29093.n636 175.546
R3693 w_13193_29093.n721 w_13193_29093.n719 175.546
R3694 w_13193_29093.n733 w_13193_29093.n719 175.546
R3695 w_13193_29093.n733 w_13193_29093.n717 175.546
R3696 w_13193_29093.n737 w_13193_29093.n717 175.546
R3697 w_13193_29093.n1149 w_13193_29093.n737 175.546
R3698 w_13193_29093.n1149 w_13193_29093.n738 175.546
R3699 w_13193_29093.n1168 w_13193_29093.n1167 175.546
R3700 w_13193_29093.n1172 w_13193_29093.n1171 175.546
R3701 w_13193_29093.n1176 w_13193_29093.n1175 175.546
R3702 w_13193_29093.n1180 w_13193_29093.n1179 175.546
R3703 w_13193_29093.n1184 w_13193_29093.n1183 175.546
R3704 w_13193_29093.n1193 w_13193_29093.n630 175.546
R3705 w_13193_29093.n1197 w_13193_29093.n1195 175.546
R3706 w_13193_29093.n1201 w_13193_29093.n628 175.546
R3707 w_13193_29093.n1205 w_13193_29093.n1203 175.546
R3708 w_13193_29093.n1209 w_13193_29093.n626 175.546
R3709 w_13193_29093.n1145 w_13193_29093.n739 175.546
R3710 w_13193_29093.n1140 w_13193_29093.n1139 175.546
R3711 w_13193_29093.n1137 w_13193_29093.n1106 175.546
R3712 w_13193_29093.n1133 w_13193_29093.n1132 175.546
R3713 w_13193_29093.n1130 w_13193_29093.n1115 175.546
R3714 w_13193_29093.n1126 w_13193_29093.n1125 175.546
R3715 w_13193_29093.n1027 w_13193_29093.n1026 175.546
R3716 w_13193_29093.n1033 w_13193_29093.n1032 175.546
R3717 w_13193_29093.n1036 w_13193_29093.n1035 175.546
R3718 w_13193_29093.n1042 w_13193_29093.n1038 175.546
R3719 w_13193_29093.n1045 w_13193_29093.n1044 175.546
R3720 w_13193_29093.n1049 w_13193_29093.n1047 175.546
R3721 w_13193_29093.n1022 w_13193_29093.n902 175.546
R3722 w_13193_29093.n1022 w_13193_29093.n903 175.546
R3723 w_13193_29093.n996 w_13193_29093.n903 175.546
R3724 w_13193_29093.n996 w_13193_29093.n985 175.546
R3725 w_13193_29093.n1000 w_13193_29093.n985 175.546
R3726 w_13193_29093.n1001 w_13193_29093.n1000 175.546
R3727 w_13193_29093.n1001 w_13193_29093.n982 175.546
R3728 w_13193_29093.n1009 w_13193_29093.n982 175.546
R3729 w_13193_29093.n1009 w_13193_29093.n980 175.546
R3730 w_13193_29093.n1013 w_13193_29093.n980 175.546
R3731 w_13193_29093.n1013 w_13193_29093.n444 175.546
R3732 w_13193_29093.n1771 w_13193_29093.n1770 175.546
R3733 w_13193_29093.n1767 w_13193_29093.n1766 175.546
R3734 w_13193_29093.n1763 w_13193_29093.n1762 175.546
R3735 w_13193_29093.n1759 w_13193_29093.n1758 175.546
R3736 w_13193_29093.n1755 w_13193_29093.n1754 175.546
R3737 w_13193_29093.n1588 w_13193_29093.n494 175.546
R3738 w_13193_29093.n1584 w_13193_29093.n494 175.546
R3739 w_13193_29093.n1584 w_13193_29093.n497 175.546
R3740 w_13193_29093.n1580 w_13193_29093.n497 175.546
R3741 w_13193_29093.n1580 w_13193_29093.n501 175.546
R3742 w_13193_29093.n1576 w_13193_29093.n501 175.546
R3743 w_13193_29093.n1576 w_13193_29093.n1575 175.546
R3744 w_13193_29093.n1575 w_13193_29093.n505 175.546
R3745 w_13193_29093.n505 w_13193_29093.n447 175.546
R3746 w_13193_29093.n1749 w_13193_29093.n447 175.546
R3747 w_13193_29093.n1750 w_13193_29093.n1749 175.546
R3748 w_13193_29093.n585 w_13193_29093.n584 175.546
R3749 w_13193_29093.n1504 w_13193_29093.n1503 175.546
R3750 w_13193_29093.n1507 w_13193_29093.n1506 175.546
R3751 w_13193_29093.n1513 w_13193_29093.n1509 175.546
R3752 w_13193_29093.n1516 w_13193_29093.n1515 175.546
R3753 w_13193_29093.n1520 w_13193_29093.n1518 175.546
R3754 w_13193_29093.n1547 w_13193_29093.n491 175.546
R3755 w_13193_29093.n1547 w_13193_29093.n498 175.546
R3756 w_13193_29093.n499 w_13193_29093.n498 175.546
R3757 w_13193_29093.n500 w_13193_29093.n499 175.546
R3758 w_13193_29093.n1560 w_13193_29093.n500 175.546
R3759 w_13193_29093.n1561 w_13193_29093.n1560 175.546
R3760 w_13193_29093.n1561 w_13193_29093.n506 175.546
R3761 w_13193_29093.n1572 w_13193_29093.n506 175.546
R3762 w_13193_29093.n1572 w_13193_29093.n450 175.546
R3763 w_13193_29093.n1747 w_13193_29093.n450 175.546
R3764 w_13193_29093.n1747 w_13193_29093.n451 175.546
R3765 w_13193_29093.n1740 w_13193_29093.n454 175.546
R3766 w_13193_29093.n1738 w_13193_29093.n1737 175.546
R3767 w_13193_29093.n1734 w_13193_29093.n1733 175.546
R3768 w_13193_29093.n1730 w_13193_29093.n1729 175.546
R3769 w_13193_29093.n1726 w_13193_29093.n1725 175.546
R3770 w_13193_29093.n1722 w_13193_29093.n431 175.546
R3771 w_13193_29093.n1657 w_13193_29093.n1656 175.546
R3772 w_13193_29093.n1661 w_13193_29093.n1657 175.546
R3773 w_13193_29093.n1661 w_13193_29093.n471 175.546
R3774 w_13193_29093.n1676 w_13193_29093.n471 175.546
R3775 w_13193_29093.n1677 w_13193_29093.n1676 175.546
R3776 w_13193_29093.n1678 w_13193_29093.n1677 175.546
R3777 w_13193_29093.n1678 w_13193_29093.n469 175.546
R3778 w_13193_29093.n1683 w_13193_29093.n469 175.546
R3779 w_13193_29093.n1683 w_13193_29093.n456 175.546
R3780 w_13193_29093.n1718 w_13193_29093.n456 175.546
R3781 w_13193_29093.n1719 w_13193_29093.n1718 175.546
R3782 w_13193_29093.n1338 w_13193_29093.n621 175.546
R3783 w_13193_29093.n1341 w_13193_29093.n1340 175.546
R3784 w_13193_29093.n1347 w_13193_29093.n1343 175.546
R3785 w_13193_29093.n1350 w_13193_29093.n1349 175.546
R3786 w_13193_29093.n1357 w_13193_29093.n1352 175.546
R3787 w_13193_29093.n1361 w_13193_29093.n1359 175.546
R3788 w_13193_29093.n1919 w_13193_29093.n1918 175.546
R3789 w_13193_29093.n1918 w_13193_29093.n323 175.546
R3790 w_13193_29093.n1914 w_13193_29093.n323 175.546
R3791 w_13193_29093.n1914 w_13193_29093.n325 175.546
R3792 w_13193_29093.n359 w_13193_29093.n325 175.546
R3793 w_13193_29093.n362 w_13193_29093.n359 175.546
R3794 w_13193_29093.n363 w_13193_29093.n362 175.546
R3795 w_13193_29093.n380 w_13193_29093.n363 175.546
R3796 w_13193_29093.n380 w_13193_29093.n356 175.546
R3797 w_13193_29093.n1841 w_13193_29093.n356 175.546
R3798 w_13193_29093.n1841 w_13193_29093.n357 175.546
R3799 w_13193_29093.n1542 w_13193_29093.n1499 175.546
R3800 w_13193_29093.n1540 w_13193_29093.n1539 175.546
R3801 w_13193_29093.n1537 w_13193_29093.n1501 175.546
R3802 w_13193_29093.n1533 w_13193_29093.n1532 175.546
R3803 w_13193_29093.n1530 w_13193_29093.n1512 175.546
R3804 w_13193_29093.n1526 w_13193_29093.n1525 175.546
R3805 w_13193_29093.n1387 w_13193_29093.n613 175.546
R3806 w_13193_29093.n1464 w_13193_29093.n613 175.546
R3807 w_13193_29093.n1464 w_13193_29093.n604 175.546
R3808 w_13193_29093.n1475 w_13193_29093.n604 175.546
R3809 w_13193_29093.n1476 w_13193_29093.n1475 175.546
R3810 w_13193_29093.n1477 w_13193_29093.n1476 175.546
R3811 w_13193_29093.n1477 w_13193_29093.n595 175.546
R3812 w_13193_29093.n1488 w_13193_29093.n595 175.546
R3813 w_13193_29093.n1488 w_13193_29093.n587 175.546
R3814 w_13193_29093.n1497 w_13193_29093.n587 175.546
R3815 w_13193_29093.n1498 w_13193_29093.n1497 175.546
R3816 w_13193_29093.n1101 w_13193_29093.n740 175.546
R3817 w_13193_29093.n1107 w_13193_29093.n1103 175.546
R3818 w_13193_29093.n1110 w_13193_29093.n1109 175.546
R3819 w_13193_29093.n1116 w_13193_29093.n1112 175.546
R3820 w_13193_29093.n1119 w_13193_29093.n1118 175.546
R3821 w_13193_29093.n1123 w_13193_29093.n1122 175.546
R3822 w_13193_29093.n1099 w_13193_29093.n743 175.546
R3823 w_13193_29093.n873 w_13193_29093.n743 175.546
R3824 w_13193_29093.n873 w_13193_29093.n812 175.546
R3825 w_13193_29093.n877 w_13193_29093.n812 175.546
R3826 w_13193_29093.n877 w_13193_29093.n809 175.546
R3827 w_13193_29093.n885 w_13193_29093.n809 175.546
R3828 w_13193_29093.n885 w_13193_29093.n807 175.546
R3829 w_13193_29093.n890 w_13193_29093.n807 175.546
R3830 w_13193_29093.n890 w_13193_29093.n808 175.546
R3831 w_13193_29093.n808 w_13193_29093.n782 175.546
R3832 w_13193_29093.n1076 w_13193_29093.n782 175.546
R3833 w_13193_29093.n1072 w_13193_29093.n783 175.546
R3834 w_13193_29093.n1070 w_13193_29093.n1069 175.546
R3835 w_13193_29093.n1067 w_13193_29093.n1030 175.546
R3836 w_13193_29093.n1063 w_13193_29093.n1062 175.546
R3837 w_13193_29093.n1060 w_13193_29093.n1041 175.546
R3838 w_13193_29093.n1056 w_13193_29093.n1055 175.546
R3839 w_13193_29093.n1385 w_13193_29093.n611 175.546
R3840 w_13193_29093.n1466 w_13193_29093.n611 175.546
R3841 w_13193_29093.n1466 w_13193_29093.n608 175.546
R3842 w_13193_29093.n1473 w_13193_29093.n608 175.546
R3843 w_13193_29093.n1473 w_13193_29093.n609 175.546
R3844 w_13193_29093.n1469 w_13193_29093.n609 175.546
R3845 w_13193_29093.n1469 w_13193_29093.n593 175.546
R3846 w_13193_29093.n1490 w_13193_29093.n593 175.546
R3847 w_13193_29093.n1490 w_13193_29093.n590 175.546
R3848 w_13193_29093.n1495 w_13193_29093.n590 175.546
R3849 w_13193_29093.n1495 w_13193_29093.n591 175.546
R3850 w_13193_29093.n2127 w_13193_29093.n2126 175.546
R3851 w_13193_29093.n2124 w_13193_29093.n309 175.546
R3852 w_13193_29093.n2120 w_13193_29093.n2119 175.546
R3853 w_13193_29093.n2117 w_13193_29093.n312 175.546
R3854 w_13193_29093.n2113 w_13193_29093.n2112 175.546
R3855 w_13193_29093.n1381 w_13193_29093.n1380 175.546
R3856 w_13193_29093.n1378 w_13193_29093.n1337 175.546
R3857 w_13193_29093.n1374 w_13193_29093.n1373 175.546
R3858 w_13193_29093.n1371 w_13193_29093.n1346 175.546
R3859 w_13193_29093.n1367 w_13193_29093.n1366 175.546
R3860 w_13193_29093.n1364 w_13193_29093.n1356 175.546
R3861 w_13193_29093.n1302 w_13193_29093.n1228 175.546
R3862 w_13193_29093.n1306 w_13193_29093.n1304 175.546
R3863 w_13193_29093.n1317 w_13193_29093.n1223 175.546
R3864 w_13193_29093.n1321 w_13193_29093.n1319 175.546
R3865 w_13193_29093.n1333 w_13193_29093.n1215 175.546
R3866 w_13193_29093.n2152 w_13193_29093.n2151 175.546
R3867 w_13193_29093.n2148 w_13193_29093.n2147 175.546
R3868 w_13193_29093.n2144 w_13193_29093.n2143 175.546
R3869 w_13193_29093.n2140 w_13193_29093.n2139 175.546
R3870 w_13193_29093.n2136 w_13193_29093.n2135 175.546
R3871 w_13193_29093.n2132 w_13193_29093.n298 175.546
R3872 w_13193_29093.t56 w_13193_29093.n222 174.089
R3873 w_13193_29093.n228 w_13193_29093.t56 174.089
R3874 w_13193_29093.n2505 w_13193_29093.t72 174.089
R3875 w_13193_29093.t72 w_13193_29093.n2504 174.089
R3876 w_13193_29093.t81 w_13193_29093.n2527 173.506
R3877 w_13193_29093.n2528 w_13193_29093.t81 173.506
R3878 w_13193_29093.t88 w_13193_29093.n2384 173.506
R3879 w_13193_29093.n2385 w_13193_29093.t88 173.506
R3880 w_13193_29093.t53 w_13193_29093.n19 173.084
R3881 w_13193_29093.t53 w_13193_29093.n18 173.084
R3882 w_13193_29093.n2555 w_13193_29093.n201 172.888
R3883 w_13193_29093.t53 w_13193_29093.n22 172.302
R3884 w_13193_29093.t53 w_13193_29093.n26 172.302
R3885 w_13193_29093.n227 w_13193_29093.n225 166.63
R3886 w_13193_29093.n2499 w_13193_29093.n2498 166.63
R3887 w_13193_29093.t187 w_13193_29093.t238 166.487
R3888 w_13193_29093.t289 w_13193_29093.t124 166.487
R3889 w_13193_29093.t291 w_13193_29093.t246 166.487
R3890 w_13193_29093.t48 w_13193_29093.t240 166.487
R3891 w_13193_29093.n1666 w_13193_29093.n486 163.333
R3892 w_13193_29093.n1903 w_13193_29093.n1898 163.333
R3893 w_13193_29093.n2026 w_13193_29093.n2024 163.333
R3894 w_13193_29093.n1551 w_13193_29093.n515 163.333
R3895 w_13193_29093.n1019 w_13193_29093.n906 163.333
R3896 w_13193_29093.n1459 w_13193_29093.n1458 163.333
R3897 w_13193_29093.n866 w_13193_29093.n865 163.333
R3898 w_13193_29093.n663 w_13193_29093.n662 163.333
R3899 w_13193_29093.n1298 w_13193_29093.n1296 163.333
R3900 w_13193_29093.t101 w_13193_29093.t272 163.281
R3901 w_13193_29093.n2201 w_13193_29093.n2200 157.601
R3902 w_13193_29093.t9 w_13193_29093.n2437 154.595
R3903 w_13193_29093.n2436 w_13193_29093.t187 154.595
R3904 w_13193_29093.t240 w_13193_29093.n2435 154.595
R3905 w_13193_29093.n1941 w_13193_29093.n303 152.643
R3906 w_13193_29093.n1695 w_13193_29093.n432 152.643
R3907 w_13193_29093.n631 w_13193_29093.n286 152.643
R3908 w_13193_29093.n1774 w_13193_29093.n443 152.643
R3909 w_13193_29093.n264 w_13193_29093.t244 151.275
R3910 w_13193_29093.n2210 w_13193_29093.t26 151.153
R3911 w_13193_29093.n2209 w_13193_29093.t179 150.885
R3912 w_13193_29093.n264 w_13193_29093.t297 150.817
R3913 w_13193_29093.n1669 w_13193_29093.n1668 150
R3914 w_13193_29093.n1671 w_13193_29093.n483 150
R3915 w_13193_29093.n1688 w_13193_29093.n465 150
R3916 w_13193_29093.n1691 w_13193_29093.n1690 150
R3917 w_13193_29093.n1649 w_13193_29093.n1647 150
R3918 w_13193_29093.n1645 w_13193_29093.n1591 150
R3919 w_13193_29093.n1641 w_13193_29093.n1639 150
R3920 w_13193_29093.n1637 w_13193_29093.n1593 150
R3921 w_13193_29093.n1633 w_13193_29093.n1631 150
R3922 w_13193_29093.n1629 w_13193_29093.n1595 150
R3923 w_13193_29093.n1625 w_13193_29093.n1624 150
R3924 w_13193_29093.n1622 w_13193_29093.n1598 150
R3925 w_13193_29093.n1693 w_13193_29093.n462 150
R3926 w_13193_29093.n1607 w_13193_29093.n1604 150
R3927 w_13193_29093.n1611 w_13193_29093.n1609 150
R3928 w_13193_29093.n1615 w_13193_29093.n1601 150
R3929 w_13193_29093.n1906 w_13193_29093.n1905 150
R3930 w_13193_29093.n1908 w_13193_29093.n331 150
R3931 w_13193_29093.n374 w_13193_29093.n372 150
R3932 w_13193_29093.n1846 w_13193_29093.n350 150
R3933 w_13193_29093.n1895 w_13193_29093.n1894 150
R3934 w_13193_29093.n1892 w_13193_29093.n336 150
R3935 w_13193_29093.n1888 w_13193_29093.n1886 150
R3936 w_13193_29093.n1884 w_13193_29093.n338 150
R3937 w_13193_29093.n1880 w_13193_29093.n1878 150
R3938 w_13193_29093.n1876 w_13193_29093.n340 150
R3939 w_13193_29093.n1872 w_13193_29093.n1871 150
R3940 w_13193_29093.n1869 w_13193_29093.n343 150
R3941 w_13193_29093.n1850 w_13193_29093.n1848 150
R3942 w_13193_29093.n1854 w_13193_29093.n348 150
R3943 w_13193_29093.n1858 w_13193_29093.n1856 150
R3944 w_13193_29093.n1862 w_13193_29093.n346 150
R3945 w_13193_29093.n2037 w_13193_29093.n1936 150
R3946 w_13193_29093.n2041 w_13193_29093.n2039 150
R3947 w_13193_29093.n2052 w_13193_29093.n1931 150
R3948 w_13193_29093.n2055 w_13193_29093.n2054 150
R3949 w_13193_29093.n2021 w_13193_29093.n2020 150
R3950 w_13193_29093.n2018 w_13193_29093.n1964 150
R3951 w_13193_29093.n2014 w_13193_29093.n2012 150
R3952 w_13193_29093.n2010 w_13193_29093.n1966 150
R3953 w_13193_29093.n2006 w_13193_29093.n2004 150
R3954 w_13193_29093.n2002 w_13193_29093.n1968 150
R3955 w_13193_29093.n1998 w_13193_29093.n1997 150
R3956 w_13193_29093.n1995 w_13193_29093.n1971 150
R3957 w_13193_29093.n2057 w_13193_29093.n1928 150
R3958 w_13193_29093.n1980 w_13193_29093.n1977 150
R3959 w_13193_29093.n1984 w_13193_29093.n1982 150
R3960 w_13193_29093.n1988 w_13193_29093.n1974 150
R3961 w_13193_29093.n1555 w_13193_29093.n1553 150
R3962 w_13193_29093.n1564 w_13193_29093.n512 150
R3963 w_13193_29093.n1567 w_13193_29093.n1566 150
R3964 w_13193_29093.n1569 w_13193_29093.n509 150
R3965 w_13193_29093.n579 w_13193_29093.n577 150
R3966 w_13193_29093.n575 w_13193_29093.n517 150
R3967 w_13193_29093.n571 w_13193_29093.n569 150
R3968 w_13193_29093.n567 w_13193_29093.n519 150
R3969 w_13193_29093.n563 w_13193_29093.n561 150
R3970 w_13193_29093.n559 w_13193_29093.n521 150
R3971 w_13193_29093.n555 w_13193_29093.n554 150
R3972 w_13193_29093.n552 w_13193_29093.n524 150
R3973 w_13193_29093.n533 w_13193_29093.n531 150
R3974 w_13193_29093.n537 w_13193_29093.n529 150
R3975 w_13193_29093.n541 w_13193_29093.n539 150
R3976 w_13193_29093.n545 w_13193_29093.n527 150
R3977 w_13193_29093.n993 w_13193_29093.n907 150
R3978 w_13193_29093.n990 w_13193_29093.n989 150
R3979 w_13193_29093.n1005 w_13193_29093.n1004 150
R3980 w_13193_29093.n1016 w_13193_29093.n925 150
R3981 w_13193_29093.n930 w_13193_29093.n929 150
R3982 w_13193_29093.n934 w_13193_29093.n933 150
R3983 w_13193_29093.n938 w_13193_29093.n937 150
R3984 w_13193_29093.n942 w_13193_29093.n941 150
R3985 w_13193_29093.n946 w_13193_29093.n945 150
R3986 w_13193_29093.n950 w_13193_29093.n949 150
R3987 w_13193_29093.n954 w_13193_29093.n953 150
R3988 w_13193_29093.n958 w_13193_29093.n957 150
R3989 w_13193_29093.n976 w_13193_29093.n924 150
R3990 w_13193_29093.n974 w_13193_29093.n973 150
R3991 w_13193_29093.n970 w_13193_29093.n969 150
R3992 w_13193_29093.n966 w_13193_29093.n965 150
R3993 w_13193_29093.n1461 w_13193_29093.n618 150
R3994 w_13193_29093.n1480 w_13193_29093.n602 150
R3995 w_13193_29093.n1483 w_13193_29093.n1482 150
R3996 w_13193_29093.n1485 w_13193_29093.n599 150
R3997 w_13193_29093.n1455 w_13193_29093.n1454 150
R3998 w_13193_29093.n1452 w_13193_29093.n1392 150
R3999 w_13193_29093.n1448 w_13193_29093.n1446 150
R4000 w_13193_29093.n1444 w_13193_29093.n1394 150
R4001 w_13193_29093.n1440 w_13193_29093.n1438 150
R4002 w_13193_29093.n1436 w_13193_29093.n1396 150
R4003 w_13193_29093.n1432 w_13193_29093.n1431 150
R4004 w_13193_29093.n1429 w_13193_29093.n1399 150
R4005 w_13193_29093.n1410 w_13193_29093.n1408 150
R4006 w_13193_29093.n1414 w_13193_29093.n1404 150
R4007 w_13193_29093.n1418 w_13193_29093.n1416 150
R4008 w_13193_29093.n1422 w_13193_29093.n1402 150
R4009 w_13193_29093.n870 w_13193_29093.n869 150
R4010 w_13193_29093.n881 w_13193_29093.n880 150
R4011 w_13193_29093.n893 w_13193_29093.n804 150
R4012 w_13193_29093.n896 w_13193_29093.n786 150
R4013 w_13193_29093.n862 w_13193_29093.n861 150
R4014 w_13193_29093.n858 w_13193_29093.n857 150
R4015 w_13193_29093.n854 w_13193_29093.n853 150
R4016 w_13193_29093.n850 w_13193_29093.n849 150
R4017 w_13193_29093.n846 w_13193_29093.n845 150
R4018 w_13193_29093.n842 w_13193_29093.n841 150
R4019 w_13193_29093.n838 w_13193_29093.n837 150
R4020 w_13193_29093.n834 w_13193_29093.n833 150
R4021 w_13193_29093.n814 w_13193_29093.n787 150
R4022 w_13193_29093.n818 w_13193_29093.n817 150
R4023 w_13193_29093.n822 w_13193_29093.n821 150
R4024 w_13193_29093.n826 w_13193_29093.n825 150
R4025 w_13193_29093.n1155 w_13193_29093.n639 150
R4026 w_13193_29093.n723 w_13193_29093.n640 150
R4027 w_13193_29093.n730 w_13193_29093.n729 150
R4028 w_13193_29093.n1152 w_13193_29093.n658 150
R4029 w_13193_29093.n667 w_13193_29093.n666 150
R4030 w_13193_29093.n671 w_13193_29093.n670 150
R4031 w_13193_29093.n675 w_13193_29093.n674 150
R4032 w_13193_29093.n679 w_13193_29093.n678 150
R4033 w_13193_29093.n683 w_13193_29093.n682 150
R4034 w_13193_29093.n687 w_13193_29093.n686 150
R4035 w_13193_29093.n691 w_13193_29093.n690 150
R4036 w_13193_29093.n695 w_13193_29093.n694 150
R4037 w_13193_29093.n713 w_13193_29093.n657 150
R4038 w_13193_29093.n711 w_13193_29093.n710 150
R4039 w_13193_29093.n707 w_13193_29093.n706 150
R4040 w_13193_29093.n703 w_13193_29093.n702 150
R4041 w_13193_29093.n1309 w_13193_29093.n1226 150
R4042 w_13193_29093.n1313 w_13193_29093.n1311 150
R4043 w_13193_29093.n1324 w_13193_29093.n1221 150
R4044 w_13193_29093.n1327 w_13193_29093.n1326 150
R4045 w_13193_29093.n1293 w_13193_29093.n1292 150
R4046 w_13193_29093.n1290 w_13193_29093.n1236 150
R4047 w_13193_29093.n1286 w_13193_29093.n1284 150
R4048 w_13193_29093.n1282 w_13193_29093.n1238 150
R4049 w_13193_29093.n1278 w_13193_29093.n1276 150
R4050 w_13193_29093.n1274 w_13193_29093.n1240 150
R4051 w_13193_29093.n1270 w_13193_29093.n1269 150
R4052 w_13193_29093.n1267 w_13193_29093.n1243 150
R4053 w_13193_29093.n1329 w_13193_29093.n1218 150
R4054 w_13193_29093.n1252 w_13193_29093.n1249 150
R4055 w_13193_29093.n1256 w_13193_29093.n1254 150
R4056 w_13193_29093.n1260 w_13193_29093.n1246 150
R4057 w_13193_29093.n2388 w_13193_29093.t189 146.095
R4058 w_13193_29093.n204 w_13193_29093.t276 146.095
R4059 w_13193_29093.t304 w_13193_29093.n2532 146.095
R4060 w_13193_29093.n1098 w_13193_29093.n24 146.041
R4061 w_13193_29093.n1921 w_13193_29093.n318 144.338
R4062 w_13193_29093.n1960 w_13193_29093.n304 144.338
R4063 w_13193_29093.n1654 w_13193_29093.n385 144.338
R4064 w_13193_29093.n1163 w_13193_29093.n285 144.338
R4065 w_13193_29093.n1026 w_13193_29093.n902 144.338
R4066 w_13193_29093.n584 w_13193_29093.n491 144.338
R4067 w_13193_29093.n1387 w_13193_29093.n621 144.338
R4068 w_13193_29093.n1099 w_13193_29093.n740 144.338
R4069 w_13193_29093.n1232 w_13193_29093.n292 144.338
R4070 w_13193_29093.n1077 w_13193_29093.n15 138.81
R4071 w_13193_29093.n1836 w_13193_29093.n354 136.536
R4072 w_13193_29093.n2106 w_13193_29093.n2063 136.536
R4073 w_13193_29093.n459 w_13193_29093.n437 136.536
R4074 w_13193_29093.n1145 w_13193_29093.n738 136.536
R4075 w_13193_29093.n1775 w_13193_29093.n444 136.536
R4076 w_13193_29093.n1742 w_13193_29093.n451 136.536
R4077 w_13193_29093.n1499 w_13193_29093.n1498 136.536
R4078 w_13193_29093.n1076 w_13193_29093.n783 136.536
R4079 w_13193_29093.n1381 w_13193_29093.n1335 136.536
R4080 w_13193_29093.n1025 w_13193_29093.t215 135.919
R4081 w_13193_29093.t139 w_13193_29093.n1146 134.474
R4082 w_13193_29093.n251 w_13193_29093.n243 134.268
R4083 w_13193_29093.n246 w_13193_29093.n243 134.268
R4084 w_13193_29093.n2542 w_13193_29093.t140 133.483
R4085 w_13193_29093.n2548 w_13193_29093.t195 133.483
R4086 w_13193_29093.n2551 w_13193_29093.t129 133.483
R4087 w_13193_29093.n2551 w_13193_29093.t31 133.483
R4088 w_13193_29093.n2709 w_13193_29093.t92 132.058
R4089 w_13193_29093.n2761 w_13193_29093.t61 132.058
R4090 w_13193_29093.n2233 w_13193_29093.t46 130.713
R4091 w_13193_29093.n2700 w_13193_29093.t213 130.314
R4092 w_13193_29093.n1160 w_13193_29093.n1159 130.136
R4093 w_13193_29093.n734 w_13193_29093.n718 130.136
R4094 w_13193_29093.n1148 w_13193_29093.n1147 130.136
R4095 w_13193_29093.n874 w_13193_29093.n744 130.136
R4096 w_13193_29093.n875 w_13193_29093.n874 130.136
R4097 w_13193_29093.n876 w_13193_29093.n875 130.136
R4098 w_13193_29093.n876 w_13193_29093.n13 130.136
R4099 w_13193_29093.n887 w_13193_29093.n886 130.136
R4100 w_13193_29093.n889 w_13193_29093.n887 130.136
R4101 w_13193_29093.n889 w_13193_29093.n888 130.136
R4102 w_13193_29093.n888 w_13193_29093.n781 130.136
R4103 w_13193_29093.n1024 w_13193_29093.n1023 130.136
R4104 w_13193_29093.n999 w_13193_29093.n998 130.136
R4105 w_13193_29093.n1011 w_13193_29093.n1010 130.136
R4106 w_13193_29093.n2224 w_13193_29093.t157 130.001
R4107 w_13193_29093.n2226 w_13193_29093.t49 130.001
R4108 w_13193_29093.n2433 w_13193_29093.t225 130.001
R4109 w_13193_29093.n66 w_13193_29093.t303 130.001
R4110 w_13193_29093.n67 w_13193_29093.t232 130.001
R4111 w_13193_29093.n2266 w_13193_29093.t144 130.001
R4112 w_13193_29093.n2270 w_13193_29093.t175 130.001
R4113 w_13193_29093.n2273 w_13193_29093.t51 130.001
R4114 w_13193_29093.n2280 w_13193_29093.t155 130.001
R4115 w_13193_29093.n2252 w_13193_29093.t163 130.001
R4116 w_13193_29093.n2342 w_13193_29093.t239 130.001
R4117 w_13193_29093.n2258 w_13193_29093.t201 130.001
R4118 w_13193_29093.n2261 w_13193_29093.t207 130.001
R4119 w_13193_29093.n260 w_13193_29093.t258 129.47
R4120 w_13193_29093.t298 w_13193_29093.t87 128.906
R4121 w_13193_29093.t164 w_13193_29093.t17 128.906
R4122 w_13193_29093.t235 w_13193_29093.t71 128.906
R4123 w_13193_29093.t160 w_13193_29093.t158 128.906
R4124 w_13193_29093.n202 w_13193_29093.t32 128.562
R4125 w_13193_29093.n2544 w_13193_29093.t196 127.754
R4126 w_13193_29093.n2538 w_13193_29093.t151 127.754
R4127 w_13193_29093.n635 w_13193_29093.t170 125.797
R4128 w_13193_29093.n735 w_13193_29093.t286 125.797
R4129 w_13193_29093.t53 w_13193_29093.n15 125.797
R4130 w_13193_29093.t53 w_13193_29093.n24 124.352
R4131 w_13193_29093.t243 w_13193_29093.t6 122.996
R4132 w_13193_29093.n2447 w_13193_29093.t169 122.501
R4133 w_13193_29093.n2459 w_13193_29093.t147 122.501
R4134 w_13193_29093.n2462 w_13193_29093.t194 122.501
R4135 w_13193_29093.n2366 w_13193_29093.t192 122.501
R4136 w_13193_29093.n2371 w_13193_29093.t114 122.501
R4137 w_13193_29093.n2390 w_13193_29093.t294 122.501
R4138 w_13193_29093.n2534 w_13193_29093.t55 120.312
R4139 w_13193_29093.t210 w_13193_29093.n997 120.013
R4140 w_13193_29093.n981 w_13193_29093.t211 120.013
R4141 w_13193_29093.t231 w_13193_29093.t205 118.919
R4142 w_13193_29093.t176 w_13193_29093.t191 118.919
R4143 w_13193_29093.n2460 w_13193_29093.n2216 117.558
R4144 w_13193_29093.t300 w_13193_29093.n63 111.719
R4145 w_13193_29093.t166 w_13193_29093.t126 108.764
R4146 w_13193_29093.t152 w_13193_29093.t115 108.764
R4147 w_13193_29093.t134 w_13193_29093.t152 108.764
R4148 w_13193_29093.n2437 w_13193_29093.t7 107.028
R4149 w_13193_29093.t311 w_13193_29093.n2436 107.028
R4150 w_13193_29093.n2435 w_13193_29093.t148 107.028
R4151 w_13193_29093.t172 w_13193_29093.n2375 107.028
R4152 w_13193_29093.t228 w_13193_29093.n2221 106.796
R4153 w_13193_29093.n256 w_13193_29093.n255 101.718
R4154 w_13193_29093.n247 w_13193_29093.n244 101.718
R4155 w_13193_29093.n768 w_13193_29093.n767 101.718
R4156 w_13193_29093.n760 w_13193_29093.n759 101.718
R4157 w_13193_29093.t53 w_13193_29093.n16 100.799
R4158 w_13193_29093.t53 w_13193_29093.n25 100.799
R4159 w_13193_29093.n2721 w_13193_29093.t83 99.9042
R4160 w_13193_29093.n2701 w_13193_29093.t108 98.8769
R4161 w_13193_29093.n56 w_13193_29093.n55 97.8707
R4162 w_13193_29093.n52 w_13193_29093.n51 97.8707
R4163 w_13193_29093.n48 w_13193_29093.n47 97.8707
R4164 w_13193_29093.n44 w_13193_29093.n43 97.8707
R4165 w_13193_29093.n38 w_13193_29093.n37 97.8707
R4166 w_13193_29093.n1012 w_13193_29093.t23 96.8786
R4167 w_13193_29093.t238 w_13193_29093.t289 95.1356
R4168 w_13193_29093.t124 w_13193_29093.t39 95.1356
R4169 w_13193_29093.t33 w_13193_29093.t291 95.1356
R4170 w_13193_29093.t246 w_13193_29093.t48 95.1356
R4171 w_13193_29093.n219 w_13193_29093.n218 92.2603
R4172 w_13193_29093.n216 w_13193_29093.n215 92.2603
R4173 w_13193_29093.n2513 w_13193_29093.n2512 92.2603
R4174 w_13193_29093.n2521 w_13193_29093.n2520 92.2603
R4175 w_13193_29093.n2476 w_13193_29093.n237 92.2603
R4176 w_13193_29093.n2470 w_13193_29093.n240 92.2603
R4177 w_13193_29093.n1161 w_13193_29093.t212 91.0948
R4178 w_13193_29093.n765 w_13193_29093.n755 91.069
R4179 w_13193_29093.n758 w_13193_29093.n755 91.069
R4180 w_13193_29093.n762 w_13193_29093.n754 91.069
R4181 w_13193_29093.n763 w_13193_29093.n762 91.069
R4182 w_13193_29093.n252 w_13193_29093.n251 91.069
R4183 w_13193_29093.n251 w_13193_29093.n250 91.069
R4184 w_13193_29093.n246 w_13193_29093.n245 91.069
R4185 w_13193_29093.t53 w_13193_29093.n16 90.2509
R4186 w_13193_29093.t53 w_13193_29093.n25 90.2509
R4187 w_13193_29093.t133 w_13193_29093.t37 86.757
R4188 w_13193_29093.t149 w_13193_29093.t2 86.757
R4189 w_13193_29093.n201 w_13193_29093.t318 86.0829
R4190 w_13193_29093.n2382 w_13193_29093.n2377 84.306
R4191 w_13193_29093.n232 w_13193_29093.n231 84.306
R4192 w_13193_29093.n2501 w_13193_29093.n205 84.306
R4193 w_13193_29093.n2525 w_13193_29093.n207 84.306
R4194 w_13193_29093.n1080 w_13193_29093.n780 84.306
R4195 w_13193_29093.n746 w_13193_29093.n745 84.306
R4196 w_13193_29093.n2529 w_13193_29093.n208 84.306
R4197 w_13193_29093.n2502 w_13193_29093.n206 84.306
R4198 w_13193_29093.n226 w_13193_29093.n223 84.306
R4199 w_13193_29093.n2386 w_13193_29093.n2378 84.306
R4200 w_13193_29093.n201 w_13193_29093.t315 82.8829
R4201 w_13193_29093.n1161 w_13193_29093.t47 82.4192
R4202 w_13193_29093.t107 w_13193_29093.n21 82.4192
R4203 w_13193_29093.n736 w_13193_29093.t130 82.4192
R4204 w_13193_29093.n1079 w_13193_29093.n1077 82.4192
R4205 w_13193_29093.t269 w_13193_29093.t185 78.7125
R4206 w_13193_29093.t185 w_13193_29093.t111 78.7125
R4207 w_13193_29093.t83 w_13193_29093.t183 78.7125
R4208 w_13193_29093.t178 w_13193_29093.t242 77.6818
R4209 w_13193_29093.t131 w_13193_29093.t25 77.6818
R4210 w_13193_29093.t214 w_13193_29093.t27 77.6818
R4211 w_13193_29093.t27 w_13193_29093.t253 77.6818
R4212 w_13193_29093.t253 w_13193_29093.t243 77.6818
R4213 w_13193_29093.t6 w_13193_29093.t24 77.6818
R4214 w_13193_29093.t24 w_13193_29093.t296 77.6818
R4215 w_13193_29093.n1098 w_13193_29093.n1097 76.6354
R4216 w_13193_29093.t310 w_13193_29093.n987 76.6354
R4217 w_13193_29093.t202 w_13193_29093.n29 76.6354
R4218 w_13193_29093.n1012 w_13193_29093.t218 76.6354
R4219 w_13193_29093.n2187 w_13193_29093.n2186 76.3222
R4220 w_13193_29093.n2192 w_13193_29093.n2191 76.3222
R4221 w_13193_29093.n2195 w_13193_29093.n2194 76.3222
R4222 w_13193_29093.n1808 w_13193_29093.n268 76.3222
R4223 w_13193_29093.n1814 w_13193_29093.n1805 76.3222
R4224 w_13193_29093.n1834 w_13193_29093.n1833 76.3222
R4225 w_13193_29093.n1829 w_13193_29093.n397 76.3222
R4226 w_13193_29093.n1827 w_13193_29093.n1826 76.3222
R4227 w_13193_29093.n1822 w_13193_29093.n406 76.3222
R4228 w_13193_29093.n1820 w_13193_29093.n1819 76.3222
R4229 w_13193_29093.n1815 w_13193_29093.n1804 76.3222
R4230 w_13193_29093.n2068 w_13193_29093.n2067 76.3222
R4231 w_13193_29093.n2071 w_13193_29093.n2070 76.3222
R4232 w_13193_29093.n2077 w_13193_29093.n2076 76.3222
R4233 w_13193_29093.n2080 w_13193_29093.n2079 76.3222
R4234 w_13193_29093.n2087 w_13193_29093.n2085 76.3222
R4235 w_13193_29093.n2184 w_13193_29093.n272 76.3222
R4236 w_13193_29093.n1956 w_13193_29093.n303 76.3222
R4237 w_13193_29093.n1952 w_13193_29093.n302 76.3222
R4238 w_13193_29093.n1948 w_13193_29093.n301 76.3222
R4239 w_13193_29093.n1944 w_13193_29093.n300 76.3222
R4240 w_13193_29093.n299 w_13193_29093.n284 76.3222
R4241 w_13193_29093.n2154 w_13193_29093.n282 76.3222
R4242 w_13193_29093.n1960 w_13193_29093.n1959 76.3222
R4243 w_13193_29093.n2031 w_13193_29093.n2030 76.3222
R4244 w_13193_29093.n2034 w_13193_29093.n2033 76.3222
R4245 w_13193_29093.n2046 w_13193_29093.n2045 76.3222
R4246 w_13193_29093.n2049 w_13193_29093.n2048 76.3222
R4247 w_13193_29093.n2062 w_13193_29093.n2061 76.3222
R4248 w_13193_29093.n2104 w_13193_29093.n2103 76.3222
R4249 w_13193_29093.n2099 w_13193_29093.n2073 76.3222
R4250 w_13193_29093.n2097 w_13193_29093.n2096 76.3222
R4251 w_13193_29093.n2092 w_13193_29093.n2082 76.3222
R4252 w_13193_29093.n2090 w_13193_29093.n2089 76.3222
R4253 w_13193_29093.n2182 w_13193_29093.n275 76.3222
R4254 w_13193_29093.n2161 w_13193_29093.n2160 76.3222
R4255 w_13193_29093.n2162 w_13193_29093.n280 76.3222
R4256 w_13193_29093.n2169 w_13193_29093.n2168 76.3222
R4257 w_13193_29093.n2170 w_13193_29093.n278 76.3222
R4258 w_13193_29093.n2177 w_13193_29093.n2176 76.3222
R4259 w_13193_29093.n2181 w_13193_29093.n276 76.3222
R4260 w_13193_29093.n392 w_13193_29093.n391 76.3222
R4261 w_13193_29093.n395 w_13193_29093.n394 76.3222
R4262 w_13193_29093.n401 w_13193_29093.n400 76.3222
R4263 w_13193_29093.n404 w_13193_29093.n403 76.3222
R4264 w_13193_29093.n410 w_13193_29093.n409 76.3222
R4265 w_13193_29093.n413 w_13193_29093.n412 76.3222
R4266 w_13193_29093.n1709 w_13193_29093.n433 76.3222
R4267 w_13193_29093.n1705 w_13193_29093.n434 76.3222
R4268 w_13193_29093.n1701 w_13193_29093.n435 76.3222
R4269 w_13193_29093.n1697 w_13193_29093.n436 76.3222
R4270 w_13193_29093.n1778 w_13193_29093.n1777 76.3222
R4271 w_13193_29093.n1800 w_13193_29093.n1799 76.3222
R4272 w_13193_29093.n1797 w_13193_29093.n1796 76.3222
R4273 w_13193_29093.n1792 w_13193_29093.n418 76.3222
R4274 w_13193_29093.n1790 w_13193_29093.n1789 76.3222
R4275 w_13193_29093.n1785 w_13193_29093.n421 76.3222
R4276 w_13193_29093.n1783 w_13193_29093.n1782 76.3222
R4277 w_13193_29093.n1167 w_13193_29093.n286 76.3222
R4278 w_13193_29093.n1171 w_13193_29093.n287 76.3222
R4279 w_13193_29093.n1175 w_13193_29093.n288 76.3222
R4280 w_13193_29093.n1179 w_13193_29093.n289 76.3222
R4281 w_13193_29093.n1183 w_13193_29093.n290 76.3222
R4282 w_13193_29093.n1187 w_13193_29093.n291 76.3222
R4283 w_13193_29093.n1188 w_13193_29093.n630 76.3222
R4284 w_13193_29093.n1195 w_13193_29093.n1194 76.3222
R4285 w_13193_29093.n1196 w_13193_29093.n628 76.3222
R4286 w_13193_29093.n1203 w_13193_29093.n1202 76.3222
R4287 w_13193_29093.n1204 w_13193_29093.n626 76.3222
R4288 w_13193_29093.n1211 w_13193_29093.n1210 76.3222
R4289 w_13193_29093.n1140 w_13193_29093.n1105 76.3222
R4290 w_13193_29093.n1138 w_13193_29093.n1137 76.3222
R4291 w_13193_29093.n1133 w_13193_29093.n1114 76.3222
R4292 w_13193_29093.n1131 w_13193_29093.n1130 76.3222
R4293 w_13193_29093.n1126 w_13193_29093.n1124 76.3222
R4294 w_13193_29093.n1212 w_13193_29093.n625 76.3222
R4295 w_13193_29093.n1032 w_13193_29093.n1031 76.3222
R4296 w_13193_29093.n1035 w_13193_29093.n1034 76.3222
R4297 w_13193_29093.n1038 w_13193_29093.n1037 76.3222
R4298 w_13193_29093.n1044 w_13193_29093.n1043 76.3222
R4299 w_13193_29093.n1047 w_13193_29093.n1046 76.3222
R4300 w_13193_29093.n1048 w_13193_29093.n493 76.3222
R4301 w_13193_29093.n1771 w_13193_29093.n443 76.3222
R4302 w_13193_29093.n1767 w_13193_29093.n442 76.3222
R4303 w_13193_29093.n1763 w_13193_29093.n441 76.3222
R4304 w_13193_29093.n1759 w_13193_29093.n440 76.3222
R4305 w_13193_29093.n1755 w_13193_29093.n439 76.3222
R4306 w_13193_29093.n1751 w_13193_29093.n438 76.3222
R4307 w_13193_29093.n1503 w_13193_29093.n1502 76.3222
R4308 w_13193_29093.n1506 w_13193_29093.n1505 76.3222
R4309 w_13193_29093.n1509 w_13193_29093.n1508 76.3222
R4310 w_13193_29093.n1515 w_13193_29093.n1514 76.3222
R4311 w_13193_29093.n1518 w_13193_29093.n1517 76.3222
R4312 w_13193_29093.n1519 w_13193_29093.n490 76.3222
R4313 w_13193_29093.n1742 w_13193_29093.n425 76.3222
R4314 w_13193_29093.n1740 w_13193_29093.n426 76.3222
R4315 w_13193_29093.n1737 w_13193_29093.n427 76.3222
R4316 w_13193_29093.n1733 w_13193_29093.n428 76.3222
R4317 w_13193_29093.n1729 w_13193_29093.n429 76.3222
R4318 w_13193_29093.n1725 w_13193_29093.n430 76.3222
R4319 w_13193_29093.n1340 w_13193_29093.n1339 76.3222
R4320 w_13193_29093.n1343 w_13193_29093.n1342 76.3222
R4321 w_13193_29093.n1349 w_13193_29093.n1348 76.3222
R4322 w_13193_29093.n1352 w_13193_29093.n1351 76.3222
R4323 w_13193_29093.n1359 w_13193_29093.n1358 76.3222
R4324 w_13193_29093.n1360 w_13193_29093.n322 76.3222
R4325 w_13193_29093.n1541 w_13193_29093.n1540 76.3222
R4326 w_13193_29093.n1538 w_13193_29093.n1537 76.3222
R4327 w_13193_29093.n1533 w_13193_29093.n1511 76.3222
R4328 w_13193_29093.n1531 w_13193_29093.n1530 76.3222
R4329 w_13193_29093.n1526 w_13193_29093.n1522 76.3222
R4330 w_13193_29093.n1524 w_13193_29093.n1523 76.3222
R4331 w_13193_29093.n1103 w_13193_29093.n1102 76.3222
R4332 w_13193_29093.n1109 w_13193_29093.n1108 76.3222
R4333 w_13193_29093.n1112 w_13193_29093.n1111 76.3222
R4334 w_13193_29093.n1118 w_13193_29093.n1117 76.3222
R4335 w_13193_29093.n1123 w_13193_29093.n1120 76.3222
R4336 w_13193_29093.n1121 w_13193_29093.n622 76.3222
R4337 w_13193_29093.n1071 w_13193_29093.n1070 76.3222
R4338 w_13193_29093.n1068 w_13193_29093.n1067 76.3222
R4339 w_13193_29093.n1063 w_13193_29093.n1040 76.3222
R4340 w_13193_29093.n1061 w_13193_29093.n1060 76.3222
R4341 w_13193_29093.n1056 w_13193_29093.n1051 76.3222
R4342 w_13193_29093.n1054 w_13193_29093.n1053 76.3222
R4343 w_13193_29093.n1049 w_13193_29093.n1048 76.3222
R4344 w_13193_29093.n1046 w_13193_29093.n1045 76.3222
R4345 w_13193_29093.n1043 w_13193_29093.n1042 76.3222
R4346 w_13193_29093.n1037 w_13193_29093.n1036 76.3222
R4347 w_13193_29093.n1034 w_13193_29093.n1033 76.3222
R4348 w_13193_29093.n1031 w_13193_29093.n1027 76.3222
R4349 w_13193_29093.n1520 w_13193_29093.n1519 76.3222
R4350 w_13193_29093.n1517 w_13193_29093.n1516 76.3222
R4351 w_13193_29093.n1514 w_13193_29093.n1513 76.3222
R4352 w_13193_29093.n1508 w_13193_29093.n1507 76.3222
R4353 w_13193_29093.n1505 w_13193_29093.n1504 76.3222
R4354 w_13193_29093.n1502 w_13193_29093.n585 76.3222
R4355 w_13193_29093.n1055 w_13193_29093.n1054 76.3222
R4356 w_13193_29093.n1051 w_13193_29093.n1041 76.3222
R4357 w_13193_29093.n1062 w_13193_29093.n1061 76.3222
R4358 w_13193_29093.n1040 w_13193_29093.n1030 76.3222
R4359 w_13193_29093.n1069 w_13193_29093.n1068 76.3222
R4360 w_13193_29093.n1072 w_13193_29093.n1071 76.3222
R4361 w_13193_29093.n1525 w_13193_29093.n1524 76.3222
R4362 w_13193_29093.n1522 w_13193_29093.n1512 76.3222
R4363 w_13193_29093.n1532 w_13193_29093.n1531 76.3222
R4364 w_13193_29093.n1511 w_13193_29093.n1501 76.3222
R4365 w_13193_29093.n1539 w_13193_29093.n1538 76.3222
R4366 w_13193_29093.n1542 w_13193_29093.n1541 76.3222
R4367 w_13193_29093.n1122 w_13193_29093.n1121 76.3222
R4368 w_13193_29093.n1120 w_13193_29093.n1119 76.3222
R4369 w_13193_29093.n1117 w_13193_29093.n1116 76.3222
R4370 w_13193_29093.n1111 w_13193_29093.n1110 76.3222
R4371 w_13193_29093.n1108 w_13193_29093.n1107 76.3222
R4372 w_13193_29093.n1102 w_13193_29093.n1101 76.3222
R4373 w_13193_29093.n1125 w_13193_29093.n625 76.3222
R4374 w_13193_29093.n1124 w_13193_29093.n1115 76.3222
R4375 w_13193_29093.n1132 w_13193_29093.n1131 76.3222
R4376 w_13193_29093.n1114 w_13193_29093.n1106 76.3222
R4377 w_13193_29093.n1139 w_13193_29093.n1138 76.3222
R4378 w_13193_29093.n1105 w_13193_29093.n739 76.3222
R4379 w_13193_29093.n1784 w_13193_29093.n1783 76.3222
R4380 w_13193_29093.n421 w_13193_29093.n419 76.3222
R4381 w_13193_29093.n1791 w_13193_29093.n1790 76.3222
R4382 w_13193_29093.n418 w_13193_29093.n416 76.3222
R4383 w_13193_29093.n1798 w_13193_29093.n1797 76.3222
R4384 w_13193_29093.n1801 w_13193_29093.n1800 76.3222
R4385 w_13193_29093.n2178 w_13193_29093.n276 76.3222
R4386 w_13193_29093.n2176 w_13193_29093.n2175 76.3222
R4387 w_13193_29093.n2171 w_13193_29093.n2170 76.3222
R4388 w_13193_29093.n2168 w_13193_29093.n2167 76.3222
R4389 w_13193_29093.n2163 w_13193_29093.n2162 76.3222
R4390 w_13193_29093.n2160 w_13193_29093.n2159 76.3222
R4391 w_13193_29093.n1754 w_13193_29093.n438 76.3222
R4392 w_13193_29093.n1758 w_13193_29093.n439 76.3222
R4393 w_13193_29093.n1762 w_13193_29093.n440 76.3222
R4394 w_13193_29093.n1766 w_13193_29093.n441 76.3222
R4395 w_13193_29093.n1770 w_13193_29093.n442 76.3222
R4396 w_13193_29093.n1775 w_13193_29093.n1774 76.3222
R4397 w_13193_29093.n1722 w_13193_29093.n430 76.3222
R4398 w_13193_29093.n1726 w_13193_29093.n429 76.3222
R4399 w_13193_29093.n1730 w_13193_29093.n428 76.3222
R4400 w_13193_29093.n1734 w_13193_29093.n427 76.3222
R4401 w_13193_29093.n1738 w_13193_29093.n426 76.3222
R4402 w_13193_29093.n454 w_13193_29093.n425 76.3222
R4403 w_13193_29093.n1777 w_13193_29093.n422 76.3222
R4404 w_13193_29093.n436 w_13193_29093.n424 76.3222
R4405 w_13193_29093.n1698 w_13193_29093.n435 76.3222
R4406 w_13193_29093.n1702 w_13193_29093.n434 76.3222
R4407 w_13193_29093.n1706 w_13193_29093.n433 76.3222
R4408 w_13193_29093.n1710 w_13193_29093.n432 76.3222
R4409 w_13193_29093.n1210 w_13193_29093.n1209 76.3222
R4410 w_13193_29093.n1205 w_13193_29093.n1204 76.3222
R4411 w_13193_29093.n1202 w_13193_29093.n1201 76.3222
R4412 w_13193_29093.n1197 w_13193_29093.n1196 76.3222
R4413 w_13193_29093.n1194 w_13193_29093.n1193 76.3222
R4414 w_13193_29093.n1189 w_13193_29093.n1188 76.3222
R4415 w_13193_29093.n1959 w_13193_29093.n1938 76.3222
R4416 w_13193_29093.n2032 w_13193_29093.n2031 76.3222
R4417 w_13193_29093.n2033 w_13193_29093.n1933 76.3222
R4418 w_13193_29093.n2047 w_13193_29093.n2046 76.3222
R4419 w_13193_29093.n2048 w_13193_29093.n1925 76.3222
R4420 w_13193_29093.n2063 w_13193_29093.n2062 76.3222
R4421 w_13193_29093.n1184 w_13193_29093.n291 76.3222
R4422 w_13193_29093.n1180 w_13193_29093.n290 76.3222
R4423 w_13193_29093.n1176 w_13193_29093.n289 76.3222
R4424 w_13193_29093.n1172 w_13193_29093.n288 76.3222
R4425 w_13193_29093.n1168 w_13193_29093.n287 76.3222
R4426 w_13193_29093.n631 w_13193_29093.n285 76.3222
R4427 w_13193_29093.n2155 w_13193_29093.n2154 76.3222
R4428 w_13193_29093.n1943 w_13193_29093.n299 76.3222
R4429 w_13193_29093.n1947 w_13193_29093.n300 76.3222
R4430 w_13193_29093.n1951 w_13193_29093.n301 76.3222
R4431 w_13193_29093.n1955 w_13193_29093.n302 76.3222
R4432 w_13193_29093.n1941 w_13193_29093.n304 76.3222
R4433 w_13193_29093.n2128 w_13193_29093.n2127 76.3222
R4434 w_13193_29093.n2125 w_13193_29093.n2124 76.3222
R4435 w_13193_29093.n2120 w_13193_29093.n311 76.3222
R4436 w_13193_29093.n2118 w_13193_29093.n2117 76.3222
R4437 w_13193_29093.n2113 w_13193_29093.n314 76.3222
R4438 w_13193_29093.n2111 w_13193_29093.n2110 76.3222
R4439 w_13193_29093.n1379 w_13193_29093.n1378 76.3222
R4440 w_13193_29093.n1374 w_13193_29093.n1345 76.3222
R4441 w_13193_29093.n1372 w_13193_29093.n1371 76.3222
R4442 w_13193_29093.n1367 w_13193_29093.n1354 76.3222
R4443 w_13193_29093.n1365 w_13193_29093.n1364 76.3222
R4444 w_13193_29093.n1355 w_13193_29093.n315 76.3222
R4445 w_13193_29093.n1232 w_13193_29093.n1231 76.3222
R4446 w_13193_29093.n1303 w_13193_29093.n1302 76.3222
R4447 w_13193_29093.n1306 w_13193_29093.n1305 76.3222
R4448 w_13193_29093.n1318 w_13193_29093.n1317 76.3222
R4449 w_13193_29093.n1321 w_13193_29093.n1320 76.3222
R4450 w_13193_29093.n1334 w_13193_29093.n1333 76.3222
R4451 w_13193_29093.n2152 w_13193_29093.n305 76.3222
R4452 w_13193_29093.n2151 w_13193_29093.n293 76.3222
R4453 w_13193_29093.n2147 w_13193_29093.n294 76.3222
R4454 w_13193_29093.n2143 w_13193_29093.n295 76.3222
R4455 w_13193_29093.n2139 w_13193_29093.n296 76.3222
R4456 w_13193_29093.n2135 w_13193_29093.n297 76.3222
R4457 w_13193_29093.n305 w_13193_29093.n292 76.3222
R4458 w_13193_29093.n1231 w_13193_29093.n1228 76.3222
R4459 w_13193_29093.n1304 w_13193_29093.n1303 76.3222
R4460 w_13193_29093.n1305 w_13193_29093.n1223 76.3222
R4461 w_13193_29093.n1319 w_13193_29093.n1318 76.3222
R4462 w_13193_29093.n1320 w_13193_29093.n1215 76.3222
R4463 w_13193_29093.n1335 w_13193_29093.n1334 76.3222
R4464 w_13193_29093.n2132 w_13193_29093.n297 76.3222
R4465 w_13193_29093.n2136 w_13193_29093.n296 76.3222
R4466 w_13193_29093.n2140 w_13193_29093.n295 76.3222
R4467 w_13193_29093.n2144 w_13193_29093.n294 76.3222
R4468 w_13193_29093.n2148 w_13193_29093.n293 76.3222
R4469 w_13193_29093.n2112 w_13193_29093.n2111 76.3222
R4470 w_13193_29093.n314 w_13193_29093.n312 76.3222
R4471 w_13193_29093.n2119 w_13193_29093.n2118 76.3222
R4472 w_13193_29093.n311 w_13193_29093.n309 76.3222
R4473 w_13193_29093.n2126 w_13193_29093.n2125 76.3222
R4474 w_13193_29093.n2129 w_13193_29093.n2128 76.3222
R4475 w_13193_29093.n1361 w_13193_29093.n1360 76.3222
R4476 w_13193_29093.n1358 w_13193_29093.n1357 76.3222
R4477 w_13193_29093.n1351 w_13193_29093.n1350 76.3222
R4478 w_13193_29093.n1348 w_13193_29093.n1347 76.3222
R4479 w_13193_29093.n1342 w_13193_29093.n1341 76.3222
R4480 w_13193_29093.n1339 w_13193_29093.n1338 76.3222
R4481 w_13193_29093.n1356 w_13193_29093.n1355 76.3222
R4482 w_13193_29093.n1366 w_13193_29093.n1365 76.3222
R4483 w_13193_29093.n1354 w_13193_29093.n1346 76.3222
R4484 w_13193_29093.n1373 w_13193_29093.n1372 76.3222
R4485 w_13193_29093.n1345 w_13193_29093.n1337 76.3222
R4486 w_13193_29093.n1380 w_13193_29093.n1379 76.3222
R4487 w_13193_29093.n2086 w_13193_29093.n272 76.3222
R4488 w_13193_29093.n2085 w_13193_29093.n2084 76.3222
R4489 w_13193_29093.n2079 w_13193_29093.n2078 76.3222
R4490 w_13193_29093.n2076 w_13193_29093.n2075 76.3222
R4491 w_13193_29093.n2070 w_13193_29093.n2069 76.3222
R4492 w_13193_29093.n2067 w_13193_29093.n2066 76.3222
R4493 w_13193_29093.n2083 w_13193_29093.n275 76.3222
R4494 w_13193_29093.n2091 w_13193_29093.n2090 76.3222
R4495 w_13193_29093.n2082 w_13193_29093.n2074 76.3222
R4496 w_13193_29093.n2098 w_13193_29093.n2097 76.3222
R4497 w_13193_29093.n2073 w_13193_29093.n2065 76.3222
R4498 w_13193_29093.n2105 w_13193_29093.n2104 76.3222
R4499 w_13193_29093.n1695 w_13193_29093.n437 76.3222
R4500 w_13193_29093.n412 w_13193_29093.n411 76.3222
R4501 w_13193_29093.n409 w_13193_29093.n408 76.3222
R4502 w_13193_29093.n403 w_13193_29093.n402 76.3222
R4503 w_13193_29093.n400 w_13193_29093.n399 76.3222
R4504 w_13193_29093.n394 w_13193_29093.n393 76.3222
R4505 w_13193_29093.n391 w_13193_29093.n390 76.3222
R4506 w_13193_29093.n1804 w_13193_29093.n407 76.3222
R4507 w_13193_29093.n1821 w_13193_29093.n1820 76.3222
R4508 w_13193_29093.n406 w_13193_29093.n398 76.3222
R4509 w_13193_29093.n1828 w_13193_29093.n1827 76.3222
R4510 w_13193_29093.n397 w_13193_29093.n389 76.3222
R4511 w_13193_29093.n1835 w_13193_29093.n1834 76.3222
R4512 w_13193_29093.n1811 w_13193_29093.n1805 76.3222
R4513 w_13193_29093.n1809 w_13193_29093.n1808 76.3222
R4514 w_13193_29093.n2196 w_13193_29093.n2195 76.3222
R4515 w_13193_29093.n2193 w_13193_29093.n2192 76.3222
R4516 w_13193_29093.n2186 w_13193_29093.n270 76.3222
R4517 w_13193_29093.n1632 w_13193_29093.n1593 74.5978
R4518 w_13193_29093.n1633 w_13193_29093.n1632 74.5978
R4519 w_13193_29093.n1879 w_13193_29093.n338 74.5978
R4520 w_13193_29093.n1880 w_13193_29093.n1879 74.5978
R4521 w_13193_29093.n2005 w_13193_29093.n1966 74.5978
R4522 w_13193_29093.n2006 w_13193_29093.n2005 74.5978
R4523 w_13193_29093.n562 w_13193_29093.n519 74.5978
R4524 w_13193_29093.n563 w_13193_29093.n562 74.5978
R4525 w_13193_29093.n942 w_13193_29093.n916 74.5978
R4526 w_13193_29093.n945 w_13193_29093.n916 74.5978
R4527 w_13193_29093.n1439 w_13193_29093.n1394 74.5978
R4528 w_13193_29093.n1440 w_13193_29093.n1439 74.5978
R4529 w_13193_29093.n849 w_13193_29093.n796 74.5978
R4530 w_13193_29093.n846 w_13193_29093.n796 74.5978
R4531 w_13193_29093.n679 w_13193_29093.n649 74.5978
R4532 w_13193_29093.n682 w_13193_29093.n649 74.5978
R4533 w_13193_29093.n1277 w_13193_29093.n1238 74.5978
R4534 w_13193_29093.n1278 w_13193_29093.n1277 74.5978
R4535 w_13193_29093.t237 w_13193_29093.t293 71.3518
R4536 w_13193_29093.n2714 w_13193_29093.n41 70.4005
R4537 w_13193_29093.n2706 w_13193_29093.n41 70.4005
R4538 w_13193_29093.n1692 w_13193_29093.n1691 69.3109
R4539 w_13193_29093.n1693 w_13193_29093.n1692 69.3109
R4540 w_13193_29093.n1847 w_13193_29093.n1846 69.3109
R4541 w_13193_29093.n1848 w_13193_29093.n1847 69.3109
R4542 w_13193_29093.n2056 w_13193_29093.n2055 69.3109
R4543 w_13193_29093.n2057 w_13193_29093.n2056 69.3109
R4544 w_13193_29093.n530 w_13193_29093.n509 69.3109
R4545 w_13193_29093.n531 w_13193_29093.n530 69.3109
R4546 w_13193_29093.n1017 w_13193_29093.n1016 69.3109
R4547 w_13193_29093.n1017 w_13193_29093.n924 69.3109
R4548 w_13193_29093.n1407 w_13193_29093.n599 69.3109
R4549 w_13193_29093.n1408 w_13193_29093.n1407 69.3109
R4550 w_13193_29093.n896 w_13193_29093.n895 69.3109
R4551 w_13193_29093.n895 w_13193_29093.n787 69.3109
R4552 w_13193_29093.n1153 w_13193_29093.n1152 69.3109
R4553 w_13193_29093.n1153 w_13193_29093.n657 69.3109
R4554 w_13193_29093.n1328 w_13193_29093.n1327 69.3109
R4555 w_13193_29093.n1329 w_13193_29093.n1328 69.3109
R4556 w_13193_29093.n2203 w_13193_29093.n2200 69.0321
R4557 w_13193_29093.t0 w_13193_29093.n159 68.7505
R4558 w_13193_29093.t220 w_13193_29093.n2533 68.7505
R4559 w_13193_29093.t79 w_13193_29093.n2531 68.7505
R4560 w_13193_29093.t53 w_13193_29093.n29 67.9598
R4561 w_13193_29093.n2712 w_13193_29093.t13 67.5444
R4562 w_13193_29093.n2763 w_13193_29093.t13 67.5444
R4563 w_13193_29093.n2354 w_13193_29093.n2226 66.69
R4564 w_13193_29093.n2433 w_13193_29093.n2432 66.69
R4565 w_13193_29093.n2426 w_13193_29093.n66 66.69
R4566 w_13193_29093.n2420 w_13193_29093.n67 66.69
R4567 w_13193_29093.n2329 w_13193_29093.n2224 66.69
R4568 w_13193_29093.n2303 w_13193_29093.n2266 66.69
R4569 w_13193_29093.n2298 w_13193_29093.n2270 66.69
R4570 w_13193_29093.n2291 w_13193_29093.n2273 66.69
R4571 w_13193_29093.n2285 w_13193_29093.n2280 66.69
R4572 w_13193_29093.n2253 w_13193_29093.n2252 66.69
R4573 w_13193_29093.n2725 w_13193_29093.n2719 66.5605
R4574 w_13193_29093.n2725 w_13193_29093.n2724 66.5605
R4575 w_13193_29093.n2726 w_13193_29093.n2725 65.9634
R4576 w_13193_29093.n2448 w_13193_29093.n2447 65.9579
R4577 w_13193_29093.n2459 w_13193_29093.n2458 65.9579
R4578 w_13193_29093.n2463 w_13193_29093.n2462 65.9579
R4579 w_13193_29093.n1616 w_13193_29093.t59 65.8183
R4580 w_13193_29093.n1610 w_13193_29093.t59 65.8183
R4581 w_13193_29093.n1608 w_13193_29093.t59 65.8183
R4582 w_13193_29093.n1603 w_13193_29093.t59 65.8183
R4583 w_13193_29093.n1600 w_13193_29093.t59 65.8183
R4584 w_13193_29093.n1623 w_13193_29093.t59 65.8183
R4585 w_13193_29093.n1597 w_13193_29093.t59 65.8183
R4586 w_13193_29093.n1630 w_13193_29093.t59 65.8183
R4587 w_13193_29093.n1638 w_13193_29093.t59 65.8183
R4588 w_13193_29093.n1640 w_13193_29093.t59 65.8183
R4589 w_13193_29093.n1646 w_13193_29093.t59 65.8183
R4590 w_13193_29093.n1648 w_13193_29093.t59 65.8183
R4591 w_13193_29093.n1863 w_13193_29093.t76 65.8183
R4592 w_13193_29093.n1857 w_13193_29093.t76 65.8183
R4593 w_13193_29093.n1855 w_13193_29093.t76 65.8183
R4594 w_13193_29093.n1849 w_13193_29093.t76 65.8183
R4595 w_13193_29093.n345 w_13193_29093.t76 65.8183
R4596 w_13193_29093.n1870 w_13193_29093.t76 65.8183
R4597 w_13193_29093.n342 w_13193_29093.t76 65.8183
R4598 w_13193_29093.n1877 w_13193_29093.t76 65.8183
R4599 w_13193_29093.n1885 w_13193_29093.t76 65.8183
R4600 w_13193_29093.n1887 w_13193_29093.t76 65.8183
R4601 w_13193_29093.n1893 w_13193_29093.t76 65.8183
R4602 w_13193_29093.n334 w_13193_29093.t76 65.8183
R4603 w_13193_29093.n1989 w_13193_29093.t75 65.8183
R4604 w_13193_29093.n1983 w_13193_29093.t75 65.8183
R4605 w_13193_29093.n1981 w_13193_29093.t75 65.8183
R4606 w_13193_29093.n1976 w_13193_29093.t75 65.8183
R4607 w_13193_29093.n1973 w_13193_29093.t75 65.8183
R4608 w_13193_29093.n1996 w_13193_29093.t75 65.8183
R4609 w_13193_29093.n1970 w_13193_29093.t75 65.8183
R4610 w_13193_29093.n2003 w_13193_29093.t75 65.8183
R4611 w_13193_29093.n2011 w_13193_29093.t75 65.8183
R4612 w_13193_29093.n2013 w_13193_29093.t75 65.8183
R4613 w_13193_29093.n2019 w_13193_29093.t75 65.8183
R4614 w_13193_29093.n1940 w_13193_29093.t75 65.8183
R4615 w_13193_29093.n2025 w_13193_29093.t75 65.8183
R4616 w_13193_29093.n2038 w_13193_29093.t75 65.8183
R4617 w_13193_29093.n2040 w_13193_29093.t75 65.8183
R4618 w_13193_29093.n2053 w_13193_29093.t75 65.8183
R4619 w_13193_29093.n546 w_13193_29093.t77 65.8183
R4620 w_13193_29093.n540 w_13193_29093.t77 65.8183
R4621 w_13193_29093.n538 w_13193_29093.t77 65.8183
R4622 w_13193_29093.n532 w_13193_29093.t77 65.8183
R4623 w_13193_29093.n526 w_13193_29093.t77 65.8183
R4624 w_13193_29093.n553 w_13193_29093.t77 65.8183
R4625 w_13193_29093.n523 w_13193_29093.t77 65.8183
R4626 w_13193_29093.n560 w_13193_29093.t77 65.8183
R4627 w_13193_29093.n568 w_13193_29093.t77 65.8183
R4628 w_13193_29093.n570 w_13193_29093.t77 65.8183
R4629 w_13193_29093.n576 w_13193_29093.t77 65.8183
R4630 w_13193_29093.n578 w_13193_29093.t77 65.8183
R4631 w_13193_29093.t99 w_13193_29093.n915 65.8183
R4632 w_13193_29093.t99 w_13193_29093.n913 65.8183
R4633 w_13193_29093.t99 w_13193_29093.n911 65.8183
R4634 w_13193_29093.t99 w_13193_29093.n909 65.8183
R4635 w_13193_29093.t99 w_13193_29093.n917 65.8183
R4636 w_13193_29093.t99 w_13193_29093.n918 65.8183
R4637 w_13193_29093.t99 w_13193_29093.n919 65.8183
R4638 w_13193_29093.t99 w_13193_29093.n920 65.8183
R4639 w_13193_29093.t99 w_13193_29093.n914 65.8183
R4640 w_13193_29093.t99 w_13193_29093.n912 65.8183
R4641 w_13193_29093.t99 w_13193_29093.n910 65.8183
R4642 w_13193_29093.t99 w_13193_29093.n908 65.8183
R4643 w_13193_29093.n1018 w_13193_29093.t99 65.8183
R4644 w_13193_29093.t99 w_13193_29093.n921 65.8183
R4645 w_13193_29093.t99 w_13193_29093.n922 65.8183
R4646 w_13193_29093.t99 w_13193_29093.n923 65.8183
R4647 w_13193_29093.n1423 w_13193_29093.t104 65.8183
R4648 w_13193_29093.n1417 w_13193_29093.t104 65.8183
R4649 w_13193_29093.n1415 w_13193_29093.t104 65.8183
R4650 w_13193_29093.n1409 w_13193_29093.t104 65.8183
R4651 w_13193_29093.n1401 w_13193_29093.t104 65.8183
R4652 w_13193_29093.n1430 w_13193_29093.t104 65.8183
R4653 w_13193_29093.n1398 w_13193_29093.t104 65.8183
R4654 w_13193_29093.n1437 w_13193_29093.t104 65.8183
R4655 w_13193_29093.n1445 w_13193_29093.t104 65.8183
R4656 w_13193_29093.n1447 w_13193_29093.t104 65.8183
R4657 w_13193_29093.n1453 w_13193_29093.t104 65.8183
R4658 w_13193_29093.n619 w_13193_29093.t104 65.8183
R4659 w_13193_29093.n1460 w_13193_29093.t104 65.8183
R4660 w_13193_29093.n616 w_13193_29093.t104 65.8183
R4661 w_13193_29093.n1481 w_13193_29093.t104 65.8183
R4662 w_13193_29093.n1484 w_13193_29093.t104 65.8183
R4663 w_13193_29093.t58 w_13193_29093.n795 65.8183
R4664 w_13193_29093.t58 w_13193_29093.n793 65.8183
R4665 w_13193_29093.t58 w_13193_29093.n791 65.8183
R4666 w_13193_29093.t58 w_13193_29093.n789 65.8183
R4667 w_13193_29093.t58 w_13193_29093.n797 65.8183
R4668 w_13193_29093.t58 w_13193_29093.n798 65.8183
R4669 w_13193_29093.t58 w_13193_29093.n799 65.8183
R4670 w_13193_29093.t58 w_13193_29093.n800 65.8183
R4671 w_13193_29093.t58 w_13193_29093.n794 65.8183
R4672 w_13193_29093.t58 w_13193_29093.n792 65.8183
R4673 w_13193_29093.t58 w_13193_29093.n790 65.8183
R4674 w_13193_29093.t58 w_13193_29093.n788 65.8183
R4675 w_13193_29093.t74 w_13193_29093.n648 65.8183
R4676 w_13193_29093.t74 w_13193_29093.n646 65.8183
R4677 w_13193_29093.t74 w_13193_29093.n644 65.8183
R4678 w_13193_29093.t74 w_13193_29093.n642 65.8183
R4679 w_13193_29093.t74 w_13193_29093.n650 65.8183
R4680 w_13193_29093.t74 w_13193_29093.n651 65.8183
R4681 w_13193_29093.t74 w_13193_29093.n652 65.8183
R4682 w_13193_29093.t74 w_13193_29093.n653 65.8183
R4683 w_13193_29093.t74 w_13193_29093.n647 65.8183
R4684 w_13193_29093.t74 w_13193_29093.n645 65.8183
R4685 w_13193_29093.t74 w_13193_29093.n643 65.8183
R4686 w_13193_29093.t74 w_13193_29093.n641 65.8183
R4687 w_13193_29093.t74 w_13193_29093.n654 65.8183
R4688 w_13193_29093.n1154 w_13193_29093.t74 65.8183
R4689 w_13193_29093.t74 w_13193_29093.n655 65.8183
R4690 w_13193_29093.t74 w_13193_29093.n656 65.8183
R4691 w_13193_29093.t58 w_13193_29093.n801 65.8183
R4692 w_13193_29093.t58 w_13193_29093.n802 65.8183
R4693 w_13193_29093.t58 w_13193_29093.n803 65.8183
R4694 w_13193_29093.t58 w_13193_29093.n894 65.8183
R4695 w_13193_29093.n1552 w_13193_29093.t77 65.8183
R4696 w_13193_29093.n1554 w_13193_29093.t77 65.8183
R4697 w_13193_29093.n1565 w_13193_29093.t77 65.8183
R4698 w_13193_29093.n1568 w_13193_29093.t77 65.8183
R4699 w_13193_29093.n1261 w_13193_29093.t52 65.8183
R4700 w_13193_29093.n1255 w_13193_29093.t52 65.8183
R4701 w_13193_29093.n1253 w_13193_29093.t52 65.8183
R4702 w_13193_29093.n1248 w_13193_29093.t52 65.8183
R4703 w_13193_29093.n1245 w_13193_29093.t52 65.8183
R4704 w_13193_29093.n1268 w_13193_29093.t52 65.8183
R4705 w_13193_29093.n1242 w_13193_29093.t52 65.8183
R4706 w_13193_29093.n1275 w_13193_29093.t52 65.8183
R4707 w_13193_29093.n1283 w_13193_29093.t52 65.8183
R4708 w_13193_29093.n1285 w_13193_29093.t52 65.8183
R4709 w_13193_29093.n1291 w_13193_29093.t52 65.8183
R4710 w_13193_29093.n1230 w_13193_29093.t52 65.8183
R4711 w_13193_29093.n1297 w_13193_29093.t52 65.8183
R4712 w_13193_29093.n1310 w_13193_29093.t52 65.8183
R4713 w_13193_29093.n1312 w_13193_29093.t52 65.8183
R4714 w_13193_29093.n1325 w_13193_29093.t52 65.8183
R4715 w_13193_29093.n1904 w_13193_29093.t76 65.8183
R4716 w_13193_29093.n1907 w_13193_29093.t76 65.8183
R4717 w_13193_29093.n371 w_13193_29093.t76 65.8183
R4718 w_13193_29093.n373 w_13193_29093.t76 65.8183
R4719 w_13193_29093.n1667 w_13193_29093.t59 65.8183
R4720 w_13193_29093.n1670 w_13193_29093.t59 65.8183
R4721 w_13193_29093.n478 w_13193_29093.t59 65.8183
R4722 w_13193_29093.n1689 w_13193_29093.t59 65.8183
R4723 w_13193_29093.n2414 w_13193_29093.n2366 65.3889
R4724 w_13193_29093.n2402 w_13193_29093.n2371 65.3889
R4725 w_13193_29093.n2391 w_13193_29093.n2390 65.3889
R4726 w_13193_29093.t53 w_13193_29093.n21 62.176
R4727 w_13193_29093.t53 w_13193_29093.n13 62.176
R4728 w_13193_29093.n2692 w_13193_29093.n2691 60.8005
R4729 w_13193_29093.n2664 w_13193_29093.n147 60.8005
R4730 w_13193_29093.n2343 w_13193_29093.n2342 60.8005
R4731 w_13193_29093.n2234 w_13193_29093.n2233 60.8005
R4732 w_13193_29093.n2316 w_13193_29093.n2258 60.8005
R4733 w_13193_29093.n2262 w_13193_29093.n2261 60.8005
R4734 w_13193_29093.t87 w_13193_29093.t284 60.1567
R4735 w_13193_29093.t55 w_13193_29093.t271 60.1567
R4736 w_13193_29093.t17 w_13193_29093.t122 60.1567
R4737 w_13193_29093.t35 w_13193_29093.t145 60.1567
R4738 w_13193_29093.t158 w_13193_29093.t120 60.1567
R4739 w_13193_29093.t103 w_13193_29093.n221 60.0005
R4740 w_13193_29093.n224 w_13193_29093.t103 60.0005
R4741 w_13193_29093.t69 w_13193_29093.n2496 60.0005
R4742 w_13193_29093.n2500 w_13193_29093.t69 60.0005
R4743 w_13193_29093.n40 w_13193_29093.t38 60.0005
R4744 w_13193_29093.n40 w_13193_29093.t110 60.0005
R4745 w_13193_29093.n2705 w_13193_29093.t241 60.0005
R4746 w_13193_29093.n2705 w_13193_29093.t94 60.0005
R4747 w_13193_29093.n2713 w_13193_29093.t65 60.0005
R4748 w_13193_29093.n2713 w_13193_29093.t252 60.0005
R4749 w_13193_29093.n58 w_13193_29093.t186 60.0005
R4750 w_13193_29093.n58 w_13193_29093.t112 60.0005
R4751 w_13193_29093.n59 w_13193_29093.t98 60.0005
R4752 w_13193_29093.n59 w_13193_29093.t270 60.0005
R4753 w_13193_29093.n2720 w_13193_29093.t184 60.0005
R4754 w_13193_29093.n2720 w_13193_29093.t84 60.0005
R4755 w_13193_29093.n2694 w_13193_29093.t197 59.46
R4756 w_13193_29093.n2389 w_13193_29093.t248 59.46
R4757 w_13193_29093.n886 w_13193_29093.t278 59.2841
R4758 w_13193_29093.n2056 w_13193_29093.t75 57.8461
R4759 w_13193_29093.t99 w_13193_29093.n1017 57.8461
R4760 w_13193_29093.n1407 w_13193_29093.t104 57.8461
R4761 w_13193_29093.t74 w_13193_29093.n1153 57.8461
R4762 w_13193_29093.n895 w_13193_29093.t58 57.8461
R4763 w_13193_29093.n530 w_13193_29093.t77 57.8461
R4764 w_13193_29093.n1328 w_13193_29093.t52 57.8461
R4765 w_13193_29093.n1847 w_13193_29093.t76 57.8461
R4766 w_13193_29093.n1692 w_13193_29093.t59 57.8461
R4767 w_13193_29093.t53 w_13193_29093.t263 57.8382
R4768 w_13193_29093.t53 w_13193_29093.t265 57.8382
R4769 w_13193_29093.t53 w_13193_29093.t111 57.5208
R4770 w_13193_29093.n1632 w_13193_29093.t59 55.2026
R4771 w_13193_29093.n1879 w_13193_29093.t76 55.2026
R4772 w_13193_29093.n2005 w_13193_29093.t75 55.2026
R4773 w_13193_29093.n562 w_13193_29093.t77 55.2026
R4774 w_13193_29093.t99 w_13193_29093.n916 55.2026
R4775 w_13193_29093.n1439 w_13193_29093.t104 55.2026
R4776 w_13193_29093.t58 w_13193_29093.n796 55.2026
R4777 w_13193_29093.t74 w_13193_29093.n649 55.2026
R4778 w_13193_29093.n1277 w_13193_29093.t52 55.2026
R4779 w_13193_29093.n2721 w_13193_29093.n30 54.4934
R4780 w_13193_29093.n2750 w_13193_29093.n41 54.4005
R4781 w_13193_29093.n1097 w_13193_29093.n744 53.5003
R4782 w_13193_29093.n997 w_13193_29093.t310 53.5003
R4783 w_13193_29093.n981 w_13193_29093.t202 53.5003
R4784 w_13193_29093.t218 w_13193_29093.n28 53.5003
R4785 w_13193_29093.n1667 w_13193_29093.n1666 53.3664
R4786 w_13193_29093.n1670 w_13193_29093.n1669 53.3664
R4787 w_13193_29093.n483 w_13193_29093.n478 53.3664
R4788 w_13193_29093.n1689 w_13193_29093.n1688 53.3664
R4789 w_13193_29093.n1648 w_13193_29093.n486 53.3664
R4790 w_13193_29093.n1647 w_13193_29093.n1646 53.3664
R4791 w_13193_29093.n1640 w_13193_29093.n1591 53.3664
R4792 w_13193_29093.n1639 w_13193_29093.n1638 53.3664
R4793 w_13193_29093.n1630 w_13193_29093.n1629 53.3664
R4794 w_13193_29093.n1625 w_13193_29093.n1597 53.3664
R4795 w_13193_29093.n1623 w_13193_29093.n1622 53.3664
R4796 w_13193_29093.n1618 w_13193_29093.n1600 53.3664
R4797 w_13193_29093.n1603 w_13193_29093.n462 53.3664
R4798 w_13193_29093.n1608 w_13193_29093.n1607 53.3664
R4799 w_13193_29093.n1611 w_13193_29093.n1610 53.3664
R4800 w_13193_29093.n1616 w_13193_29093.n1615 53.3664
R4801 w_13193_29093.n1617 w_13193_29093.n1616 53.3664
R4802 w_13193_29093.n1610 w_13193_29093.n1601 53.3664
R4803 w_13193_29093.n1609 w_13193_29093.n1608 53.3664
R4804 w_13193_29093.n1604 w_13193_29093.n1603 53.3664
R4805 w_13193_29093.n1600 w_13193_29093.n1598 53.3664
R4806 w_13193_29093.n1624 w_13193_29093.n1623 53.3664
R4807 w_13193_29093.n1597 w_13193_29093.n1595 53.3664
R4808 w_13193_29093.n1631 w_13193_29093.n1630 53.3664
R4809 w_13193_29093.n1638 w_13193_29093.n1637 53.3664
R4810 w_13193_29093.n1641 w_13193_29093.n1640 53.3664
R4811 w_13193_29093.n1646 w_13193_29093.n1645 53.3664
R4812 w_13193_29093.n1649 w_13193_29093.n1648 53.3664
R4813 w_13193_29093.n1904 w_13193_29093.n1903 53.3664
R4814 w_13193_29093.n1907 w_13193_29093.n1906 53.3664
R4815 w_13193_29093.n371 w_13193_29093.n331 53.3664
R4816 w_13193_29093.n374 w_13193_29093.n373 53.3664
R4817 w_13193_29093.n1898 w_13193_29093.n334 53.3664
R4818 w_13193_29093.n1894 w_13193_29093.n1893 53.3664
R4819 w_13193_29093.n1887 w_13193_29093.n336 53.3664
R4820 w_13193_29093.n1886 w_13193_29093.n1885 53.3664
R4821 w_13193_29093.n1877 w_13193_29093.n1876 53.3664
R4822 w_13193_29093.n1872 w_13193_29093.n342 53.3664
R4823 w_13193_29093.n1870 w_13193_29093.n1869 53.3664
R4824 w_13193_29093.n1865 w_13193_29093.n345 53.3664
R4825 w_13193_29093.n1850 w_13193_29093.n1849 53.3664
R4826 w_13193_29093.n1855 w_13193_29093.n1854 53.3664
R4827 w_13193_29093.n1858 w_13193_29093.n1857 53.3664
R4828 w_13193_29093.n1863 w_13193_29093.n1862 53.3664
R4829 w_13193_29093.n1864 w_13193_29093.n1863 53.3664
R4830 w_13193_29093.n1857 w_13193_29093.n346 53.3664
R4831 w_13193_29093.n1856 w_13193_29093.n1855 53.3664
R4832 w_13193_29093.n1849 w_13193_29093.n348 53.3664
R4833 w_13193_29093.n345 w_13193_29093.n343 53.3664
R4834 w_13193_29093.n1871 w_13193_29093.n1870 53.3664
R4835 w_13193_29093.n342 w_13193_29093.n340 53.3664
R4836 w_13193_29093.n1878 w_13193_29093.n1877 53.3664
R4837 w_13193_29093.n1885 w_13193_29093.n1884 53.3664
R4838 w_13193_29093.n1888 w_13193_29093.n1887 53.3664
R4839 w_13193_29093.n1893 w_13193_29093.n1892 53.3664
R4840 w_13193_29093.n1895 w_13193_29093.n334 53.3664
R4841 w_13193_29093.n2026 w_13193_29093.n2025 53.3664
R4842 w_13193_29093.n2038 w_13193_29093.n2037 53.3664
R4843 w_13193_29093.n2041 w_13193_29093.n2040 53.3664
R4844 w_13193_29093.n2053 w_13193_29093.n2052 53.3664
R4845 w_13193_29093.n2024 w_13193_29093.n1940 53.3664
R4846 w_13193_29093.n2020 w_13193_29093.n2019 53.3664
R4847 w_13193_29093.n2013 w_13193_29093.n1964 53.3664
R4848 w_13193_29093.n2012 w_13193_29093.n2011 53.3664
R4849 w_13193_29093.n2003 w_13193_29093.n2002 53.3664
R4850 w_13193_29093.n1998 w_13193_29093.n1970 53.3664
R4851 w_13193_29093.n1996 w_13193_29093.n1995 53.3664
R4852 w_13193_29093.n1991 w_13193_29093.n1973 53.3664
R4853 w_13193_29093.n1976 w_13193_29093.n1928 53.3664
R4854 w_13193_29093.n1981 w_13193_29093.n1980 53.3664
R4855 w_13193_29093.n1984 w_13193_29093.n1983 53.3664
R4856 w_13193_29093.n1989 w_13193_29093.n1988 53.3664
R4857 w_13193_29093.n1990 w_13193_29093.n1989 53.3664
R4858 w_13193_29093.n1983 w_13193_29093.n1974 53.3664
R4859 w_13193_29093.n1982 w_13193_29093.n1981 53.3664
R4860 w_13193_29093.n1977 w_13193_29093.n1976 53.3664
R4861 w_13193_29093.n1973 w_13193_29093.n1971 53.3664
R4862 w_13193_29093.n1997 w_13193_29093.n1996 53.3664
R4863 w_13193_29093.n1970 w_13193_29093.n1968 53.3664
R4864 w_13193_29093.n2004 w_13193_29093.n2003 53.3664
R4865 w_13193_29093.n2011 w_13193_29093.n2010 53.3664
R4866 w_13193_29093.n2014 w_13193_29093.n2013 53.3664
R4867 w_13193_29093.n2019 w_13193_29093.n2018 53.3664
R4868 w_13193_29093.n2021 w_13193_29093.n1940 53.3664
R4869 w_13193_29093.n2025 w_13193_29093.n1936 53.3664
R4870 w_13193_29093.n2039 w_13193_29093.n2038 53.3664
R4871 w_13193_29093.n2040 w_13193_29093.n1931 53.3664
R4872 w_13193_29093.n2054 w_13193_29093.n2053 53.3664
R4873 w_13193_29093.n1552 w_13193_29093.n1551 53.3664
R4874 w_13193_29093.n1555 w_13193_29093.n1554 53.3664
R4875 w_13193_29093.n1565 w_13193_29093.n1564 53.3664
R4876 w_13193_29093.n1568 w_13193_29093.n1567 53.3664
R4877 w_13193_29093.n578 w_13193_29093.n515 53.3664
R4878 w_13193_29093.n577 w_13193_29093.n576 53.3664
R4879 w_13193_29093.n570 w_13193_29093.n517 53.3664
R4880 w_13193_29093.n569 w_13193_29093.n568 53.3664
R4881 w_13193_29093.n560 w_13193_29093.n559 53.3664
R4882 w_13193_29093.n555 w_13193_29093.n523 53.3664
R4883 w_13193_29093.n553 w_13193_29093.n552 53.3664
R4884 w_13193_29093.n548 w_13193_29093.n526 53.3664
R4885 w_13193_29093.n533 w_13193_29093.n532 53.3664
R4886 w_13193_29093.n538 w_13193_29093.n537 53.3664
R4887 w_13193_29093.n541 w_13193_29093.n540 53.3664
R4888 w_13193_29093.n546 w_13193_29093.n545 53.3664
R4889 w_13193_29093.n547 w_13193_29093.n546 53.3664
R4890 w_13193_29093.n540 w_13193_29093.n527 53.3664
R4891 w_13193_29093.n539 w_13193_29093.n538 53.3664
R4892 w_13193_29093.n532 w_13193_29093.n529 53.3664
R4893 w_13193_29093.n526 w_13193_29093.n524 53.3664
R4894 w_13193_29093.n554 w_13193_29093.n553 53.3664
R4895 w_13193_29093.n523 w_13193_29093.n521 53.3664
R4896 w_13193_29093.n561 w_13193_29093.n560 53.3664
R4897 w_13193_29093.n568 w_13193_29093.n567 53.3664
R4898 w_13193_29093.n571 w_13193_29093.n570 53.3664
R4899 w_13193_29093.n576 w_13193_29093.n575 53.3664
R4900 w_13193_29093.n579 w_13193_29093.n578 53.3664
R4901 w_13193_29093.n1019 w_13193_29093.n1018 53.3664
R4902 w_13193_29093.n993 w_13193_29093.n921 53.3664
R4903 w_13193_29093.n989 w_13193_29093.n922 53.3664
R4904 w_13193_29093.n1005 w_13193_29093.n923 53.3664
R4905 w_13193_29093.n908 w_13193_29093.n906 53.3664
R4906 w_13193_29093.n930 w_13193_29093.n910 53.3664
R4907 w_13193_29093.n934 w_13193_29093.n912 53.3664
R4908 w_13193_29093.n938 w_13193_29093.n914 53.3664
R4909 w_13193_29093.n949 w_13193_29093.n920 53.3664
R4910 w_13193_29093.n953 w_13193_29093.n919 53.3664
R4911 w_13193_29093.n957 w_13193_29093.n918 53.3664
R4912 w_13193_29093.n961 w_13193_29093.n917 53.3664
R4913 w_13193_29093.n976 w_13193_29093.n909 53.3664
R4914 w_13193_29093.n973 w_13193_29093.n911 53.3664
R4915 w_13193_29093.n969 w_13193_29093.n913 53.3664
R4916 w_13193_29093.n965 w_13193_29093.n915 53.3664
R4917 w_13193_29093.n962 w_13193_29093.n915 53.3664
R4918 w_13193_29093.n966 w_13193_29093.n913 53.3664
R4919 w_13193_29093.n970 w_13193_29093.n911 53.3664
R4920 w_13193_29093.n974 w_13193_29093.n909 53.3664
R4921 w_13193_29093.n958 w_13193_29093.n917 53.3664
R4922 w_13193_29093.n954 w_13193_29093.n918 53.3664
R4923 w_13193_29093.n950 w_13193_29093.n919 53.3664
R4924 w_13193_29093.n946 w_13193_29093.n920 53.3664
R4925 w_13193_29093.n941 w_13193_29093.n914 53.3664
R4926 w_13193_29093.n937 w_13193_29093.n912 53.3664
R4927 w_13193_29093.n933 w_13193_29093.n910 53.3664
R4928 w_13193_29093.n929 w_13193_29093.n908 53.3664
R4929 w_13193_29093.n1018 w_13193_29093.n907 53.3664
R4930 w_13193_29093.n990 w_13193_29093.n921 53.3664
R4931 w_13193_29093.n1004 w_13193_29093.n922 53.3664
R4932 w_13193_29093.n925 w_13193_29093.n923 53.3664
R4933 w_13193_29093.n1460 w_13193_29093.n1459 53.3664
R4934 w_13193_29093.n618 w_13193_29093.n616 53.3664
R4935 w_13193_29093.n1481 w_13193_29093.n1480 53.3664
R4936 w_13193_29093.n1484 w_13193_29093.n1483 53.3664
R4937 w_13193_29093.n1458 w_13193_29093.n619 53.3664
R4938 w_13193_29093.n1454 w_13193_29093.n1453 53.3664
R4939 w_13193_29093.n1447 w_13193_29093.n1392 53.3664
R4940 w_13193_29093.n1446 w_13193_29093.n1445 53.3664
R4941 w_13193_29093.n1437 w_13193_29093.n1436 53.3664
R4942 w_13193_29093.n1432 w_13193_29093.n1398 53.3664
R4943 w_13193_29093.n1430 w_13193_29093.n1429 53.3664
R4944 w_13193_29093.n1425 w_13193_29093.n1401 53.3664
R4945 w_13193_29093.n1410 w_13193_29093.n1409 53.3664
R4946 w_13193_29093.n1415 w_13193_29093.n1414 53.3664
R4947 w_13193_29093.n1418 w_13193_29093.n1417 53.3664
R4948 w_13193_29093.n1423 w_13193_29093.n1422 53.3664
R4949 w_13193_29093.n1424 w_13193_29093.n1423 53.3664
R4950 w_13193_29093.n1417 w_13193_29093.n1402 53.3664
R4951 w_13193_29093.n1416 w_13193_29093.n1415 53.3664
R4952 w_13193_29093.n1409 w_13193_29093.n1404 53.3664
R4953 w_13193_29093.n1401 w_13193_29093.n1399 53.3664
R4954 w_13193_29093.n1431 w_13193_29093.n1430 53.3664
R4955 w_13193_29093.n1398 w_13193_29093.n1396 53.3664
R4956 w_13193_29093.n1438 w_13193_29093.n1437 53.3664
R4957 w_13193_29093.n1445 w_13193_29093.n1444 53.3664
R4958 w_13193_29093.n1448 w_13193_29093.n1447 53.3664
R4959 w_13193_29093.n1453 w_13193_29093.n1452 53.3664
R4960 w_13193_29093.n1455 w_13193_29093.n619 53.3664
R4961 w_13193_29093.n1461 w_13193_29093.n1460 53.3664
R4962 w_13193_29093.n616 w_13193_29093.n602 53.3664
R4963 w_13193_29093.n1482 w_13193_29093.n1481 53.3664
R4964 w_13193_29093.n1485 w_13193_29093.n1484 53.3664
R4965 w_13193_29093.n866 w_13193_29093.n801 53.3664
R4966 w_13193_29093.n869 w_13193_29093.n802 53.3664
R4967 w_13193_29093.n881 w_13193_29093.n803 53.3664
R4968 w_13193_29093.n894 w_13193_29093.n893 53.3664
R4969 w_13193_29093.n865 w_13193_29093.n788 53.3664
R4970 w_13193_29093.n861 w_13193_29093.n790 53.3664
R4971 w_13193_29093.n857 w_13193_29093.n792 53.3664
R4972 w_13193_29093.n853 w_13193_29093.n794 53.3664
R4973 w_13193_29093.n842 w_13193_29093.n800 53.3664
R4974 w_13193_29093.n838 w_13193_29093.n799 53.3664
R4975 w_13193_29093.n834 w_13193_29093.n798 53.3664
R4976 w_13193_29093.n830 w_13193_29093.n797 53.3664
R4977 w_13193_29093.n814 w_13193_29093.n789 53.3664
R4978 w_13193_29093.n818 w_13193_29093.n791 53.3664
R4979 w_13193_29093.n822 w_13193_29093.n793 53.3664
R4980 w_13193_29093.n826 w_13193_29093.n795 53.3664
R4981 w_13193_29093.n829 w_13193_29093.n795 53.3664
R4982 w_13193_29093.n825 w_13193_29093.n793 53.3664
R4983 w_13193_29093.n821 w_13193_29093.n791 53.3664
R4984 w_13193_29093.n817 w_13193_29093.n789 53.3664
R4985 w_13193_29093.n833 w_13193_29093.n797 53.3664
R4986 w_13193_29093.n837 w_13193_29093.n798 53.3664
R4987 w_13193_29093.n841 w_13193_29093.n799 53.3664
R4988 w_13193_29093.n845 w_13193_29093.n800 53.3664
R4989 w_13193_29093.n850 w_13193_29093.n794 53.3664
R4990 w_13193_29093.n854 w_13193_29093.n792 53.3664
R4991 w_13193_29093.n858 w_13193_29093.n790 53.3664
R4992 w_13193_29093.n862 w_13193_29093.n788 53.3664
R4993 w_13193_29093.n662 w_13193_29093.n654 53.3664
R4994 w_13193_29093.n1155 w_13193_29093.n1154 53.3664
R4995 w_13193_29093.n723 w_13193_29093.n655 53.3664
R4996 w_13193_29093.n730 w_13193_29093.n656 53.3664
R4997 w_13193_29093.n663 w_13193_29093.n641 53.3664
R4998 w_13193_29093.n667 w_13193_29093.n643 53.3664
R4999 w_13193_29093.n671 w_13193_29093.n645 53.3664
R5000 w_13193_29093.n675 w_13193_29093.n647 53.3664
R5001 w_13193_29093.n686 w_13193_29093.n653 53.3664
R5002 w_13193_29093.n690 w_13193_29093.n652 53.3664
R5003 w_13193_29093.n694 w_13193_29093.n651 53.3664
R5004 w_13193_29093.n698 w_13193_29093.n650 53.3664
R5005 w_13193_29093.n713 w_13193_29093.n642 53.3664
R5006 w_13193_29093.n710 w_13193_29093.n644 53.3664
R5007 w_13193_29093.n706 w_13193_29093.n646 53.3664
R5008 w_13193_29093.n702 w_13193_29093.n648 53.3664
R5009 w_13193_29093.n699 w_13193_29093.n648 53.3664
R5010 w_13193_29093.n703 w_13193_29093.n646 53.3664
R5011 w_13193_29093.n707 w_13193_29093.n644 53.3664
R5012 w_13193_29093.n711 w_13193_29093.n642 53.3664
R5013 w_13193_29093.n695 w_13193_29093.n650 53.3664
R5014 w_13193_29093.n691 w_13193_29093.n651 53.3664
R5015 w_13193_29093.n687 w_13193_29093.n652 53.3664
R5016 w_13193_29093.n683 w_13193_29093.n653 53.3664
R5017 w_13193_29093.n678 w_13193_29093.n647 53.3664
R5018 w_13193_29093.n674 w_13193_29093.n645 53.3664
R5019 w_13193_29093.n670 w_13193_29093.n643 53.3664
R5020 w_13193_29093.n666 w_13193_29093.n641 53.3664
R5021 w_13193_29093.n654 w_13193_29093.n639 53.3664
R5022 w_13193_29093.n1154 w_13193_29093.n640 53.3664
R5023 w_13193_29093.n729 w_13193_29093.n655 53.3664
R5024 w_13193_29093.n658 w_13193_29093.n656 53.3664
R5025 w_13193_29093.n870 w_13193_29093.n801 53.3664
R5026 w_13193_29093.n880 w_13193_29093.n802 53.3664
R5027 w_13193_29093.n804 w_13193_29093.n803 53.3664
R5028 w_13193_29093.n894 w_13193_29093.n786 53.3664
R5029 w_13193_29093.n1553 w_13193_29093.n1552 53.3664
R5030 w_13193_29093.n1554 w_13193_29093.n512 53.3664
R5031 w_13193_29093.n1566 w_13193_29093.n1565 53.3664
R5032 w_13193_29093.n1569 w_13193_29093.n1568 53.3664
R5033 w_13193_29093.n1298 w_13193_29093.n1297 53.3664
R5034 w_13193_29093.n1310 w_13193_29093.n1309 53.3664
R5035 w_13193_29093.n1313 w_13193_29093.n1312 53.3664
R5036 w_13193_29093.n1325 w_13193_29093.n1324 53.3664
R5037 w_13193_29093.n1296 w_13193_29093.n1230 53.3664
R5038 w_13193_29093.n1292 w_13193_29093.n1291 53.3664
R5039 w_13193_29093.n1285 w_13193_29093.n1236 53.3664
R5040 w_13193_29093.n1284 w_13193_29093.n1283 53.3664
R5041 w_13193_29093.n1275 w_13193_29093.n1274 53.3664
R5042 w_13193_29093.n1270 w_13193_29093.n1242 53.3664
R5043 w_13193_29093.n1268 w_13193_29093.n1267 53.3664
R5044 w_13193_29093.n1263 w_13193_29093.n1245 53.3664
R5045 w_13193_29093.n1248 w_13193_29093.n1218 53.3664
R5046 w_13193_29093.n1253 w_13193_29093.n1252 53.3664
R5047 w_13193_29093.n1256 w_13193_29093.n1255 53.3664
R5048 w_13193_29093.n1261 w_13193_29093.n1260 53.3664
R5049 w_13193_29093.n1262 w_13193_29093.n1261 53.3664
R5050 w_13193_29093.n1255 w_13193_29093.n1246 53.3664
R5051 w_13193_29093.n1254 w_13193_29093.n1253 53.3664
R5052 w_13193_29093.n1249 w_13193_29093.n1248 53.3664
R5053 w_13193_29093.n1245 w_13193_29093.n1243 53.3664
R5054 w_13193_29093.n1269 w_13193_29093.n1268 53.3664
R5055 w_13193_29093.n1242 w_13193_29093.n1240 53.3664
R5056 w_13193_29093.n1276 w_13193_29093.n1275 53.3664
R5057 w_13193_29093.n1283 w_13193_29093.n1282 53.3664
R5058 w_13193_29093.n1286 w_13193_29093.n1285 53.3664
R5059 w_13193_29093.n1291 w_13193_29093.n1290 53.3664
R5060 w_13193_29093.n1293 w_13193_29093.n1230 53.3664
R5061 w_13193_29093.n1297 w_13193_29093.n1226 53.3664
R5062 w_13193_29093.n1311 w_13193_29093.n1310 53.3664
R5063 w_13193_29093.n1312 w_13193_29093.n1221 53.3664
R5064 w_13193_29093.n1326 w_13193_29093.n1325 53.3664
R5065 w_13193_29093.n1905 w_13193_29093.n1904 53.3664
R5066 w_13193_29093.n1908 w_13193_29093.n1907 53.3664
R5067 w_13193_29093.n372 w_13193_29093.n371 53.3664
R5068 w_13193_29093.n373 w_13193_29093.n350 53.3664
R5069 w_13193_29093.n1668 w_13193_29093.n1667 53.3664
R5070 w_13193_29093.n1671 w_13193_29093.n1670 53.3664
R5071 w_13193_29093.n478 w_13193_29093.n465 53.3664
R5072 w_13193_29093.n1690 w_13193_29093.n1689 53.3664
R5073 w_13193_29093.n88 w_13193_29093.t307 48.0005
R5074 w_13193_29093.n88 w_13193_29093.t10 48.0005
R5075 w_13193_29093.n86 w_13193_29093.t8 48.0005
R5076 w_13193_29093.n86 w_13193_29093.t137 48.0005
R5077 w_13193_29093.n81 w_13193_29093.t312 48.0005
R5078 w_13193_29093.n81 w_13193_29093.t188 48.0005
R5079 w_13193_29093.n105 w_13193_29093.t290 48.0005
R5080 w_13193_29093.n105 w_13193_29093.t40 48.0005
R5081 w_13193_29093.n113 w_13193_29093.t34 48.0005
R5082 w_13193_29093.n113 w_13193_29093.t247 48.0005
R5083 w_13193_29093.n125 w_13193_29093.t119 48.0005
R5084 w_13193_29093.n125 w_13193_29093.t20 48.0005
R5085 w_13193_29093.n72 w_13193_29093.t16 48.0005
R5086 w_13193_29093.n72 w_13193_29093.t44 48.0005
R5087 w_13193_29093.n141 w_13193_29093.t173 48.0005
R5088 w_13193_29093.n141 w_13193_29093.t217 48.0005
R5089 w_13193_29093.n144 w_13193_29093.t181 48.0005
R5090 w_13193_29093.n144 w_13193_29093.t42 48.0005
R5091 w_13193_29093.n150 w_13193_29093.t309 48.0005
R5092 w_13193_29093.n150 w_13193_29093.t223 48.0005
R5093 w_13193_29093.n153 w_13193_29093.t204 48.0005
R5094 w_13193_29093.n153 w_13193_29093.t190 48.0005
R5095 w_13193_29093.n156 w_13193_29093.t299 48.0005
R5096 w_13193_29093.n156 w_13193_29093.t285 48.0005
R5097 w_13193_29093.n162 w_13193_29093.t106 48.0005
R5098 w_13193_29093.n162 w_13193_29093.t273 48.0005
R5099 w_13193_29093.n163 w_13193_29093.t275 48.0005
R5100 w_13193_29093.n163 w_13193_29093.t277 48.0005
R5101 w_13193_29093.n168 w_13193_29093.t165 48.0005
R5102 w_13193_29093.n168 w_13193_29093.t123 48.0005
R5103 w_13193_29093.n173 w_13193_29093.t251 48.0005
R5104 w_13193_29093.n173 w_13193_29093.t305 48.0005
R5105 w_13193_29093.n176 w_13193_29093.t30 48.0005
R5106 w_13193_29093.n176 w_13193_29093.t236 48.0005
R5107 w_13193_29093.n180 w_13193_29093.t161 48.0005
R5108 w_13193_29093.n180 w_13193_29093.t121 48.0005
R5109 w_13193_29093.n185 w_13193_29093.t301 48.0005
R5110 w_13193_29093.n185 w_13193_29093.t127 48.0005
R5111 w_13193_29093.n188 w_13193_29093.t167 48.0005
R5112 w_13193_29093.n188 w_13193_29093.t109 48.0005
R5113 w_13193_29093.n2581 w_13193_29093.t153 48.0005
R5114 w_13193_29093.n2581 w_13193_29093.t135 48.0005
R5115 w_13193_29093.n2697 w_13193_29093.t306 47.9388
R5116 w_13193_29093.t47 w_13193_29093.n20 47.7166
R5117 w_13193_29093.n635 w_13193_29093.t107 47.7166
R5118 w_13193_29093.t130 w_13193_29093.n735 47.7166
R5119 w_13193_29093.n1079 w_13193_29093.n781 47.7166
R5120 w_13193_29093.t156 w_13193_29093.t136 47.5681
R5121 w_13193_29093.t254 w_13193_29093.t261 47.5681
R5122 w_13193_29093.t53 w_13193_29093.n14 47.5454
R5123 w_13193_29093.t53 w_13193_29093.n23 47.5454
R5124 w_13193_29093.t126 w_13193_29093.n63 44.4949
R5125 w_13193_29093.t203 w_13193_29093.n2388 42.9693
R5126 w_13193_29093.n2387 w_13193_29093.t132 42.9693
R5127 w_13193_29093.n2532 w_13193_29093.t29 42.9693
R5128 w_13193_29093.n2530 w_13193_29093.t300 42.9693
R5129 w_13193_29093.t53 w_13193_29093.t131 42.7252
R5130 w_13193_29093.n2756 w_13193_29093.n34 39.5027
R5131 w_13193_29093.n2726 w_13193_29093.n54 39.4985
R5132 w_13193_29093.n2764 w_13193_29093.t269 39.3565
R5133 w_13193_29093.t212 w_13193_29093.n1160 39.0409
R5134 w_13193_29093.n718 w_13193_29093.t21 39.0409
R5135 w_13193_29093.n1148 w_13193_29093.t133 39.0409
R5136 w_13193_29093.n1146 w_13193_29093.t295 39.0409
R5137 w_13193_29093.n1025 w_13193_29093.t22 37.595
R5138 w_13193_29093.n2700 w_13193_29093.n2699 36.8449
R5139 w_13193_29093.n2438 w_13193_29093.t9 35.6762
R5140 w_13193_29093.n2696 w_13193_29093.t302 35.6762
R5141 w_13193_29093.n2546 w_13193_29093.n2545 35.6576
R5142 w_13193_29093.n2565 w_13193_29093.n197 35.6576
R5143 w_13193_29093.n2540 w_13193_29093.n2539 35.6576
R5144 w_13193_29093.n2537 w_13193_29093.n193 35.6576
R5145 w_13193_29093.t53 w_13193_29093.t242 34.9571
R5146 w_13193_29093.t53 w_13193_29093.n20 34.7031
R5147 w_13193_29093.t53 w_13193_29093.n17 34.4319
R5148 w_13193_29093.n2549 w_13193_29093.n203 34.3278
R5149 w_13193_29093.n2554 w_13193_29093.n2553 34.3278
R5150 w_13193_29093.t53 w_13193_29093.n27 33.9847
R5151 w_13193_29093.n1023 w_13193_29093.t149 33.2572
R5152 w_13193_29093.n999 w_13193_29093.t219 33.2572
R5153 w_13193_29093.t23 w_13193_29093.n1011 33.2572
R5154 w_13193_29093.n774 w_13193_29093.n769 33.0535
R5155 w_13193_29093.n258 w_13193_29093.n257 32.3962
R5156 w_13193_29093.n2483 w_13193_29093.n2482 32.0005
R5157 w_13193_29093.n2484 w_13193_29093.n2483 32.0005
R5158 w_13193_29093.n2488 w_13193_29093.n219 32.0005
R5159 w_13193_29093.n2489 w_13193_29093.n2488 32.0005
R5160 w_13193_29093.n2490 w_13193_29093.n2489 32.0005
R5161 w_13193_29093.n2495 w_13193_29093.n2494 32.0005
R5162 w_13193_29093.n2511 w_13193_29093.n213 32.0005
R5163 w_13193_29093.n2513 w_13193_29093.n2511 32.0005
R5164 w_13193_29093.n2514 w_13193_29093.n211 32.0005
R5165 w_13193_29093.n2518 w_13193_29093.n211 32.0005
R5166 w_13193_29093.n2519 w_13193_29093.n2518 32.0005
R5167 w_13193_29093.n2478 w_13193_29093.n2477 32.0005
R5168 w_13193_29093.n2478 w_13193_29093.n234 32.0005
R5169 w_13193_29093.n2471 w_13193_29093.n238 32.0005
R5170 w_13193_29093.n2475 w_13193_29093.n238 32.0005
R5171 w_13193_29093.n2469 w_13193_29093.n241 32.0005
R5172 w_13193_29093.n92 w_13193_29093.n91 32.0005
R5173 w_13193_29093.n93 w_13193_29093.n92 32.0005
R5174 w_13193_29093.n93 w_13193_29093.n84 32.0005
R5175 w_13193_29093.n98 w_13193_29093.n97 32.0005
R5176 w_13193_29093.n99 w_13193_29093.n98 32.0005
R5177 w_13193_29093.n99 w_13193_29093.n82 32.0005
R5178 w_13193_29093.n104 w_13193_29093.n103 32.0005
R5179 w_13193_29093.n107 w_13193_29093.n79 32.0005
R5180 w_13193_29093.n111 w_13193_29093.n79 32.0005
R5181 w_13193_29093.n112 w_13193_29093.n111 32.0005
R5182 w_13193_29093.n114 w_13193_29093.n77 32.0005
R5183 w_13193_29093.n118 w_13193_29093.n77 32.0005
R5184 w_13193_29093.n119 w_13193_29093.n118 32.0005
R5185 w_13193_29093.n120 w_13193_29093.n119 32.0005
R5186 w_13193_29093.n120 w_13193_29093.n75 32.0005
R5187 w_13193_29093.n124 w_13193_29093.n75 32.0005
R5188 w_13193_29093.n128 w_13193_29093.n127 32.0005
R5189 w_13193_29093.n132 w_13193_29093.n73 32.0005
R5190 w_13193_29093.n133 w_13193_29093.n132 32.0005
R5191 w_13193_29093.n134 w_13193_29093.n133 32.0005
R5192 w_13193_29093.n134 w_13193_29093.n69 32.0005
R5193 w_13193_29093.n2690 w_13193_29093.n70 32.0005
R5194 w_13193_29093.n2686 w_13193_29093.n70 32.0005
R5195 w_13193_29093.n2686 w_13193_29093.n2685 32.0005
R5196 w_13193_29093.n2683 w_13193_29093.n139 32.0005
R5197 w_13193_29093.n2679 w_13193_29093.n139 32.0005
R5198 w_13193_29093.n2677 w_13193_29093.n2676 32.0005
R5199 w_13193_29093.n2672 w_13193_29093.n2671 32.0005
R5200 w_13193_29093.n2669 w_13193_29093.n145 32.0005
R5201 w_13193_29093.n2665 w_13193_29093.n145 32.0005
R5202 w_13193_29093.n2663 w_13193_29093.n2662 32.0005
R5203 w_13193_29093.n2662 w_13193_29093.n148 32.0005
R5204 w_13193_29093.n2658 w_13193_29093.n148 32.0005
R5205 w_13193_29093.n2658 w_13193_29093.n2657 32.0005
R5206 w_13193_29093.n2657 w_13193_29093.n2656 32.0005
R5207 w_13193_29093.n2656 w_13193_29093.n151 32.0005
R5208 w_13193_29093.n2652 w_13193_29093.n2651 32.0005
R5209 w_13193_29093.n2649 w_13193_29093.n154 32.0005
R5210 w_13193_29093.n2645 w_13193_29093.n154 32.0005
R5211 w_13193_29093.n2645 w_13193_29093.n2644 32.0005
R5212 w_13193_29093.n2644 w_13193_29093.n2643 32.0005
R5213 w_13193_29093.n2639 w_13193_29093.n2638 32.0005
R5214 w_13193_29093.n2636 w_13193_29093.n160 32.0005
R5215 w_13193_29093.n2632 w_13193_29093.n160 32.0005
R5216 w_13193_29093.n2631 w_13193_29093.n2630 32.0005
R5217 w_13193_29093.n2627 w_13193_29093.n2626 32.0005
R5218 w_13193_29093.n2626 w_13193_29093.n2625 32.0005
R5219 w_13193_29093.n2625 w_13193_29093.n166 32.0005
R5220 w_13193_29093.n2621 w_13193_29093.n166 32.0005
R5221 w_13193_29093.n2619 w_13193_29093.n169 32.0005
R5222 w_13193_29093.n2615 w_13193_29093.n2614 32.0005
R5223 w_13193_29093.n2614 w_13193_29093.n2613 32.0005
R5224 w_13193_29093.n2612 w_13193_29093.n174 32.0005
R5225 w_13193_29093.n2608 w_13193_29093.n2607 32.0005
R5226 w_13193_29093.n2607 w_13193_29093.n2606 32.0005
R5227 w_13193_29093.n2606 w_13193_29093.n178 32.0005
R5228 w_13193_29093.n2602 w_13193_29093.n178 32.0005
R5229 w_13193_29093.n2600 w_13193_29093.n181 32.0005
R5230 w_13193_29093.n2596 w_13193_29093.n2595 32.0005
R5231 w_13193_29093.n2595 w_13193_29093.n2594 32.0005
R5232 w_13193_29093.n2593 w_13193_29093.n186 32.0005
R5233 w_13193_29093.n2589 w_13193_29093.n2588 32.0005
R5234 w_13193_29093.n2588 w_13193_29093.n2587 32.0005
R5235 w_13193_29093.n2587 w_13193_29093.n190 32.0005
R5236 w_13193_29093.n2583 w_13193_29093.n190 32.0005
R5237 w_13193_29093.n2564 w_13193_29093.n198 32.0005
R5238 w_13193_29093.n2560 w_13193_29093.n198 32.0005
R5239 w_13193_29093.n2560 w_13193_29093.n2559 32.0005
R5240 w_13193_29093.n2559 w_13193_29093.n2558 32.0005
R5241 w_13193_29093.n2558 w_13193_29093.n200 32.0005
R5242 w_13193_29093.n2572 w_13193_29093.n2571 32.0005
R5243 w_13193_29093.n2571 w_13193_29093.n2570 32.0005
R5244 w_13193_29093.n2570 w_13193_29093.n195 32.0005
R5245 w_13193_29093.n2566 w_13193_29093.n195 32.0005
R5246 w_13193_29093.n2566 w_13193_29093.n2565 32.0005
R5247 w_13193_29093.n2577 w_13193_29093.n2576 32.0005
R5248 w_13193_29093.n2576 w_13193_29093.n193 32.0005
R5249 w_13193_29093.n2344 w_13193_29093.n2343 32.0005
R5250 w_13193_29093.n2349 w_13193_29093.n2348 32.0005
R5251 w_13193_29093.n2354 w_13193_29093.n2229 32.0005
R5252 w_13193_29093.n2356 w_13193_29093.n2355 32.0005
R5253 w_13193_29093.n2356 w_13193_29093.n2227 32.0005
R5254 w_13193_29093.n2432 w_13193_29093.n2227 32.0005
R5255 w_13193_29093.n2431 w_13193_29093.n2360 32.0005
R5256 w_13193_29093.n2427 w_13193_29093.n2360 32.0005
R5257 w_13193_29093.n2425 w_13193_29093.n2424 32.0005
R5258 w_13193_29093.n2424 w_13193_29093.n2362 32.0005
R5259 w_13193_29093.n2420 w_13193_29093.n2419 32.0005
R5260 w_13193_29093.n2419 w_13193_29093.n2418 32.0005
R5261 w_13193_29093.n2418 w_13193_29093.n2364 32.0005
R5262 w_13193_29093.n2414 w_13193_29093.n2364 32.0005
R5263 w_13193_29093.n2413 w_13193_29093.n2412 32.0005
R5264 w_13193_29093.n2412 w_13193_29093.n2367 32.0005
R5265 w_13193_29093.n2408 w_13193_29093.n2367 32.0005
R5266 w_13193_29093.n2408 w_13193_29093.n2407 32.0005
R5267 w_13193_29093.n2407 w_13193_29093.n2369 32.0005
R5268 w_13193_29093.n2403 w_13193_29093.n2369 32.0005
R5269 w_13193_29093.n2401 w_13193_29093.n2372 32.0005
R5270 w_13193_29093.n2397 w_13193_29093.n2372 32.0005
R5271 w_13193_29093.n2397 w_13193_29093.n2396 32.0005
R5272 w_13193_29093.n2396 w_13193_29093.n2395 32.0005
R5273 w_13193_29093.n2395 w_13193_29093.n2374 32.0005
R5274 w_13193_29093.n2338 w_13193_29093.n2337 32.0005
R5275 w_13193_29093.n2335 w_13193_29093.n2237 32.0005
R5276 w_13193_29093.n2330 w_13193_29093.n2329 32.0005
R5277 w_13193_29093.n2302 w_13193_29093.n2268 32.0005
R5278 w_13193_29093.n2298 w_13193_29093.n2268 32.0005
R5279 w_13193_29093.n2297 w_13193_29093.n2296 32.0005
R5280 w_13193_29093.n2296 w_13193_29093.n2271 32.0005
R5281 w_13193_29093.n2292 w_13193_29093.n2271 32.0005
R5282 w_13193_29093.n2290 w_13193_29093.n2289 32.0005
R5283 w_13193_29093.n2289 w_13193_29093.n2274 32.0005
R5284 w_13193_29093.n2284 w_13193_29093.n2283 32.0005
R5285 w_13193_29093.n2283 w_13193_29093.n2219 32.0005
R5286 w_13193_29093.n2448 w_13193_29093.n2219 32.0005
R5287 w_13193_29093.n2450 w_13193_29093.n2449 32.0005
R5288 w_13193_29093.n2450 w_13193_29093.n2217 32.0005
R5289 w_13193_29093.n2457 w_13193_29093.n2454 32.0005
R5290 w_13193_29093.n2454 w_13193_29093.n2215 32.0005
R5291 w_13193_29093.n2324 w_13193_29093.n2253 32.0005
R5292 w_13193_29093.n2322 w_13193_29093.n2255 32.0005
R5293 w_13193_29093.n2317 w_13193_29093.n2316 32.0005
R5294 w_13193_29093.n2304 w_13193_29093.n2303 32.0005
R5295 w_13193_29093.n2309 w_13193_29093.n2264 32.0005
R5296 w_13193_29093.n2311 w_13193_29093.n2262 32.0005
R5297 w_13193_29093.n2756 w_13193_29093.n2755 32.0005
R5298 w_13193_29093.n2755 w_13193_29093.n2754 32.0005
R5299 w_13193_29093.n2754 w_13193_29093.n36 32.0005
R5300 w_13193_29093.n2750 w_13193_29093.n2749 32.0005
R5301 w_13193_29093.n2749 w_13193_29093.n2748 32.0005
R5302 w_13193_29093.n2748 w_13193_29093.n42 32.0005
R5303 w_13193_29093.n2744 w_13193_29093.n42 32.0005
R5304 w_13193_29093.n2744 w_13193_29093.n2743 32.0005
R5305 w_13193_29093.n2743 w_13193_29093.n2742 32.0005
R5306 w_13193_29093.n2742 w_13193_29093.n46 32.0005
R5307 w_13193_29093.n2738 w_13193_29093.n46 32.0005
R5308 w_13193_29093.n2738 w_13193_29093.n2737 32.0005
R5309 w_13193_29093.n2737 w_13193_29093.n2736 32.0005
R5310 w_13193_29093.n2736 w_13193_29093.n50 32.0005
R5311 w_13193_29093.n2732 w_13193_29093.n50 32.0005
R5312 w_13193_29093.n2732 w_13193_29093.n2731 32.0005
R5313 w_13193_29093.n2731 w_13193_29093.n2730 32.0005
R5314 w_13193_29093.n2730 w_13193_29093.n54 32.0005
R5315 w_13193_29093.n2578 w_13193_29093.n2577 29.4625
R5316 w_13193_29093.n260 w_13193_29093.t178 29.131
R5317 w_13193_29093.n234 w_13193_29093.n233 29.0291
R5318 w_13193_29093.n2507 w_13193_29093.n2506 29.0291
R5319 w_13193_29093.t53 w_13193_29093.t21 28.9193
R5320 w_13193_29093.t295 w_13193_29093.t263 28.9193
R5321 w_13193_29093.t22 w_13193_29093.t265 28.9193
R5322 w_13193_29093.t53 w_13193_29093.t219 28.9193
R5323 w_13193_29093.t53 w_13193_29093.n28 28.9193
R5324 w_13193_29093.n2685 w_13193_29093.n2684 28.8005
R5325 w_13193_29093.n2676 w_13193_29093.n142 28.8005
R5326 w_13193_29093.n2643 w_13193_29093.n157 28.8005
R5327 w_13193_29093.n2620 w_13193_29093.n2619 28.8005
R5328 w_13193_29093.n2601 w_13193_29093.n2600 28.8005
R5329 w_13193_29093.n2285 w_13193_29093.n2284 28.8005
R5330 w_13193_29093.n2458 w_13193_29093.n2217 28.8005
R5331 w_13193_29093.n1619 w_13193_29093.n1599 27.5561
R5332 w_13193_29093.n1866 w_13193_29093.n344 27.5561
R5333 w_13193_29093.n1992 w_13193_29093.n1972 27.5561
R5334 w_13193_29093.n549 w_13193_29093.n525 27.5561
R5335 w_13193_29093.n963 w_13193_29093.n960 27.5561
R5336 w_13193_29093.n1426 w_13193_29093.n1400 27.5561
R5337 w_13193_29093.n831 w_13193_29093.n828 27.5561
R5338 w_13193_29093.n700 w_13193_29093.n697 27.5561
R5339 w_13193_29093.n1264 w_13193_29093.n1244 27.5561
R5340 w_13193_29093.n2718 w_13193_29093.n2717 27.2005
R5341 w_13193_29093.n2723 w_13193_29093.n2722 27.2005
R5342 w_13193_29093.n1635 w_13193_29093.n1634 26.6672
R5343 w_13193_29093.n1882 w_13193_29093.n1881 26.6672
R5344 w_13193_29093.n2008 w_13193_29093.n2007 26.6672
R5345 w_13193_29093.n565 w_13193_29093.n564 26.6672
R5346 w_13193_29093.n944 w_13193_29093.n943 26.6672
R5347 w_13193_29093.n1442 w_13193_29093.n1441 26.6672
R5348 w_13193_29093.n848 w_13193_29093.n847 26.6672
R5349 w_13193_29093.n681 w_13193_29093.n680 26.6672
R5350 w_13193_29093.n1280 w_13193_29093.n1279 26.6672
R5351 w_13193_29093.t105 w_13193_29093.t116 25.7817
R5352 w_13193_29093.t274 w_13193_29093.t101 25.7817
R5353 w_13193_29093.t67 w_13193_29093.t250 25.7817
R5354 w_13193_29093.n2507 w_13193_29093.n2495 25.6005
R5355 w_13193_29093.n2471 w_13193_29093.n2470 25.6005
R5356 w_13193_29093.n2476 w_13193_29093.n2475 25.6005
R5357 w_13193_29093.n2554 w_13193_29093.n200 25.6005
R5358 w_13193_29093.n2344 w_13193_29093.n2231 25.6005
R5359 w_13193_29093.n2348 w_13193_29093.n2231 25.6005
R5360 w_13193_29093.n2350 w_13193_29093.n2349 25.6005
R5361 w_13193_29093.n2350 w_13193_29093.n2229 25.6005
R5362 w_13193_29093.n2403 w_13193_29093.n2402 25.6005
R5363 w_13193_29093.n2402 w_13193_29093.n2401 25.6005
R5364 w_13193_29093.n2337 w_13193_29093.n2336 25.6005
R5365 w_13193_29093.n2331 w_13193_29093.n2237 25.6005
R5366 w_13193_29093.n2336 w_13193_29093.n2335 25.6005
R5367 w_13193_29093.n2331 w_13193_29093.n2330 25.6005
R5368 w_13193_29093.n2463 w_13193_29093.n2215 25.6005
R5369 w_13193_29093.n2324 w_13193_29093.n2323 25.6005
R5370 w_13193_29093.n2323 w_13193_29093.n2322 25.6005
R5371 w_13193_29093.n2318 w_13193_29093.n2255 25.6005
R5372 w_13193_29093.n2318 w_13193_29093.n2317 25.6005
R5373 w_13193_29093.n2305 w_13193_29093.n2304 25.6005
R5374 w_13193_29093.n2310 w_13193_29093.n2309 25.6005
R5375 w_13193_29093.n2305 w_13193_29093.n2264 25.6005
R5376 w_13193_29093.n2311 w_13193_29093.n2310 25.6005
R5377 w_13193_29093.n2708 w_13193_29093.n2707 25.6005
R5378 w_13193_29093.n2716 w_13193_29093.n2715 25.6005
R5379 w_13193_29093.n257 w_13193_29093.n243 25.3679
R5380 w_13193_29093.t115 w_13193_29093.n2535 24.7196
R5381 w_13193_29093.n55 w_13193_29093.t227 24.0005
R5382 w_13193_29093.n55 w_13193_29093.t91 24.0005
R5383 w_13193_29093.n51 w_13193_29093.t182 24.0005
R5384 w_13193_29093.n51 w_13193_29093.t280 24.0005
R5385 w_13193_29093.n47 w_13193_29093.t28 24.0005
R5386 w_13193_29093.n47 w_13193_29093.t171 24.0005
R5387 w_13193_29093.n43 w_13193_29093.t279 24.0005
R5388 w_13193_29093.n43 w_13193_29093.t14 24.0005
R5389 w_13193_29093.n37 w_13193_29093.t62 24.0005
R5390 w_13193_29093.n37 w_13193_29093.t226 24.0005
R5391 w_13193_29093.t113 w_13193_29093.t216 23.7843
R5392 w_13193_29093.n2580 w_13193_29093.n2579 23.1805
R5393 w_13193_29093.n91 w_13193_29093.n87 22.4005
R5394 w_13193_29093.n2684 w_13193_29093.n2683 22.4005
R5395 w_13193_29093.n2672 w_13193_29093.n142 22.4005
R5396 w_13193_29093.n2639 w_13193_29093.n157 22.4005
R5397 w_13193_29093.n2621 w_13193_29093.n2620 22.4005
R5398 w_13193_29093.n2602 w_13193_29093.n2601 22.4005
R5399 w_13193_29093.n2583 w_13193_29093.n2582 22.4005
R5400 w_13193_29093.n2285 w_13193_29093.n2274 22.4005
R5401 w_13193_29093.n2458 w_13193_29093.n2457 22.4005
R5402 w_13193_29093.n2710 w_13193_29093.n57 22.4005
R5403 w_13193_29093.n2760 w_13193_29093.n2759 22.4005
R5404 w_13193_29093.t53 w_13193_29093.t183 21.1922
R5405 w_13193_29093.n2523 w_13193_29093.n2522 20.9665
R5406 w_13193_29093.n2490 w_13193_29093.n216 19.2005
R5407 w_13193_29093.n2494 w_13193_29093.n216 19.2005
R5408 w_13193_29093.n97 w_13193_29093.n84 19.2005
R5409 w_13193_29093.n103 w_13193_29093.n82 19.2005
R5410 w_13193_29093.n114 w_13193_29093.n112 19.2005
R5411 w_13193_29093.n128 w_13193_29093.n73 19.2005
R5412 w_13193_29093.n2652 w_13193_29093.n151 19.2005
R5413 w_13193_29093.n2632 w_13193_29093.n2631 19.2005
R5414 w_13193_29093.n2613 w_13193_29093.n2612 19.2005
R5415 w_13193_29093.n2594 w_13193_29093.n2593 19.2005
R5416 w_13193_29093.n2355 w_13193_29093.n2354 19.2005
R5417 w_13193_29093.n2432 w_13193_29093.n2431 19.2005
R5418 w_13193_29093.n2420 w_13193_29093.n2362 19.2005
R5419 w_13193_29093.n2414 w_13193_29093.n2413 19.2005
R5420 w_13193_29093.n2391 w_13193_29093.n2374 19.2005
R5421 w_13193_29093.n2343 w_13193_29093.n2341 19.2005
R5422 w_13193_29093.n2303 w_13193_29093.n2302 19.2005
R5423 w_13193_29093.n2298 w_13193_29093.n2297 19.2005
R5424 w_13193_29093.n2449 w_13193_29093.n2448 19.2005
R5425 w_13193_29093.n2316 w_13193_29093.n2315 19.2005
R5426 w_13193_29093.n2315 w_13193_29093.n2262 19.2005
R5427 w_13193_29093.n2750 w_13193_29093.n36 19.2005
R5428 w_13193_29093.n2158 w_13193_29093.n2157 17.5843
R5429 w_13193_29093.n1190 w_13193_29093.n1186 17.5843
R5430 w_13193_29093.n2131 w_13193_29093.n2130 17.5843
R5431 w_13193_29093.n1781 w_13193_29093.n1780 17.0672
R5432 w_13193_29093.n1752 w_13193_29093.n446 17.0672
R5433 w_13193_29093.n1721 w_13193_29093.n1720 17.0672
R5434 w_13193_29093.n2199 w_13193_29093.n2198 16.9605
R5435 w_13193_29093.n1838 w_13193_29093.n1837 16.7235
R5436 w_13193_29093.n1383 w_13193_29093.n1382 16.7235
R5437 w_13193_29093.n583 w_13193_29093.n495 16.7235
R5438 w_13193_29093.n2108 w_13193_29093.n2107 16.7235
R5439 w_13193_29093.n2578 w_13193_29093.n192 16.0525
R5440 w_13193_29093.n2670 w_13193_29093.n2669 16.0005
R5441 w_13193_29093.n2638 w_13193_29093.n2637 16.0005
R5442 w_13193_29093.n171 w_13193_29093.n169 16.0005
R5443 w_13193_29093.n183 w_13193_29093.n181 16.0005
R5444 w_13193_29093.n2341 w_13193_29093.n2234 16.0005
R5445 w_13193_29093.n1694 w_13193_29093.n461 16.0005
R5446 w_13193_29093.n1605 w_13193_29093.n461 16.0005
R5447 w_13193_29093.n1606 w_13193_29093.n1605 16.0005
R5448 w_13193_29093.n1606 w_13193_29093.n1602 16.0005
R5449 w_13193_29093.n1612 w_13193_29093.n1602 16.0005
R5450 w_13193_29093.n1613 w_13193_29093.n1612 16.0005
R5451 w_13193_29093.n1614 w_13193_29093.n1613 16.0005
R5452 w_13193_29093.n1614 w_13193_29093.n1599 16.0005
R5453 w_13193_29093.n1634 w_13193_29093.n1594 16.0005
R5454 w_13193_29093.n1628 w_13193_29093.n1594 16.0005
R5455 w_13193_29093.n1628 w_13193_29093.n1627 16.0005
R5456 w_13193_29093.n1627 w_13193_29093.n1626 16.0005
R5457 w_13193_29093.n1626 w_13193_29093.n1596 16.0005
R5458 w_13193_29093.n1621 w_13193_29093.n1596 16.0005
R5459 w_13193_29093.n1621 w_13193_29093.n1620 16.0005
R5460 w_13193_29093.n1620 w_13193_29093.n1619 16.0005
R5461 w_13193_29093.n1651 w_13193_29093.n1650 16.0005
R5462 w_13193_29093.n1650 w_13193_29093.n1590 16.0005
R5463 w_13193_29093.n1644 w_13193_29093.n1590 16.0005
R5464 w_13193_29093.n1644 w_13193_29093.n1643 16.0005
R5465 w_13193_29093.n1643 w_13193_29093.n1642 16.0005
R5466 w_13193_29093.n1642 w_13193_29093.n1592 16.0005
R5467 w_13193_29093.n1636 w_13193_29093.n1592 16.0005
R5468 w_13193_29093.n1636 w_13193_29093.n1635 16.0005
R5469 w_13193_29093.n1851 w_13193_29093.n349 16.0005
R5470 w_13193_29093.n1852 w_13193_29093.n1851 16.0005
R5471 w_13193_29093.n1853 w_13193_29093.n1852 16.0005
R5472 w_13193_29093.n1853 w_13193_29093.n347 16.0005
R5473 w_13193_29093.n1859 w_13193_29093.n347 16.0005
R5474 w_13193_29093.n1860 w_13193_29093.n1859 16.0005
R5475 w_13193_29093.n1861 w_13193_29093.n1860 16.0005
R5476 w_13193_29093.n1861 w_13193_29093.n344 16.0005
R5477 w_13193_29093.n1881 w_13193_29093.n339 16.0005
R5478 w_13193_29093.n1875 w_13193_29093.n339 16.0005
R5479 w_13193_29093.n1875 w_13193_29093.n1874 16.0005
R5480 w_13193_29093.n1874 w_13193_29093.n1873 16.0005
R5481 w_13193_29093.n1873 w_13193_29093.n341 16.0005
R5482 w_13193_29093.n1868 w_13193_29093.n341 16.0005
R5483 w_13193_29093.n1868 w_13193_29093.n1867 16.0005
R5484 w_13193_29093.n1867 w_13193_29093.n1866 16.0005
R5485 w_13193_29093.n1897 w_13193_29093.n1896 16.0005
R5486 w_13193_29093.n1896 w_13193_29093.n335 16.0005
R5487 w_13193_29093.n1891 w_13193_29093.n335 16.0005
R5488 w_13193_29093.n1891 w_13193_29093.n1890 16.0005
R5489 w_13193_29093.n1890 w_13193_29093.n1889 16.0005
R5490 w_13193_29093.n1889 w_13193_29093.n337 16.0005
R5491 w_13193_29093.n1883 w_13193_29093.n337 16.0005
R5492 w_13193_29093.n1883 w_13193_29093.n1882 16.0005
R5493 w_13193_29093.n2058 w_13193_29093.n1927 16.0005
R5494 w_13193_29093.n1978 w_13193_29093.n1927 16.0005
R5495 w_13193_29093.n1979 w_13193_29093.n1978 16.0005
R5496 w_13193_29093.n1979 w_13193_29093.n1975 16.0005
R5497 w_13193_29093.n1985 w_13193_29093.n1975 16.0005
R5498 w_13193_29093.n1986 w_13193_29093.n1985 16.0005
R5499 w_13193_29093.n1987 w_13193_29093.n1986 16.0005
R5500 w_13193_29093.n1987 w_13193_29093.n1972 16.0005
R5501 w_13193_29093.n2007 w_13193_29093.n1967 16.0005
R5502 w_13193_29093.n2001 w_13193_29093.n1967 16.0005
R5503 w_13193_29093.n2001 w_13193_29093.n2000 16.0005
R5504 w_13193_29093.n2000 w_13193_29093.n1999 16.0005
R5505 w_13193_29093.n1999 w_13193_29093.n1969 16.0005
R5506 w_13193_29093.n1994 w_13193_29093.n1969 16.0005
R5507 w_13193_29093.n1994 w_13193_29093.n1993 16.0005
R5508 w_13193_29093.n1993 w_13193_29093.n1992 16.0005
R5509 w_13193_29093.n2023 w_13193_29093.n2022 16.0005
R5510 w_13193_29093.n2022 w_13193_29093.n1963 16.0005
R5511 w_13193_29093.n2017 w_13193_29093.n1963 16.0005
R5512 w_13193_29093.n2017 w_13193_29093.n2016 16.0005
R5513 w_13193_29093.n2016 w_13193_29093.n2015 16.0005
R5514 w_13193_29093.n2015 w_13193_29093.n1965 16.0005
R5515 w_13193_29093.n2009 w_13193_29093.n1965 16.0005
R5516 w_13193_29093.n2009 w_13193_29093.n2008 16.0005
R5517 w_13193_29093.n534 w_13193_29093.n453 16.0005
R5518 w_13193_29093.n535 w_13193_29093.n534 16.0005
R5519 w_13193_29093.n536 w_13193_29093.n535 16.0005
R5520 w_13193_29093.n536 w_13193_29093.n528 16.0005
R5521 w_13193_29093.n542 w_13193_29093.n528 16.0005
R5522 w_13193_29093.n543 w_13193_29093.n542 16.0005
R5523 w_13193_29093.n544 w_13193_29093.n543 16.0005
R5524 w_13193_29093.n544 w_13193_29093.n525 16.0005
R5525 w_13193_29093.n564 w_13193_29093.n520 16.0005
R5526 w_13193_29093.n558 w_13193_29093.n520 16.0005
R5527 w_13193_29093.n558 w_13193_29093.n557 16.0005
R5528 w_13193_29093.n557 w_13193_29093.n556 16.0005
R5529 w_13193_29093.n556 w_13193_29093.n522 16.0005
R5530 w_13193_29093.n551 w_13193_29093.n522 16.0005
R5531 w_13193_29093.n551 w_13193_29093.n550 16.0005
R5532 w_13193_29093.n550 w_13193_29093.n549 16.0005
R5533 w_13193_29093.n581 w_13193_29093.n580 16.0005
R5534 w_13193_29093.n580 w_13193_29093.n516 16.0005
R5535 w_13193_29093.n574 w_13193_29093.n516 16.0005
R5536 w_13193_29093.n574 w_13193_29093.n573 16.0005
R5537 w_13193_29093.n573 w_13193_29093.n572 16.0005
R5538 w_13193_29093.n572 w_13193_29093.n518 16.0005
R5539 w_13193_29093.n566 w_13193_29093.n518 16.0005
R5540 w_13193_29093.n566 w_13193_29093.n565 16.0005
R5541 w_13193_29093.n978 w_13193_29093.n977 16.0005
R5542 w_13193_29093.n977 w_13193_29093.n975 16.0005
R5543 w_13193_29093.n975 w_13193_29093.n972 16.0005
R5544 w_13193_29093.n972 w_13193_29093.n971 16.0005
R5545 w_13193_29093.n971 w_13193_29093.n968 16.0005
R5546 w_13193_29093.n968 w_13193_29093.n967 16.0005
R5547 w_13193_29093.n967 w_13193_29093.n964 16.0005
R5548 w_13193_29093.n964 w_13193_29093.n963 16.0005
R5549 w_13193_29093.n947 w_13193_29093.n944 16.0005
R5550 w_13193_29093.n948 w_13193_29093.n947 16.0005
R5551 w_13193_29093.n951 w_13193_29093.n948 16.0005
R5552 w_13193_29093.n952 w_13193_29093.n951 16.0005
R5553 w_13193_29093.n955 w_13193_29093.n952 16.0005
R5554 w_13193_29093.n956 w_13193_29093.n955 16.0005
R5555 w_13193_29093.n959 w_13193_29093.n956 16.0005
R5556 w_13193_29093.n960 w_13193_29093.n959 16.0005
R5557 w_13193_29093.n928 w_13193_29093.n927 16.0005
R5558 w_13193_29093.n931 w_13193_29093.n928 16.0005
R5559 w_13193_29093.n932 w_13193_29093.n931 16.0005
R5560 w_13193_29093.n935 w_13193_29093.n932 16.0005
R5561 w_13193_29093.n936 w_13193_29093.n935 16.0005
R5562 w_13193_29093.n939 w_13193_29093.n936 16.0005
R5563 w_13193_29093.n940 w_13193_29093.n939 16.0005
R5564 w_13193_29093.n943 w_13193_29093.n940 16.0005
R5565 w_13193_29093.n1411 w_13193_29093.n1406 16.0005
R5566 w_13193_29093.n1412 w_13193_29093.n1411 16.0005
R5567 w_13193_29093.n1413 w_13193_29093.n1412 16.0005
R5568 w_13193_29093.n1413 w_13193_29093.n1403 16.0005
R5569 w_13193_29093.n1419 w_13193_29093.n1403 16.0005
R5570 w_13193_29093.n1420 w_13193_29093.n1419 16.0005
R5571 w_13193_29093.n1421 w_13193_29093.n1420 16.0005
R5572 w_13193_29093.n1421 w_13193_29093.n1400 16.0005
R5573 w_13193_29093.n1441 w_13193_29093.n1395 16.0005
R5574 w_13193_29093.n1435 w_13193_29093.n1395 16.0005
R5575 w_13193_29093.n1435 w_13193_29093.n1434 16.0005
R5576 w_13193_29093.n1434 w_13193_29093.n1433 16.0005
R5577 w_13193_29093.n1433 w_13193_29093.n1397 16.0005
R5578 w_13193_29093.n1428 w_13193_29093.n1397 16.0005
R5579 w_13193_29093.n1428 w_13193_29093.n1427 16.0005
R5580 w_13193_29093.n1427 w_13193_29093.n1426 16.0005
R5581 w_13193_29093.n1457 w_13193_29093.n1456 16.0005
R5582 w_13193_29093.n1456 w_13193_29093.n1391 16.0005
R5583 w_13193_29093.n1451 w_13193_29093.n1391 16.0005
R5584 w_13193_29093.n1451 w_13193_29093.n1450 16.0005
R5585 w_13193_29093.n1450 w_13193_29093.n1449 16.0005
R5586 w_13193_29093.n1449 w_13193_29093.n1393 16.0005
R5587 w_13193_29093.n1443 w_13193_29093.n1393 16.0005
R5588 w_13193_29093.n1443 w_13193_29093.n1442 16.0005
R5589 w_13193_29093.n815 w_13193_29093.n784 16.0005
R5590 w_13193_29093.n816 w_13193_29093.n815 16.0005
R5591 w_13193_29093.n819 w_13193_29093.n816 16.0005
R5592 w_13193_29093.n820 w_13193_29093.n819 16.0005
R5593 w_13193_29093.n823 w_13193_29093.n820 16.0005
R5594 w_13193_29093.n824 w_13193_29093.n823 16.0005
R5595 w_13193_29093.n827 w_13193_29093.n824 16.0005
R5596 w_13193_29093.n828 w_13193_29093.n827 16.0005
R5597 w_13193_29093.n847 w_13193_29093.n844 16.0005
R5598 w_13193_29093.n844 w_13193_29093.n843 16.0005
R5599 w_13193_29093.n843 w_13193_29093.n840 16.0005
R5600 w_13193_29093.n840 w_13193_29093.n839 16.0005
R5601 w_13193_29093.n839 w_13193_29093.n836 16.0005
R5602 w_13193_29093.n836 w_13193_29093.n835 16.0005
R5603 w_13193_29093.n835 w_13193_29093.n832 16.0005
R5604 w_13193_29093.n832 w_13193_29093.n831 16.0005
R5605 w_13193_29093.n864 w_13193_29093.n863 16.0005
R5606 w_13193_29093.n863 w_13193_29093.n860 16.0005
R5607 w_13193_29093.n860 w_13193_29093.n859 16.0005
R5608 w_13193_29093.n859 w_13193_29093.n856 16.0005
R5609 w_13193_29093.n856 w_13193_29093.n855 16.0005
R5610 w_13193_29093.n855 w_13193_29093.n852 16.0005
R5611 w_13193_29093.n852 w_13193_29093.n851 16.0005
R5612 w_13193_29093.n851 w_13193_29093.n848 16.0005
R5613 w_13193_29093.n715 w_13193_29093.n714 16.0005
R5614 w_13193_29093.n714 w_13193_29093.n712 16.0005
R5615 w_13193_29093.n712 w_13193_29093.n709 16.0005
R5616 w_13193_29093.n709 w_13193_29093.n708 16.0005
R5617 w_13193_29093.n708 w_13193_29093.n705 16.0005
R5618 w_13193_29093.n705 w_13193_29093.n704 16.0005
R5619 w_13193_29093.n704 w_13193_29093.n701 16.0005
R5620 w_13193_29093.n701 w_13193_29093.n700 16.0005
R5621 w_13193_29093.n684 w_13193_29093.n681 16.0005
R5622 w_13193_29093.n685 w_13193_29093.n684 16.0005
R5623 w_13193_29093.n688 w_13193_29093.n685 16.0005
R5624 w_13193_29093.n689 w_13193_29093.n688 16.0005
R5625 w_13193_29093.n692 w_13193_29093.n689 16.0005
R5626 w_13193_29093.n693 w_13193_29093.n692 16.0005
R5627 w_13193_29093.n696 w_13193_29093.n693 16.0005
R5628 w_13193_29093.n697 w_13193_29093.n696 16.0005
R5629 w_13193_29093.n665 w_13193_29093.n664 16.0005
R5630 w_13193_29093.n668 w_13193_29093.n665 16.0005
R5631 w_13193_29093.n669 w_13193_29093.n668 16.0005
R5632 w_13193_29093.n672 w_13193_29093.n669 16.0005
R5633 w_13193_29093.n673 w_13193_29093.n672 16.0005
R5634 w_13193_29093.n676 w_13193_29093.n673 16.0005
R5635 w_13193_29093.n677 w_13193_29093.n676 16.0005
R5636 w_13193_29093.n680 w_13193_29093.n677 16.0005
R5637 w_13193_29093.n1330 w_13193_29093.n1217 16.0005
R5638 w_13193_29093.n1250 w_13193_29093.n1217 16.0005
R5639 w_13193_29093.n1251 w_13193_29093.n1250 16.0005
R5640 w_13193_29093.n1251 w_13193_29093.n1247 16.0005
R5641 w_13193_29093.n1257 w_13193_29093.n1247 16.0005
R5642 w_13193_29093.n1258 w_13193_29093.n1257 16.0005
R5643 w_13193_29093.n1259 w_13193_29093.n1258 16.0005
R5644 w_13193_29093.n1259 w_13193_29093.n1244 16.0005
R5645 w_13193_29093.n1279 w_13193_29093.n1239 16.0005
R5646 w_13193_29093.n1273 w_13193_29093.n1239 16.0005
R5647 w_13193_29093.n1273 w_13193_29093.n1272 16.0005
R5648 w_13193_29093.n1272 w_13193_29093.n1271 16.0005
R5649 w_13193_29093.n1271 w_13193_29093.n1241 16.0005
R5650 w_13193_29093.n1266 w_13193_29093.n1241 16.0005
R5651 w_13193_29093.n1266 w_13193_29093.n1265 16.0005
R5652 w_13193_29093.n1265 w_13193_29093.n1264 16.0005
R5653 w_13193_29093.n1295 w_13193_29093.n1294 16.0005
R5654 w_13193_29093.n1294 w_13193_29093.n1235 16.0005
R5655 w_13193_29093.n1289 w_13193_29093.n1235 16.0005
R5656 w_13193_29093.n1289 w_13193_29093.n1288 16.0005
R5657 w_13193_29093.n1288 w_13193_29093.n1287 16.0005
R5658 w_13193_29093.n1287 w_13193_29093.n1237 16.0005
R5659 w_13193_29093.n1281 w_13193_29093.n1237 16.0005
R5660 w_13193_29093.n1281 w_13193_29093.n1280 16.0005
R5661 w_13193_29093.n2381 w_13193_29093.n2380 15.6449
R5662 w_13193_29093.n2524 w_13193_29093.n2523 15.6449
R5663 w_13193_29093.n2213 w_13193_29093.n34 15.567
R5664 w_13193_29093.n2202 w_13193_29093.n31 15.4471
R5665 w_13193_29093.n2467 w_13193_29093.n2466 15.3497
R5666 w_13193_29093.n218 w_13193_29093.t57 15.0005
R5667 w_13193_29093.n218 w_13193_29093.t18 15.0005
R5668 w_13193_29093.n215 w_13193_29093.t221 15.0005
R5669 w_13193_29093.n215 w_13193_29093.t68 15.0005
R5670 w_13193_29093.n2512 w_13193_29093.t73 15.0005
R5671 w_13193_29093.n2512 w_13193_29093.t36 15.0005
R5672 w_13193_29093.n2520 w_13193_29093.t159 15.0005
R5673 w_13193_29093.n2520 w_13193_29093.t80 15.0005
R5674 w_13193_29093.n237 w_13193_29093.t117 15.0005
R5675 w_13193_29093.n237 w_13193_29093.t102 15.0005
R5676 w_13193_29093.n240 w_13193_29093.t89 15.0005
R5677 w_13193_29093.n240 w_13193_29093.t1 15.0005
R5678 w_13193_29093.n2380 w_13193_29093.n241 14.4005
R5679 w_13193_29093.n2719 w_13193_29093.n2718 14.0805
R5680 w_13193_29093.n2724 w_13193_29093.n2723 14.0805
R5681 w_13193_29093.n2328 w_13193_29093.n2327 13.0271
R5682 w_13193_29093.n2507 w_13193_29093.n213 12.8005
R5683 w_13193_29093.n2521 w_13193_29093.n2519 12.8005
R5684 w_13193_29093.n2477 w_13193_29093.n2476 12.8005
R5685 w_13193_29093.n2470 w_13193_29093.n2469 12.8005
R5686 w_13193_29093.n107 w_13193_29093.n106 12.8005
R5687 w_13193_29093.n126 w_13193_29093.n124 12.8005
R5688 w_13193_29093.n2679 w_13193_29093.n2678 12.8005
R5689 w_13193_29093.n2665 w_13193_29093.n2664 12.8005
R5690 w_13193_29093.n2650 w_13193_29093.n2649 12.8005
R5691 w_13193_29093.n2627 w_13193_29093.n164 12.8005
R5692 w_13193_29093.n2608 w_13193_29093.n177 12.8005
R5693 w_13193_29093.n2589 w_13193_29093.n189 12.8005
R5694 w_13193_29093.n2565 w_13193_29093.n2564 12.8005
R5695 w_13193_29093.n2572 w_13193_29093.n193 12.8005
R5696 w_13193_29093.n2292 w_13193_29093.n2291 12.8005
R5697 w_13193_29093.n1095 w_13193_29093.n1094 12.8005
R5698 w_13193_29093.n1094 w_13193_29093.n748 12.8005
R5699 w_13193_29093.n1082 w_13193_29093.n779 12.8005
R5700 w_13193_29093.n1082 w_13193_29093.n1081 12.8005
R5701 w_13193_29093.n2205 w_13193_29093.n2199 12.8005
R5702 w_13193_29093.n2205 w_13193_29093.n2204 12.8005
R5703 w_13193_29093.n2327 w_13193_29093.n2326 11.9273
R5704 w_13193_29093.t118 w_13193_29093.n2434 11.8924
R5705 w_13193_29093.n2696 w_13193_29093.t15 11.8924
R5706 w_13193_29093.t43 w_13193_29093.n2695 11.8924
R5707 w_13193_29093.n1957 w_13193_29093.n1954 11.6369
R5708 w_13193_29093.n1954 w_13193_29093.n1953 11.6369
R5709 w_13193_29093.n1953 w_13193_29093.n1950 11.6369
R5710 w_13193_29093.n1950 w_13193_29093.n1949 11.6369
R5711 w_13193_29093.n1949 w_13193_29093.n1946 11.6369
R5712 w_13193_29093.n1946 w_13193_29093.n1945 11.6369
R5713 w_13193_29093.n1945 w_13193_29093.n1942 11.6369
R5714 w_13193_29093.n1942 w_13193_29093.n283 11.6369
R5715 w_13193_29093.n2156 w_13193_29093.n283 11.6369
R5716 w_13193_29093.n2157 w_13193_29093.n2156 11.6369
R5717 w_13193_29093.n2158 w_13193_29093.n281 11.6369
R5718 w_13193_29093.n2164 w_13193_29093.n281 11.6369
R5719 w_13193_29093.n2165 w_13193_29093.n2164 11.6369
R5720 w_13193_29093.n2166 w_13193_29093.n2165 11.6369
R5721 w_13193_29093.n2166 w_13193_29093.n279 11.6369
R5722 w_13193_29093.n2172 w_13193_29093.n279 11.6369
R5723 w_13193_29093.n2173 w_13193_29093.n2172 11.6369
R5724 w_13193_29093.n2174 w_13193_29093.n2173 11.6369
R5725 w_13193_29093.n2174 w_13193_29093.n277 11.6369
R5726 w_13193_29093.n2179 w_13193_29093.n277 11.6369
R5727 w_13193_29093.n2180 w_13193_29093.n2179 11.6369
R5728 w_13193_29093.n1711 w_13193_29093.n1708 11.6369
R5729 w_13193_29093.n1708 w_13193_29093.n1707 11.6369
R5730 w_13193_29093.n1707 w_13193_29093.n1704 11.6369
R5731 w_13193_29093.n1704 w_13193_29093.n1703 11.6369
R5732 w_13193_29093.n1703 w_13193_29093.n1700 11.6369
R5733 w_13193_29093.n1700 w_13193_29093.n1699 11.6369
R5734 w_13193_29093.n1699 w_13193_29093.n1696 11.6369
R5735 w_13193_29093.n1696 w_13193_29093.n423 11.6369
R5736 w_13193_29093.n1779 w_13193_29093.n423 11.6369
R5737 w_13193_29093.n1780 w_13193_29093.n1779 11.6369
R5738 w_13193_29093.n1802 w_13193_29093.n414 11.6369
R5739 w_13193_29093.n415 w_13193_29093.n414 11.6369
R5740 w_13193_29093.n1795 w_13193_29093.n415 11.6369
R5741 w_13193_29093.n1795 w_13193_29093.n1794 11.6369
R5742 w_13193_29093.n1794 w_13193_29093.n1793 11.6369
R5743 w_13193_29093.n1793 w_13193_29093.n417 11.6369
R5744 w_13193_29093.n1788 w_13193_29093.n417 11.6369
R5745 w_13193_29093.n1788 w_13193_29093.n1787 11.6369
R5746 w_13193_29093.n1787 w_13193_29093.n1786 11.6369
R5747 w_13193_29093.n1786 w_13193_29093.n420 11.6369
R5748 w_13193_29093.n1781 w_13193_29093.n420 11.6369
R5749 w_13193_29093.n1772 w_13193_29093.n1769 11.6369
R5750 w_13193_29093.n1769 w_13193_29093.n1768 11.6369
R5751 w_13193_29093.n1768 w_13193_29093.n1765 11.6369
R5752 w_13193_29093.n1765 w_13193_29093.n1764 11.6369
R5753 w_13193_29093.n1764 w_13193_29093.n1761 11.6369
R5754 w_13193_29093.n1761 w_13193_29093.n1760 11.6369
R5755 w_13193_29093.n1760 w_13193_29093.n1757 11.6369
R5756 w_13193_29093.n1757 w_13193_29093.n1756 11.6369
R5757 w_13193_29093.n1756 w_13193_29093.n1753 11.6369
R5758 w_13193_29093.n1753 w_13193_29093.n1752 11.6369
R5759 w_13193_29093.n1169 w_13193_29093.n1166 11.6369
R5760 w_13193_29093.n1170 w_13193_29093.n1169 11.6369
R5761 w_13193_29093.n1173 w_13193_29093.n1170 11.6369
R5762 w_13193_29093.n1174 w_13193_29093.n1173 11.6369
R5763 w_13193_29093.n1177 w_13193_29093.n1174 11.6369
R5764 w_13193_29093.n1178 w_13193_29093.n1177 11.6369
R5765 w_13193_29093.n1181 w_13193_29093.n1178 11.6369
R5766 w_13193_29093.n1182 w_13193_29093.n1181 11.6369
R5767 w_13193_29093.n1185 w_13193_29093.n1182 11.6369
R5768 w_13193_29093.n1186 w_13193_29093.n1185 11.6369
R5769 w_13193_29093.n1191 w_13193_29093.n1190 11.6369
R5770 w_13193_29093.n1192 w_13193_29093.n1191 11.6369
R5771 w_13193_29093.n1192 w_13193_29093.n629 11.6369
R5772 w_13193_29093.n1198 w_13193_29093.n629 11.6369
R5773 w_13193_29093.n1199 w_13193_29093.n1198 11.6369
R5774 w_13193_29093.n1200 w_13193_29093.n1199 11.6369
R5775 w_13193_29093.n1200 w_13193_29093.n627 11.6369
R5776 w_13193_29093.n1206 w_13193_29093.n627 11.6369
R5777 w_13193_29093.n1207 w_13193_29093.n1206 11.6369
R5778 w_13193_29093.n1208 w_13193_29093.n1207 11.6369
R5779 w_13193_29093.n1208 w_13193_29093.n623 11.6369
R5780 w_13193_29093.n1384 w_13193_29093.n610 11.6369
R5781 w_13193_29093.n1467 w_13193_29093.n610 11.6369
R5782 w_13193_29093.n1468 w_13193_29093.n1467 11.6369
R5783 w_13193_29093.n1472 w_13193_29093.n1468 11.6369
R5784 w_13193_29093.n1472 w_13193_29093.n1471 11.6369
R5785 w_13193_29093.n1471 w_13193_29093.n1470 11.6369
R5786 w_13193_29093.n1470 w_13193_29093.n592 11.6369
R5787 w_13193_29093.n1491 w_13193_29093.n592 11.6369
R5788 w_13193_29093.n1492 w_13193_29093.n1491 11.6369
R5789 w_13193_29093.n1494 w_13193_29093.n1492 11.6369
R5790 w_13193_29093.n1494 w_13193_29093.n1493 11.6369
R5791 w_13193_29093.n1587 w_13193_29093.n1586 11.6369
R5792 w_13193_29093.n1586 w_13193_29093.n1585 11.6369
R5793 w_13193_29093.n1585 w_13193_29093.n496 11.6369
R5794 w_13193_29093.n1579 w_13193_29093.n496 11.6369
R5795 w_13193_29093.n1579 w_13193_29093.n1578 11.6369
R5796 w_13193_29093.n1578 w_13193_29093.n1577 11.6369
R5797 w_13193_29093.n1577 w_13193_29093.n502 11.6369
R5798 w_13193_29093.n504 w_13193_29093.n502 11.6369
R5799 w_13193_29093.n504 w_13193_29093.n503 11.6369
R5800 w_13193_29093.n503 w_13193_29093.n448 11.6369
R5801 w_13193_29093.n448 w_13193_29093.n446 11.6369
R5802 w_13193_29093.n1741 w_13193_29093.n1739 11.6369
R5803 w_13193_29093.n1739 w_13193_29093.n1736 11.6369
R5804 w_13193_29093.n1736 w_13193_29093.n1735 11.6369
R5805 w_13193_29093.n1735 w_13193_29093.n1732 11.6369
R5806 w_13193_29093.n1732 w_13193_29093.n1731 11.6369
R5807 w_13193_29093.n1731 w_13193_29093.n1728 11.6369
R5808 w_13193_29093.n1728 w_13193_29093.n1727 11.6369
R5809 w_13193_29093.n1727 w_13193_29093.n1724 11.6369
R5810 w_13193_29093.n1724 w_13193_29093.n1723 11.6369
R5811 w_13193_29093.n1723 w_13193_29093.n1721 11.6369
R5812 w_13193_29093.n1658 w_13193_29093.n384 11.6369
R5813 w_13193_29093.n1660 w_13193_29093.n1658 11.6369
R5814 w_13193_29093.n1660 w_13193_29093.n1659 11.6369
R5815 w_13193_29093.n1659 w_13193_29093.n472 11.6369
R5816 w_13193_29093.n472 w_13193_29093.n470 11.6369
R5817 w_13193_29093.n1679 w_13193_29093.n470 11.6369
R5818 w_13193_29093.n1680 w_13193_29093.n1679 11.6369
R5819 w_13193_29093.n1682 w_13193_29093.n1680 11.6369
R5820 w_13193_29093.n1682 w_13193_29093.n1681 11.6369
R5821 w_13193_29093.n1681 w_13193_29093.n455 11.6369
R5822 w_13193_29093.n1720 w_13193_29093.n455 11.6369
R5823 w_13193_29093.n2150 w_13193_29093.n2149 11.6369
R5824 w_13193_29093.n2149 w_13193_29093.n2146 11.6369
R5825 w_13193_29093.n2146 w_13193_29093.n2145 11.6369
R5826 w_13193_29093.n2145 w_13193_29093.n2142 11.6369
R5827 w_13193_29093.n2142 w_13193_29093.n2141 11.6369
R5828 w_13193_29093.n2141 w_13193_29093.n2138 11.6369
R5829 w_13193_29093.n2138 w_13193_29093.n2137 11.6369
R5830 w_13193_29093.n2137 w_13193_29093.n2134 11.6369
R5831 w_13193_29093.n2134 w_13193_29093.n2133 11.6369
R5832 w_13193_29093.n2133 w_13193_29093.n2131 11.6369
R5833 w_13193_29093.n2130 w_13193_29093.n307 11.6369
R5834 w_13193_29093.n308 w_13193_29093.n307 11.6369
R5835 w_13193_29093.n2123 w_13193_29093.n308 11.6369
R5836 w_13193_29093.n2123 w_13193_29093.n2122 11.6369
R5837 w_13193_29093.n2122 w_13193_29093.n2121 11.6369
R5838 w_13193_29093.n2121 w_13193_29093.n310 11.6369
R5839 w_13193_29093.n2116 w_13193_29093.n310 11.6369
R5840 w_13193_29093.n2116 w_13193_29093.n2115 11.6369
R5841 w_13193_29093.n2115 w_13193_29093.n2114 11.6369
R5842 w_13193_29093.n2114 w_13193_29093.n313 11.6369
R5843 w_13193_29093.n2109 w_13193_29093.n313 11.6369
R5844 w_13193_29093.n1917 w_13193_29093.n316 11.6369
R5845 w_13193_29093.n1917 w_13193_29093.n1916 11.6369
R5846 w_13193_29093.n1916 w_13193_29093.n1915 11.6369
R5847 w_13193_29093.n1915 w_13193_29093.n324 11.6369
R5848 w_13193_29093.n360 w_13193_29093.n324 11.6369
R5849 w_13193_29093.n361 w_13193_29093.n360 11.6369
R5850 w_13193_29093.n361 w_13193_29093.n358 11.6369
R5851 w_13193_29093.n381 w_13193_29093.n358 11.6369
R5852 w_13193_29093.n382 w_13193_29093.n381 11.6369
R5853 w_13193_29093.n1840 w_13193_29093.n382 11.6369
R5854 w_13193_29093.n1840 w_13193_29093.n1839 11.6369
R5855 w_13193_29093.n2188 w_13193_29093.n271 11.6369
R5856 w_13193_29093.n2189 w_13193_29093.n2188 11.6369
R5857 w_13193_29093.n2190 w_13193_29093.n2189 11.6369
R5858 w_13193_29093.n2190 w_13193_29093.n269 11.6369
R5859 w_13193_29093.n269 w_13193_29093.n266 11.6369
R5860 w_13193_29093.n2197 w_13193_29093.n267 11.6369
R5861 w_13193_29093.n1807 w_13193_29093.n267 11.6369
R5862 w_13193_29093.n1807 w_13193_29093.n1806 11.6369
R5863 w_13193_29093.n1812 w_13193_29093.n1806 11.6369
R5864 w_13193_29093.n1813 w_13193_29093.n1812 11.6369
R5865 w_13193_29093.t215 w_13193_29093.n1024 10.1221
R5866 w_13193_29093.n987 w_13193_29093.t2 10.1221
R5867 w_13193_29093.n998 w_13193_29093.t210 10.1221
R5868 w_13193_29093.n1010 w_13193_29093.t211 10.1221
R5869 w_13193_29093.n2701 w_13193_29093.t166 9.88814
R5870 w_13193_29093.n2691 w_13193_29093.n69 9.6005
R5871 w_13193_29093.n2691 w_13193_29093.n2690 9.6005
R5872 w_13193_29093.n2427 w_13193_29093.n2426 9.6005
R5873 w_13193_29093.n2426 w_13193_29093.n2425 9.6005
R5874 w_13193_29093.n246 w_13193_29093.t259 9.6005
R5875 w_13193_29093.n251 w_13193_29093.t266 9.6005
R5876 w_13193_29093.n762 w_13193_29093.t268 9.6005
R5877 w_13193_29093.n755 w_13193_29093.t264 9.6005
R5878 w_13193_29093.n2727 w_13193_29093.n57 9.58175
R5879 w_13193_29093.n2759 w_13193_29093.n2758 9.58175
R5880 w_13193_29093.n2465 w_13193_29093.n2464 9.40114
R5881 w_13193_29093.n1095 w_13193_29093.n747 9.36264
R5882 w_13193_29093.n1084 w_13193_29093.n779 9.36264
R5883 w_13193_29093.n2207 w_13193_29093.n2199 9.36264
R5884 w_13193_29093.n2584 w_13193_29093.n2583 9.3005
R5885 w_13193_29093.n2585 w_13193_29093.n190 9.3005
R5886 w_13193_29093.n2587 w_13193_29093.n2586 9.3005
R5887 w_13193_29093.n2588 w_13193_29093.n187 9.3005
R5888 w_13193_29093.n2590 w_13193_29093.n2589 9.3005
R5889 w_13193_29093.n2591 w_13193_29093.n186 9.3005
R5890 w_13193_29093.n2593 w_13193_29093.n2592 9.3005
R5891 w_13193_29093.n2594 w_13193_29093.n184 9.3005
R5892 w_13193_29093.n2595 w_13193_29093.n182 9.3005
R5893 w_13193_29093.n2597 w_13193_29093.n2596 9.3005
R5894 w_13193_29093.n2598 w_13193_29093.n181 9.3005
R5895 w_13193_29093.n2600 w_13193_29093.n2599 9.3005
R5896 w_13193_29093.n2601 w_13193_29093.n179 9.3005
R5897 w_13193_29093.n2603 w_13193_29093.n2602 9.3005
R5898 w_13193_29093.n2604 w_13193_29093.n178 9.3005
R5899 w_13193_29093.n2606 w_13193_29093.n2605 9.3005
R5900 w_13193_29093.n2607 w_13193_29093.n175 9.3005
R5901 w_13193_29093.n2609 w_13193_29093.n2608 9.3005
R5902 w_13193_29093.n2610 w_13193_29093.n174 9.3005
R5903 w_13193_29093.n2612 w_13193_29093.n2611 9.3005
R5904 w_13193_29093.n2613 w_13193_29093.n172 9.3005
R5905 w_13193_29093.n2614 w_13193_29093.n170 9.3005
R5906 w_13193_29093.n2616 w_13193_29093.n2615 9.3005
R5907 w_13193_29093.n2617 w_13193_29093.n169 9.3005
R5908 w_13193_29093.n2619 w_13193_29093.n2618 9.3005
R5909 w_13193_29093.n2620 w_13193_29093.n167 9.3005
R5910 w_13193_29093.n2622 w_13193_29093.n2621 9.3005
R5911 w_13193_29093.n2623 w_13193_29093.n166 9.3005
R5912 w_13193_29093.n2625 w_13193_29093.n2624 9.3005
R5913 w_13193_29093.n2626 w_13193_29093.n165 9.3005
R5914 w_13193_29093.n2628 w_13193_29093.n2627 9.3005
R5915 w_13193_29093.n2630 w_13193_29093.n2629 9.3005
R5916 w_13193_29093.n2631 w_13193_29093.n161 9.3005
R5917 w_13193_29093.n2633 w_13193_29093.n2632 9.3005
R5918 w_13193_29093.n2634 w_13193_29093.n160 9.3005
R5919 w_13193_29093.n2636 w_13193_29093.n2635 9.3005
R5920 w_13193_29093.n2638 w_13193_29093.n158 9.3005
R5921 w_13193_29093.n2640 w_13193_29093.n2639 9.3005
R5922 w_13193_29093.n2641 w_13193_29093.n157 9.3005
R5923 w_13193_29093.n2643 w_13193_29093.n2642 9.3005
R5924 w_13193_29093.n2644 w_13193_29093.n155 9.3005
R5925 w_13193_29093.n2646 w_13193_29093.n2645 9.3005
R5926 w_13193_29093.n2647 w_13193_29093.n154 9.3005
R5927 w_13193_29093.n2649 w_13193_29093.n2648 9.3005
R5928 w_13193_29093.n2651 w_13193_29093.n152 9.3005
R5929 w_13193_29093.n2653 w_13193_29093.n2652 9.3005
R5930 w_13193_29093.n2654 w_13193_29093.n151 9.3005
R5931 w_13193_29093.n2656 w_13193_29093.n2655 9.3005
R5932 w_13193_29093.n2657 w_13193_29093.n149 9.3005
R5933 w_13193_29093.n2659 w_13193_29093.n2658 9.3005
R5934 w_13193_29093.n2660 w_13193_29093.n148 9.3005
R5935 w_13193_29093.n2662 w_13193_29093.n2661 9.3005
R5936 w_13193_29093.n2663 w_13193_29093.n146 9.3005
R5937 w_13193_29093.n2666 w_13193_29093.n2665 9.3005
R5938 w_13193_29093.n2667 w_13193_29093.n145 9.3005
R5939 w_13193_29093.n2669 w_13193_29093.n2668 9.3005
R5940 w_13193_29093.n2671 w_13193_29093.n143 9.3005
R5941 w_13193_29093.n2673 w_13193_29093.n2672 9.3005
R5942 w_13193_29093.n2674 w_13193_29093.n142 9.3005
R5943 w_13193_29093.n2676 w_13193_29093.n2675 9.3005
R5944 w_13193_29093.n2677 w_13193_29093.n140 9.3005
R5945 w_13193_29093.n2680 w_13193_29093.n2679 9.3005
R5946 w_13193_29093.n2681 w_13193_29093.n139 9.3005
R5947 w_13193_29093.n2683 w_13193_29093.n2682 9.3005
R5948 w_13193_29093.n2684 w_13193_29093.n138 9.3005
R5949 w_13193_29093.n2685 w_13193_29093.n137 9.3005
R5950 w_13193_29093.n2687 w_13193_29093.n2686 9.3005
R5951 w_13193_29093.n2688 w_13193_29093.n70 9.3005
R5952 w_13193_29093.n2690 w_13193_29093.n2689 9.3005
R5953 w_13193_29093.n136 w_13193_29093.n69 9.3005
R5954 w_13193_29093.n135 w_13193_29093.n134 9.3005
R5955 w_13193_29093.n133 w_13193_29093.n71 9.3005
R5956 w_13193_29093.n132 w_13193_29093.n131 9.3005
R5957 w_13193_29093.n130 w_13193_29093.n73 9.3005
R5958 w_13193_29093.n129 w_13193_29093.n128 9.3005
R5959 w_13193_29093.n127 w_13193_29093.n74 9.3005
R5960 w_13193_29093.n124 w_13193_29093.n123 9.3005
R5961 w_13193_29093.n122 w_13193_29093.n75 9.3005
R5962 w_13193_29093.n121 w_13193_29093.n120 9.3005
R5963 w_13193_29093.n119 w_13193_29093.n76 9.3005
R5964 w_13193_29093.n118 w_13193_29093.n117 9.3005
R5965 w_13193_29093.n116 w_13193_29093.n77 9.3005
R5966 w_13193_29093.n115 w_13193_29093.n114 9.3005
R5967 w_13193_29093.n112 w_13193_29093.n78 9.3005
R5968 w_13193_29093.n111 w_13193_29093.n110 9.3005
R5969 w_13193_29093.n109 w_13193_29093.n79 9.3005
R5970 w_13193_29093.n108 w_13193_29093.n107 9.3005
R5971 w_13193_29093.n104 w_13193_29093.n80 9.3005
R5972 w_13193_29093.n103 w_13193_29093.n102 9.3005
R5973 w_13193_29093.n101 w_13193_29093.n82 9.3005
R5974 w_13193_29093.n100 w_13193_29093.n99 9.3005
R5975 w_13193_29093.n98 w_13193_29093.n83 9.3005
R5976 w_13193_29093.n97 w_13193_29093.n96 9.3005
R5977 w_13193_29093.n95 w_13193_29093.n84 9.3005
R5978 w_13193_29093.n94 w_13193_29093.n93 9.3005
R5979 w_13193_29093.n92 w_13193_29093.n85 9.3005
R5980 w_13193_29093.n91 w_13193_29093.n90 9.3005
R5981 w_13193_29093.n2577 w_13193_29093.n191 9.3005
R5982 w_13193_29093.n2576 w_13193_29093.n2575 9.3005
R5983 w_13193_29093.n2574 w_13193_29093.n193 9.3005
R5984 w_13193_29093.n2556 w_13193_29093.n200 9.3005
R5985 w_13193_29093.n2558 w_13193_29093.n2557 9.3005
R5986 w_13193_29093.n2559 w_13193_29093.n199 9.3005
R5987 w_13193_29093.n2561 w_13193_29093.n2560 9.3005
R5988 w_13193_29093.n2562 w_13193_29093.n198 9.3005
R5989 w_13193_29093.n2564 w_13193_29093.n2563 9.3005
R5990 w_13193_29093.n2565 w_13193_29093.n196 9.3005
R5991 w_13193_29093.n2567 w_13193_29093.n2566 9.3005
R5992 w_13193_29093.n2568 w_13193_29093.n195 9.3005
R5993 w_13193_29093.n2570 w_13193_29093.n2569 9.3005
R5994 w_13193_29093.n2571 w_13193_29093.n194 9.3005
R5995 w_13193_29093.n2573 w_13193_29093.n2572 9.3005
R5996 w_13193_29093.n2315 w_13193_29093.n2314 9.3005
R5997 w_13193_29093.n2215 w_13193_29093.n2214 9.3005
R5998 w_13193_29093.n2455 w_13193_29093.n2454 9.3005
R5999 w_13193_29093.n2457 w_13193_29093.n2456 9.3005
R6000 w_13193_29093.n2458 w_13193_29093.n2453 9.3005
R6001 w_13193_29093.n2452 w_13193_29093.n2217 9.3005
R6002 w_13193_29093.n2451 w_13193_29093.n2450 9.3005
R6003 w_13193_29093.n2449 w_13193_29093.n2218 9.3005
R6004 w_13193_29093.n2448 w_13193_29093.n2220 9.3005
R6005 w_13193_29093.n2281 w_13193_29093.n2219 9.3005
R6006 w_13193_29093.n2283 w_13193_29093.n2282 9.3005
R6007 w_13193_29093.n2284 w_13193_29093.n2275 9.3005
R6008 w_13193_29093.n2286 w_13193_29093.n2285 9.3005
R6009 w_13193_29093.n2287 w_13193_29093.n2274 9.3005
R6010 w_13193_29093.n2289 w_13193_29093.n2288 9.3005
R6011 w_13193_29093.n2290 w_13193_29093.n2272 9.3005
R6012 w_13193_29093.n2293 w_13193_29093.n2292 9.3005
R6013 w_13193_29093.n2294 w_13193_29093.n2271 9.3005
R6014 w_13193_29093.n2296 w_13193_29093.n2295 9.3005
R6015 w_13193_29093.n2297 w_13193_29093.n2269 9.3005
R6016 w_13193_29093.n2299 w_13193_29093.n2298 9.3005
R6017 w_13193_29093.n2300 w_13193_29093.n2268 9.3005
R6018 w_13193_29093.n2302 w_13193_29093.n2301 9.3005
R6019 w_13193_29093.n2303 w_13193_29093.n2267 9.3005
R6020 w_13193_29093.n2304 w_13193_29093.n2265 9.3005
R6021 w_13193_29093.n2306 w_13193_29093.n2305 9.3005
R6022 w_13193_29093.n2307 w_13193_29093.n2264 9.3005
R6023 w_13193_29093.n2309 w_13193_29093.n2308 9.3005
R6024 w_13193_29093.n2310 w_13193_29093.n2263 9.3005
R6025 w_13193_29093.n2312 w_13193_29093.n2311 9.3005
R6026 w_13193_29093.n2313 w_13193_29093.n2262 9.3005
R6027 w_13193_29093.n2316 w_13193_29093.n2257 9.3005
R6028 w_13193_29093.n2317 w_13193_29093.n2256 9.3005
R6029 w_13193_29093.n2319 w_13193_29093.n2318 9.3005
R6030 w_13193_29093.n2320 w_13193_29093.n2255 9.3005
R6031 w_13193_29093.n2322 w_13193_29093.n2321 9.3005
R6032 w_13193_29093.n2323 w_13193_29093.n2254 9.3005
R6033 w_13193_29093.n2325 w_13193_29093.n2324 9.3005
R6034 w_13193_29093.n2393 w_13193_29093.n2374 9.3005
R6035 w_13193_29093.n2395 w_13193_29093.n2394 9.3005
R6036 w_13193_29093.n2396 w_13193_29093.n2373 9.3005
R6037 w_13193_29093.n2398 w_13193_29093.n2397 9.3005
R6038 w_13193_29093.n2399 w_13193_29093.n2372 9.3005
R6039 w_13193_29093.n2401 w_13193_29093.n2400 9.3005
R6040 w_13193_29093.n2402 w_13193_29093.n2370 9.3005
R6041 w_13193_29093.n2404 w_13193_29093.n2403 9.3005
R6042 w_13193_29093.n2405 w_13193_29093.n2369 9.3005
R6043 w_13193_29093.n2407 w_13193_29093.n2406 9.3005
R6044 w_13193_29093.n2409 w_13193_29093.n2408 9.3005
R6045 w_13193_29093.n2410 w_13193_29093.n2367 9.3005
R6046 w_13193_29093.n2412 w_13193_29093.n2411 9.3005
R6047 w_13193_29093.n2413 w_13193_29093.n2365 9.3005
R6048 w_13193_29093.n2415 w_13193_29093.n2414 9.3005
R6049 w_13193_29093.n2416 w_13193_29093.n2364 9.3005
R6050 w_13193_29093.n2418 w_13193_29093.n2417 9.3005
R6051 w_13193_29093.n2419 w_13193_29093.n2363 9.3005
R6052 w_13193_29093.n2421 w_13193_29093.n2420 9.3005
R6053 w_13193_29093.n2422 w_13193_29093.n2362 9.3005
R6054 w_13193_29093.n2424 w_13193_29093.n2423 9.3005
R6055 w_13193_29093.n2425 w_13193_29093.n2361 9.3005
R6056 w_13193_29093.n2428 w_13193_29093.n2427 9.3005
R6057 w_13193_29093.n2429 w_13193_29093.n2360 9.3005
R6058 w_13193_29093.n2431 w_13193_29093.n2430 9.3005
R6059 w_13193_29093.n2432 w_13193_29093.n2359 9.3005
R6060 w_13193_29093.n2358 w_13193_29093.n2227 9.3005
R6061 w_13193_29093.n2357 w_13193_29093.n2356 9.3005
R6062 w_13193_29093.n2355 w_13193_29093.n2228 9.3005
R6063 w_13193_29093.n2354 w_13193_29093.n2353 9.3005
R6064 w_13193_29093.n2352 w_13193_29093.n2229 9.3005
R6065 w_13193_29093.n2351 w_13193_29093.n2350 9.3005
R6066 w_13193_29093.n2349 w_13193_29093.n2230 9.3005
R6067 w_13193_29093.n2348 w_13193_29093.n2347 9.3005
R6068 w_13193_29093.n2346 w_13193_29093.n2231 9.3005
R6069 w_13193_29093.n2345 w_13193_29093.n2344 9.3005
R6070 w_13193_29093.n2343 w_13193_29093.n2232 9.3005
R6071 w_13193_29093.n2341 w_13193_29093.n2340 9.3005
R6072 w_13193_29093.n2339 w_13193_29093.n2338 9.3005
R6073 w_13193_29093.n2337 w_13193_29093.n2235 9.3005
R6074 w_13193_29093.n2336 w_13193_29093.n2236 9.3005
R6075 w_13193_29093.n2335 w_13193_29093.n2334 9.3005
R6076 w_13193_29093.n2333 w_13193_29093.n2237 9.3005
R6077 w_13193_29093.n2332 w_13193_29093.n2331 9.3005
R6078 w_13193_29093.n2330 w_13193_29093.n2238 9.3005
R6079 w_13193_29093.n1094 w_13193_29093.n1093 9.3005
R6080 w_13193_29093.n1092 w_13193_29093.n748 9.3005
R6081 w_13193_29093.n1083 w_13193_29093.n1082 9.3005
R6082 w_13193_29093.n1081 w_13193_29093.n778 9.3005
R6083 w_13193_29093.n2206 w_13193_29093.n2205 9.3005
R6084 w_13193_29093.n2204 w_13193_29093.n265 9.3005
R6085 w_13193_29093.n2728 w_13193_29093.n54 9.3005
R6086 w_13193_29093.n2730 w_13193_29093.n2729 9.3005
R6087 w_13193_29093.n2731 w_13193_29093.n53 9.3005
R6088 w_13193_29093.n2733 w_13193_29093.n2732 9.3005
R6089 w_13193_29093.n2734 w_13193_29093.n50 9.3005
R6090 w_13193_29093.n2736 w_13193_29093.n2735 9.3005
R6091 w_13193_29093.n2737 w_13193_29093.n49 9.3005
R6092 w_13193_29093.n2739 w_13193_29093.n2738 9.3005
R6093 w_13193_29093.n2740 w_13193_29093.n46 9.3005
R6094 w_13193_29093.n2742 w_13193_29093.n2741 9.3005
R6095 w_13193_29093.n2743 w_13193_29093.n45 9.3005
R6096 w_13193_29093.n2745 w_13193_29093.n2744 9.3005
R6097 w_13193_29093.n2746 w_13193_29093.n42 9.3005
R6098 w_13193_29093.n2748 w_13193_29093.n2747 9.3005
R6099 w_13193_29093.n2749 w_13193_29093.n39 9.3005
R6100 w_13193_29093.n2751 w_13193_29093.n2750 9.3005
R6101 w_13193_29093.n2752 w_13193_29093.n36 9.3005
R6102 w_13193_29093.n2754 w_13193_29093.n2753 9.3005
R6103 w_13193_29093.n2755 w_13193_29093.n35 9.3005
R6104 w_13193_29093.n2757 w_13193_29093.n2756 9.3005
R6105 w_13193_29093.n2519 w_13193_29093.n210 9.3005
R6106 w_13193_29093.n2518 w_13193_29093.n2517 9.3005
R6107 w_13193_29093.n2516 w_13193_29093.n211 9.3005
R6108 w_13193_29093.n2515 w_13193_29093.n2514 9.3005
R6109 w_13193_29093.n2513 w_13193_29093.n212 9.3005
R6110 w_13193_29093.n2511 w_13193_29093.n2510 9.3005
R6111 w_13193_29093.n2509 w_13193_29093.n213 9.3005
R6112 w_13193_29093.n2508 w_13193_29093.n2507 9.3005
R6113 w_13193_29093.n2495 w_13193_29093.n214 9.3005
R6114 w_13193_29093.n2494 w_13193_29093.n2493 9.3005
R6115 w_13193_29093.n2492 w_13193_29093.n216 9.3005
R6116 w_13193_29093.n2491 w_13193_29093.n2490 9.3005
R6117 w_13193_29093.n2489 w_13193_29093.n217 9.3005
R6118 w_13193_29093.n2488 w_13193_29093.n2487 9.3005
R6119 w_13193_29093.n2486 w_13193_29093.n219 9.3005
R6120 w_13193_29093.n2485 w_13193_29093.n2484 9.3005
R6121 w_13193_29093.n2483 w_13193_29093.n220 9.3005
R6122 w_13193_29093.n2482 w_13193_29093.n2481 9.3005
R6123 w_13193_29093.n2480 w_13193_29093.n234 9.3005
R6124 w_13193_29093.n2479 w_13193_29093.n2478 9.3005
R6125 w_13193_29093.n2477 w_13193_29093.n235 9.3005
R6126 w_13193_29093.n2476 w_13193_29093.n236 9.3005
R6127 w_13193_29093.n2475 w_13193_29093.n2474 9.3005
R6128 w_13193_29093.n2473 w_13193_29093.n238 9.3005
R6129 w_13193_29093.n2472 w_13193_29093.n2471 9.3005
R6130 w_13193_29093.n2470 w_13193_29093.n239 9.3005
R6131 w_13193_29093.n2469 w_13193_29093.n2468 9.3005
R6132 w_13193_29093.n2440 w_13193_29093.n2439 9.21941
R6133 w_13193_29093.t53 w_13193_29093.t278 8.67615
R6134 w_13193_29093.n2392 w_13193_29093.n192 8.31939
R6135 w_13193_29093.t53 w_13193_29093.n31 7.77365
R6136 w_13193_29093.n2392 w_13193_29093.n2391 7.56834
R6137 w_13193_29093.n2582 w_13193_29093.n2580 7.37605
R6138 w_13193_29093.n2464 w_13193_29093.n2463 7.22808
R6139 w_13193_29093.n2383 w_13193_29093.n2379 7.11161
R6140 w_13193_29093.n2526 w_13193_29093.n209 7.11161
R6141 w_13193_29093.n89 w_13193_29093.n87 7.07105
R6142 w_13193_29093.n2329 w_13193_29093.n2328 6.86155
R6143 w_13193_29093.n2326 w_13193_29093.n2253 6.86155
R6144 w_13193_29093.n2555 w_13193_29093.n2554 6.86152
R6145 w_13193_29093.n1803 w_13193_29093.n1802 6.72373
R6146 w_13193_29093.n1384 w_13193_29093.n1383 6.72373
R6147 w_13193_29093.n1587 w_13193_29093.n495 6.72373
R6148 w_13193_29093.n1838 w_13193_29093.n384 6.72373
R6149 w_13193_29093.n2108 w_13193_29093.n316 6.72373
R6150 w_13193_29093.n274 w_13193_29093.n271 6.72373
R6151 w_13193_29093.n2522 w_13193_29093.n2521 6.69883
R6152 w_13193_29093.n2482 w_13193_29093.n234 6.4005
R6153 w_13193_29093.n2484 w_13193_29093.n219 6.4005
R6154 w_13193_29093.n2514 w_13193_29093.n2513 6.4005
R6155 w_13193_29093.n106 w_13193_29093.n104 6.4005
R6156 w_13193_29093.n127 w_13193_29093.n126 6.4005
R6157 w_13193_29093.n2678 w_13193_29093.n2677 6.4005
R6158 w_13193_29093.n2664 w_13193_29093.n2663 6.4005
R6159 w_13193_29093.n2651 w_13193_29093.n2650 6.4005
R6160 w_13193_29093.n2630 w_13193_29093.n164 6.4005
R6161 w_13193_29093.n177 w_13193_29093.n174 6.4005
R6162 w_13193_29093.n189 w_13193_29093.n186 6.4005
R6163 w_13193_29093.n2291 w_13193_29093.n2290 6.4005
R6164 w_13193_29093.n2707 w_13193_29093.n2706 6.4005
R6165 w_13193_29093.n2715 w_13193_29093.n2714 6.4005
R6166 w_13193_29093.n2211 w_13193_29093.n263 6.36829
R6167 w_13193_29093.n2180 w_13193_29093.n274 6.20656
R6168 w_13193_29093.n1383 w_13193_29093.n623 6.20656
R6169 w_13193_29093.n1493 w_13193_29093.n495 6.20656
R6170 w_13193_29093.n2109 w_13193_29093.n2108 6.20656
R6171 w_13193_29093.n1839 w_13193_29093.n1838 6.20656
R6172 w_13193_29093.n1813 w_13193_29093.n1803 6.20656
R6173 w_13193_29093.n2198 w_13193_29093.n2197 6.07727
R6174 w_13193_29093.n257 w_13193_29093.n242 5.81868
R6175 w_13193_29093.n2467 w_13193_29093.n241 5.80512
R6176 w_13193_29093.n2342 w_13193_29093.n2225 5.68939
R6177 w_13193_29093.n2260 w_13193_29093.n2258 5.68939
R6178 w_13193_29093.n2261 w_13193_29093.n2260 5.68939
R6179 w_13193_29093.n2211 w_13193_29093.n2210 5.6447
R6180 w_13193_29093.n2198 w_13193_29093.n266 5.5601
R6181 w_13193_29093.n1652 w_13193_29093.n1651 5.51161
R6182 w_13193_29093.n1897 w_13193_29093.n319 5.51161
R6183 w_13193_29093.n2023 w_13193_29093.n1962 5.51161
R6184 w_13193_29093.n1546 w_13193_29093.n581 5.51161
R6185 w_13193_29093.n927 w_13193_29093.n904 5.51161
R6186 w_13193_29093.n1457 w_13193_29093.n1390 5.51161
R6187 w_13193_29093.n864 w_13193_29093.n742 5.51161
R6188 w_13193_29093.n664 w_13193_29093.n632 5.51161
R6189 w_13193_29093.n1295 w_13193_29093.n1234 5.51161
R6190 w_13193_29093.n1961 w_13193_29093.n1958 5.1717
R6191 w_13193_29093.n1165 w_13193_29093.n1164 5.1717
R6192 w_13193_29093.n1233 w_13193_29093.n306 5.1717
R6193 w_13193_29093.n2327 w_13193_29093.n2251 5.13092
R6194 w_13193_29093.n2233 w_13193_29093.n2225 4.97828
R6195 w_13193_29093.n1773 w_13193_29093.n445 4.9157
R6196 w_13193_29093.n1744 w_13193_29093.n1743 4.9157
R6197 w_13193_29093.n1713 w_13193_29093.n1712 4.9157
R6198 w_13193_29093.n2710 w_13193_29093.n2709 4.88834
R6199 w_13193_29093.n2761 w_13193_29093.n2760 4.88834
R6200 w_13193_29093.n230 w_13193_29093.n229 4.57193
R6201 w_13193_29093.n2503 w_13193_29093.n2497 4.57193
R6202 w_13193_29093.n1085 w_13193_29093.n778 4.5005
R6203 w_13193_29093.n1092 w_13193_29093.n1091 4.5005
R6204 w_13193_29093.n1086 w_13193_29093.n750 4.5005
R6205 w_13193_29093.n1088 w_13193_29093.n1087 4.5005
R6206 w_13193_29093.n1087 w_13193_29093.n1086 4.5005
R6207 w_13193_29093.n770 w_13193_29093.n753 4.5005
R6208 w_13193_29093.n2208 w_13193_29093.n265 4.5005
R6209 w_13193_29093.n2544 w_13193_29093.n197 4.49344
R6210 w_13193_29093.n2545 w_13193_29093.n2544 4.49344
R6211 w_13193_29093.n2538 w_13193_29093.n2537 4.49344
R6212 w_13193_29093.n2539 w_13193_29093.n2538 4.49344
R6213 w_13193_29093.n2212 w_13193_29093.n2211 4.42387
R6214 w_13193_29093.n2384 w_13193_29093.n2381 4.36399
R6215 w_13193_29093.n2527 w_13193_29093.n2524 4.36399
R6216 w_13193_29093.n1159 w_13193_29093.t170 4.33832
R6217 w_13193_29093.t286 w_13193_29093.n734 4.33832
R6218 w_13193_29093.n736 w_13193_29093.t37 4.33832
R6219 w_13193_29093.n1147 w_13193_29093.t139 4.33832
R6220 w_13193_29093.n1142 w_13193_29093.n1141 4.26717
R6221 w_13193_29093.n1141 w_13193_29093.n1104 4.26717
R6222 w_13193_29093.n1136 w_13193_29093.n1104 4.26717
R6223 w_13193_29093.n1136 w_13193_29093.n1135 4.26717
R6224 w_13193_29093.n1135 w_13193_29093.n1134 4.26717
R6225 w_13193_29093.n1134 w_13193_29093.n1113 4.26717
R6226 w_13193_29093.n1129 w_13193_29093.n1113 4.26717
R6227 w_13193_29093.n1129 w_13193_29093.n1128 4.26717
R6228 w_13193_29093.n1128 w_13193_29093.n1127 4.26717
R6229 w_13193_29093.n1127 w_13193_29093.n624 4.26717
R6230 w_13193_29093.n1213 w_13193_29093.n624 4.26717
R6231 w_13193_29093.n1073 w_13193_29093.n1028 4.26717
R6232 w_13193_29093.n1029 w_13193_29093.n1028 4.26717
R6233 w_13193_29093.n1066 w_13193_29093.n1029 4.26717
R6234 w_13193_29093.n1066 w_13193_29093.n1065 4.26717
R6235 w_13193_29093.n1065 w_13193_29093.n1064 4.26717
R6236 w_13193_29093.n1064 w_13193_29093.n1039 4.26717
R6237 w_13193_29093.n1059 w_13193_29093.n1039 4.26717
R6238 w_13193_29093.n1059 w_13193_29093.n1058 4.26717
R6239 w_13193_29093.n1058 w_13193_29093.n1057 4.26717
R6240 w_13193_29093.n1057 w_13193_29093.n1050 4.26717
R6241 w_13193_29093.n1052 w_13193_29093.n1050 4.26717
R6242 w_13193_29093.n1543 w_13193_29093.n586 4.26717
R6243 w_13193_29093.n1500 w_13193_29093.n586 4.26717
R6244 w_13193_29093.n1536 w_13193_29093.n1500 4.26717
R6245 w_13193_29093.n1536 w_13193_29093.n1535 4.26717
R6246 w_13193_29093.n1535 w_13193_29093.n1534 4.26717
R6247 w_13193_29093.n1534 w_13193_29093.n1510 4.26717
R6248 w_13193_29093.n1529 w_13193_29093.n1510 4.26717
R6249 w_13193_29093.n1529 w_13193_29093.n1528 4.26717
R6250 w_13193_29093.n1528 w_13193_29093.n1527 4.26717
R6251 w_13193_29093.n1527 w_13193_29093.n1521 4.26717
R6252 w_13193_29093.n1521 w_13193_29093.n383 4.26717
R6253 w_13193_29093.n1377 w_13193_29093.n1336 4.26717
R6254 w_13193_29093.n1377 w_13193_29093.n1376 4.26717
R6255 w_13193_29093.n1376 w_13193_29093.n1375 4.26717
R6256 w_13193_29093.n1375 w_13193_29093.n1344 4.26717
R6257 w_13193_29093.n1370 w_13193_29093.n1344 4.26717
R6258 w_13193_29093.n1370 w_13193_29093.n1369 4.26717
R6259 w_13193_29093.n1369 w_13193_29093.n1368 4.26717
R6260 w_13193_29093.n1368 w_13193_29093.n1353 4.26717
R6261 w_13193_29093.n1363 w_13193_29093.n1353 4.26717
R6262 w_13193_29093.n1363 w_13193_29093.n1362 4.26717
R6263 w_13193_29093.n1362 w_13193_29093.n317 4.26717
R6264 w_13193_29093.n2102 w_13193_29093.n2064 4.26717
R6265 w_13193_29093.n2102 w_13193_29093.n2101 4.26717
R6266 w_13193_29093.n2101 w_13193_29093.n2100 4.26717
R6267 w_13193_29093.n2100 w_13193_29093.n2072 4.26717
R6268 w_13193_29093.n2095 w_13193_29093.n2072 4.26717
R6269 w_13193_29093.n2095 w_13193_29093.n2094 4.26717
R6270 w_13193_29093.n2094 w_13193_29093.n2093 4.26717
R6271 w_13193_29093.n2093 w_13193_29093.n2081 4.26717
R6272 w_13193_29093.n2088 w_13193_29093.n2081 4.26717
R6273 w_13193_29093.n2088 w_13193_29093.n273 4.26717
R6274 w_13193_29093.n2183 w_13193_29093.n273 4.26717
R6275 w_13193_29093.n1832 w_13193_29093.n388 4.26717
R6276 w_13193_29093.n1832 w_13193_29093.n1831 4.26717
R6277 w_13193_29093.n1831 w_13193_29093.n1830 4.26717
R6278 w_13193_29093.n1830 w_13193_29093.n396 4.26717
R6279 w_13193_29093.n1825 w_13193_29093.n396 4.26717
R6280 w_13193_29093.n1825 w_13193_29093.n1824 4.26717
R6281 w_13193_29093.n1824 w_13193_29093.n1823 4.26717
R6282 w_13193_29093.n1823 w_13193_29093.n405 4.26717
R6283 w_13193_29093.n1818 w_13193_29093.n405 4.26717
R6284 w_13193_29093.n1818 w_13193_29093.n1817 4.26717
R6285 w_13193_29093.n1817 w_13193_29093.n1816 4.26717
R6286 w_13193_29093.n2250 VGND 4.1224
R6287 w_13193_29093.n1383 w_13193_29093.n1213 3.98272
R6288 w_13193_29093.n1052 w_13193_29093.n495 3.98272
R6289 w_13193_29093.n1838 w_13193_29093.n383 3.98272
R6290 w_13193_29093.n2108 w_13193_29093.n317 3.98272
R6291 w_13193_29093.n2183 w_13193_29093.n274 3.98272
R6292 w_13193_29093.n1816 w_13193_29093.n1803 3.98272
R6293 w_13193_29093.n2547 w_13193_29093.n2546 3.8278
R6294 w_13193_29093.n2550 w_13193_29093.n2549 3.8278
R6295 w_13193_29093.n2541 w_13193_29093.n2540 3.8278
R6296 w_13193_29093.n2029 w_13193_29093.n2027 3.7893
R6297 w_13193_29093.n2028 w_13193_29093.n1937 3.7893
R6298 w_13193_29093.n2036 w_13193_29093.n2035 3.7893
R6299 w_13193_29093.n1935 w_13193_29093.n1934 3.7893
R6300 w_13193_29093.n2044 w_13193_29093.n2042 3.7893
R6301 w_13193_29093.n2043 w_13193_29093.n1932 3.7893
R6302 w_13193_29093.n2051 w_13193_29093.n2050 3.7893
R6303 w_13193_29093.n1930 w_13193_29093.n1929 3.7893
R6304 w_13193_29093.n2060 w_13193_29093.n1926 3.7893
R6305 w_13193_29093.n1020 w_13193_29093.n905 3.7893
R6306 w_13193_29093.n995 w_13193_29093.n988 3.7893
R6307 w_13193_29093.n994 w_13193_29093.n992 3.7893
R6308 w_13193_29093.n991 w_13193_29093.n986 3.7893
R6309 w_13193_29093.n1002 w_13193_29093.n984 3.7893
R6310 w_13193_29093.n1003 w_13193_29093.n983 3.7893
R6311 w_13193_29093.n1008 w_13193_29093.n1006 3.7893
R6312 w_13193_29093.n1007 w_13193_29093.n926 3.7893
R6313 w_13193_29093.n1015 w_13193_29093.n1014 3.7893
R6314 w_13193_29093.n1463 w_13193_29093.n614 3.7893
R6315 w_13193_29093.n1462 w_13193_29093.n615 3.7893
R6316 w_13193_29093.n617 w_13193_29093.n606 3.7893
R6317 w_13193_29093.n605 w_13193_29093.n603 3.7893
R6318 w_13193_29093.n1479 w_13193_29093.n1478 3.7893
R6319 w_13193_29093.n601 w_13193_29093.n600 3.7893
R6320 w_13193_29093.n1487 w_13193_29093.n596 3.7893
R6321 w_13193_29093.n1486 w_13193_29093.n597 3.7893
R6322 w_13193_29093.n598 w_13193_29093.n588 3.7893
R6323 w_13193_29093.n661 w_13193_29093.n660 3.7893
R6324 w_13193_29093.n1157 w_13193_29093.n637 3.7893
R6325 w_13193_29093.n1156 w_13193_29093.n638 3.7893
R6326 w_13193_29093.n722 w_13193_29093.n720 3.7893
R6327 w_13193_29093.n725 w_13193_29093.n724 3.7893
R6328 w_13193_29093.n732 w_13193_29093.n726 3.7893
R6329 w_13193_29093.n731 w_13193_29093.n728 3.7893
R6330 w_13193_29093.n727 w_13193_29093.n659 3.7893
R6331 w_13193_29093.n1151 w_13193_29093.n1150 3.7893
R6332 w_13193_29093.n872 w_13193_29093.n867 3.7893
R6333 w_13193_29093.n871 w_13193_29093.n868 3.7893
R6334 w_13193_29093.n878 w_13193_29093.n811 3.7893
R6335 w_13193_29093.n879 w_13193_29093.n810 3.7893
R6336 w_13193_29093.n884 w_13193_29093.n882 3.7893
R6337 w_13193_29093.n883 w_13193_29093.n805 3.7893
R6338 w_13193_29093.n892 w_13193_29093.n891 3.7893
R6339 w_13193_29093.n806 w_13193_29093.n785 3.7893
R6340 w_13193_29093.n898 w_13193_29093.n897 3.7893
R6341 w_13193_29093.n1550 w_13193_29093.n1549 3.7893
R6342 w_13193_29093.n514 w_13193_29093.n513 3.7893
R6343 w_13193_29093.n1557 w_13193_29093.n1556 3.7893
R6344 w_13193_29093.n1559 w_13193_29093.n1558 3.7893
R6345 w_13193_29093.n1563 w_13193_29093.n1562 3.7893
R6346 w_13193_29093.n511 w_13193_29093.n510 3.7893
R6347 w_13193_29093.n1571 w_13193_29093.n507 3.7893
R6348 w_13193_29093.n1570 w_13193_29093.n508 3.7893
R6349 w_13193_29093.n1746 w_13193_29093.n452 3.7893
R6350 w_13193_29093.n1301 w_13193_29093.n1299 3.7893
R6351 w_13193_29093.n1300 w_13193_29093.n1227 3.7893
R6352 w_13193_29093.n1308 w_13193_29093.n1307 3.7893
R6353 w_13193_29093.n1225 w_13193_29093.n1224 3.7893
R6354 w_13193_29093.n1316 w_13193_29093.n1314 3.7893
R6355 w_13193_29093.n1315 w_13193_29093.n1222 3.7893
R6356 w_13193_29093.n1323 w_13193_29093.n1322 3.7893
R6357 w_13193_29093.n1220 w_13193_29093.n1219 3.7893
R6358 w_13193_29093.n1332 w_13193_29093.n1216 3.7893
R6359 w_13193_29093.n1902 w_13193_29093.n1901 3.7893
R6360 w_13193_29093.n333 w_13193_29093.n332 3.7893
R6361 w_13193_29093.n1910 w_13193_29093.n329 3.7893
R6362 w_13193_29093.n1909 w_13193_29093.n330 3.7893
R6363 w_13193_29093.n369 w_13193_29093.n367 3.7893
R6364 w_13193_29093.n370 w_13193_29093.n366 3.7893
R6365 w_13193_29093.n377 w_13193_29093.n375 3.7893
R6366 w_13193_29093.n376 w_13193_29093.n351 3.7893
R6367 w_13193_29093.n1845 w_13193_29093.n1844 3.7893
R6368 w_13193_29093.n1665 w_13193_29093.n1664 3.7893
R6369 w_13193_29093.n485 w_13193_29093.n484 3.7893
R6370 w_13193_29093.n1673 w_13193_29093.n476 3.7893
R6371 w_13193_29093.n1672 w_13193_29093.n477 3.7893
R6372 w_13193_29093.n482 w_13193_29093.n481 3.7893
R6373 w_13193_29093.n479 w_13193_29093.n466 3.7893
R6374 w_13193_29093.n1687 w_13193_29093.n1686 3.7893
R6375 w_13193_29093.n464 w_13193_29093.n463 3.7893
R6376 w_13193_29093.n1715 w_13193_29093.n460 3.7893
R6377 w_13193_29093.n2246 w_13193_29093.n2245 3.4105
R6378 w_13193_29093.n2245 w_13193_29093.n2241 3.4105
R6379 w_13193_29093.n2251 w_13193_29093.n2241 3.4105
R6380 w_13193_29093.n2248 w_13193_29093.n2239 3.4105
R6381 w_13193_29093.n2251 w_13193_29093.n2239 3.4105
R6382 w_13193_29093.n2251 w_13193_29093.n2250 3.4105
R6383 w_13193_29093.n2671 w_13193_29093.n2670 3.2005
R6384 w_13193_29093.n2637 w_13193_29093.n2636 3.2005
R6385 w_13193_29093.n2615 w_13193_29093.n171 3.2005
R6386 w_13193_29093.n2596 w_13193_29093.n183 3.2005
R6387 w_13193_29093.n2338 w_13193_29093.n2234 3.2005
R6388 w_13193_29093.t258 w_13193_29093.n27 3.13108
R6389 w_13193_29093.n2212 w_13193_29093.n258 2.986
R6390 w_13193_29093.n2553 w_13193_29093.n202 2.8779
R6391 w_13193_29093.n203 w_13193_29093.n202 2.8779
R6392 w_13193_29093.n761 w_13193_29093.n758 2.86505
R6393 w_13193_29093.n763 w_13193_29093.n757 2.86505
R6394 w_13193_29093.n765 w_13193_29093.n764 2.86505
R6395 w_13193_29093.n766 w_13193_29093.n754 2.86505
R6396 w_13193_29093.n766 w_13193_29093.n765 2.86505
R6397 w_13193_29093.n758 w_13193_29093.n757 2.86505
R6398 w_13193_29093.n769 w_13193_29093.n754 2.86505
R6399 w_13193_29093.n764 w_13193_29093.n763 2.86505
R6400 w_13193_29093.n250 w_13193_29093.n248 2.86505
R6401 w_13193_29093.n249 w_13193_29093.n245 2.86505
R6402 w_13193_29093.n253 w_13193_29093.n252 2.86505
R6403 w_13193_29093.n252 w_13193_29093.n242 2.86505
R6404 w_13193_29093.n250 w_13193_29093.n249 2.86505
R6405 w_13193_29093.n253 w_13193_29093.n245 2.86505
R6406 w_13193_29093.n233 w_13193_29093.n222 2.82018
R6407 w_13193_29093.n228 w_13193_29093.n227 2.82018
R6408 w_13193_29093.n2506 w_13193_29093.n2505 2.82018
R6409 w_13193_29093.n2504 w_13193_29093.n2499 2.82018
R6410 w_13193_29093.t267 w_13193_29093.n17 2.68393
R6411 w_13193_29093.n2059 w_13193_29093.n1924 2.6629
R6412 w_13193_29093.n1074 w_13193_29093.n900 2.6629
R6413 w_13193_29093.n979 w_13193_29093.n445 2.6629
R6414 w_13193_29093.n1388 w_13193_29093.n620 2.6629
R6415 w_13193_29093.n1405 w_13193_29093.n582 2.6629
R6416 w_13193_29093.n741 w_13193_29093.n716 2.6629
R6417 w_13193_29093.n1143 w_13193_29093.n1100 2.6629
R6418 w_13193_29093.n1075 w_13193_29093.n899 2.6629
R6419 w_13193_29093.n1545 w_13193_29093.n1544 2.6629
R6420 w_13193_29093.n1745 w_13193_29093.n1744 2.6629
R6421 w_13193_29093.n1331 w_13193_29093.n1214 2.6629
R6422 w_13193_29093.n1923 w_13193_29093.n1922 2.6629
R6423 w_13193_29093.n386 w_13193_29093.n352 2.6629
R6424 w_13193_29093.n1653 w_13193_29093.n387 2.6629
R6425 w_13193_29093.n1714 w_13193_29093.n1713 2.6629
R6426 w_13193_29093.n2385 w_13193_29093.n2379 2.6474
R6427 w_13193_29093.n2384 w_13193_29093.n2383 2.6474
R6428 w_13193_29093.n2528 w_13193_29093.n209 2.6474
R6429 w_13193_29093.n2527 w_13193_29093.n2526 2.6474
R6430 w_13193_29093.n1962 w_13193_29093.n1961 2.4581
R6431 w_13193_29093.n1924 w_13193_29093.n1923 2.4581
R6432 w_13193_29093.n904 w_13193_29093.n900 2.4581
R6433 w_13193_29093.n1390 w_13193_29093.n1388 2.4581
R6434 w_13193_29093.n1544 w_13193_29093.n582 2.4581
R6435 w_13193_29093.n1164 w_13193_29093.n632 2.4581
R6436 w_13193_29093.n1143 w_13193_29093.n741 2.4581
R6437 w_13193_29093.n1100 w_13193_29093.n742 2.4581
R6438 w_13193_29093.n1075 w_13193_29093.n1074 2.4581
R6439 w_13193_29093.n1546 w_13193_29093.n1545 2.4581
R6440 w_13193_29093.n1234 w_13193_29093.n1233 2.4581
R6441 w_13193_29093.n1214 w_13193_29093.n620 2.4581
R6442 w_13193_29093.n1922 w_13193_29093.n319 2.4581
R6443 w_13193_29093.n387 w_13193_29093.n386 2.4581
R6444 w_13193_29093.n1653 w_13193_29093.n1652 2.4581
R6445 w_13193_29093.n263 w_13193_29093.n262 2.44675
R6446 w_13193_29093.n263 w_13193_29093.n259 2.44675
R6447 w_13193_29093.n773 w_13193_29093.n772 2.26187
R6448 w_13193_29093.n1089 w_13193_29093.n1088 2.24063
R6449 w_13193_29093.n777 w_13193_29093.n751 2.24063
R6450 w_13193_29093.n776 w_13193_29093.n752 2.24063
R6451 w_13193_29093.n772 w_13193_29093.n771 2.24063
R6452 w_13193_29093.n1090 w_13193_29093.n749 2.24063
R6453 w_13193_29093.n775 w_13193_29093.n774 2.24063
R6454 w_13193_29093.n1085 w_13193_29093.n1084 2.22018
R6455 w_13193_29093.n1091 w_13193_29093.n747 2.22018
R6456 w_13193_29093.n2208 w_13193_29093.n2207 2.22018
R6457 w_13193_29093.n1143 w_13193_29093.n1142 2.18124
R6458 w_13193_29093.n1074 w_13193_29093.n1073 2.18124
R6459 w_13193_29093.n1544 w_13193_29093.n1543 2.18124
R6460 w_13193_29093.n1336 w_13193_29093.n620 2.18124
R6461 w_13193_29093.n2064 w_13193_29093.n1923 2.18124
R6462 w_13193_29093.n388 w_13193_29093.n387 2.18124
R6463 w_13193_29093.n1962 w_13193_29093.n1939 2.1509
R6464 w_13193_29093.n1021 w_13193_29093.n904 2.1509
R6465 w_13193_29093.n1390 w_13193_29093.n1389 2.1509
R6466 w_13193_29093.n634 w_13193_29093.n632 2.1509
R6467 w_13193_29093.n813 w_13193_29093.n742 2.1509
R6468 w_13193_29093.n1548 w_13193_29093.n1546 2.1509
R6469 w_13193_29093.n1234 w_13193_29093.n1229 2.1509
R6470 w_13193_29093.n1899 w_13193_29093.n319 2.1509
R6471 w_13193_29093.n1652 w_13193_29093.n487 2.1509
R6472 w_13193_29093.n1714 w_13193_29093.n1694 2.13383
R6473 w_13193_29093.n352 w_13193_29093.n349 2.13383
R6474 w_13193_29093.n2059 w_13193_29093.n2058 2.13383
R6475 w_13193_29093.n1745 w_13193_29093.n453 2.13383
R6476 w_13193_29093.n979 w_13193_29093.n978 2.13383
R6477 w_13193_29093.n1406 w_13193_29093.n1405 2.13383
R6478 w_13193_29093.n899 w_13193_29093.n784 2.13383
R6479 w_13193_29093.n716 w_13193_29093.n715 2.13383
R6480 w_13193_29093.n1331 w_13193_29093.n1330 2.13383
R6481 w_13193_29093.n1144 w_13193_29093.n1143 2.08643
R6482 w_13193_29093.n1074 w_13193_29093.n901 2.08643
R6483 w_13193_29093.n1544 w_13193_29093.n583 2.08643
R6484 w_13193_29093.n1382 w_13193_29093.n620 2.08643
R6485 w_13193_29093.n2107 w_13193_29093.n1923 2.08643
R6486 w_13193_29093.n1837 w_13193_29093.n387 2.08643
R6487 w_13193_29093.n2060 w_13193_29093.n2059 1.9461
R6488 w_13193_29093.n1014 w_13193_29093.n979 1.9461
R6489 w_13193_29093.n1405 w_13193_29093.n588 1.9461
R6490 w_13193_29093.n1150 w_13193_29093.n716 1.9461
R6491 w_13193_29093.n899 w_13193_29093.n898 1.9461
R6492 w_13193_29093.n1746 w_13193_29093.n1745 1.9461
R6493 w_13193_29093.n1332 w_13193_29093.n1331 1.9461
R6494 w_13193_29093.n1844 w_13193_29093.n352 1.9461
R6495 w_13193_29093.n1715 w_13193_29093.n1714 1.9461
R6496 w_13193_29093.n229 w_13193_29093.n228 1.71099
R6497 w_13193_29093.n230 w_13193_29093.n222 1.71099
R6498 w_13193_29093.n2504 w_13193_29093.n2503 1.71099
R6499 w_13193_29093.n2505 w_13193_29093.n2497 1.71099
R6500 w_13193_29093.n2246 w_13193_29093.n2240 1.70307
R6501 w_13193_29093.n2248 w_13193_29093.n2247 1.70307
R6502 w_13193_29093.n2244 w_13193_29093.n2243 1.70307
R6503 w_13193_29093.n2245 w_13193_29093.n2242 1.70307
R6504 w_13193_29093.n2250 w_13193_29093.n2249 1.70307
R6505 w_13193_29093.n1712 w_13193_29093.n1711 1.52512
R6506 w_13193_29093.n1773 w_13193_29093.n1772 1.52512
R6507 w_13193_29093.n1743 w_13193_29093.n1741 1.52512
R6508 w_13193_29093.n2465 w_13193_29093.n2213 1.5139
R6509 w_13193_29093.n1958 w_13193_29093.n1957 1.42272
R6510 w_13193_29093.n1166 w_13193_29093.n1165 1.42272
R6511 w_13193_29093.n2150 w_13193_29093.n306 1.42272
R6512 w_13193_29093.n1776 w_13193_29093.n27 1.28415
R6513 w_13193_29093.n2208 w_13193_29093.n264 1.20883
R6514 w_13193_29093.n2209 w_13193_29093.n2208 1.14633
R6515 w_13193_29093.n2153 w_13193_29093.n17 1.11531
R6516 w_13193_29093.n2466 w_13193_29093.n2465 0.9781
R6517 w_13193_29093.n2027 w_13193_29093.n1939 0.8197
R6518 w_13193_29093.n2029 w_13193_29093.n2028 0.8197
R6519 w_13193_29093.n2036 w_13193_29093.n1937 0.8197
R6520 w_13193_29093.n2035 w_13193_29093.n1935 0.8197
R6521 w_13193_29093.n2042 w_13193_29093.n1934 0.8197
R6522 w_13193_29093.n2044 w_13193_29093.n2043 0.8197
R6523 w_13193_29093.n2051 w_13193_29093.n1932 0.8197
R6524 w_13193_29093.n2050 w_13193_29093.n1930 0.8197
R6525 w_13193_29093.n1929 w_13193_29093.n1926 0.8197
R6526 w_13193_29093.n1021 w_13193_29093.n1020 0.8197
R6527 w_13193_29093.n988 w_13193_29093.n905 0.8197
R6528 w_13193_29093.n995 w_13193_29093.n994 0.8197
R6529 w_13193_29093.n992 w_13193_29093.n991 0.8197
R6530 w_13193_29093.n986 w_13193_29093.n984 0.8197
R6531 w_13193_29093.n1003 w_13193_29093.n1002 0.8197
R6532 w_13193_29093.n1006 w_13193_29093.n983 0.8197
R6533 w_13193_29093.n1008 w_13193_29093.n1007 0.8197
R6534 w_13193_29093.n1015 w_13193_29093.n926 0.8197
R6535 w_13193_29093.n1389 w_13193_29093.n614 0.8197
R6536 w_13193_29093.n1463 w_13193_29093.n1462 0.8197
R6537 w_13193_29093.n617 w_13193_29093.n615 0.8197
R6538 w_13193_29093.n606 w_13193_29093.n605 0.8197
R6539 w_13193_29093.n1479 w_13193_29093.n603 0.8197
R6540 w_13193_29093.n1478 w_13193_29093.n601 0.8197
R6541 w_13193_29093.n600 w_13193_29093.n596 0.8197
R6542 w_13193_29093.n1487 w_13193_29093.n1486 0.8197
R6543 w_13193_29093.n598 w_13193_29093.n597 0.8197
R6544 w_13193_29093.n661 w_13193_29093.n634 0.8197
R6545 w_13193_29093.n660 w_13193_29093.n637 0.8197
R6546 w_13193_29093.n1157 w_13193_29093.n1156 0.8197
R6547 w_13193_29093.n720 w_13193_29093.n638 0.8197
R6548 w_13193_29093.n724 w_13193_29093.n722 0.8197
R6549 w_13193_29093.n726 w_13193_29093.n725 0.8197
R6550 w_13193_29093.n732 w_13193_29093.n731 0.8197
R6551 w_13193_29093.n728 w_13193_29093.n727 0.8197
R6552 w_13193_29093.n1151 w_13193_29093.n659 0.8197
R6553 w_13193_29093.n867 w_13193_29093.n813 0.8197
R6554 w_13193_29093.n872 w_13193_29093.n871 0.8197
R6555 w_13193_29093.n868 w_13193_29093.n811 0.8197
R6556 w_13193_29093.n879 w_13193_29093.n878 0.8197
R6557 w_13193_29093.n882 w_13193_29093.n810 0.8197
R6558 w_13193_29093.n884 w_13193_29093.n883 0.8197
R6559 w_13193_29093.n892 w_13193_29093.n805 0.8197
R6560 w_13193_29093.n891 w_13193_29093.n806 0.8197
R6561 w_13193_29093.n897 w_13193_29093.n785 0.8197
R6562 w_13193_29093.n1550 w_13193_29093.n1548 0.8197
R6563 w_13193_29093.n1549 w_13193_29093.n514 0.8197
R6564 w_13193_29093.n1556 w_13193_29093.n513 0.8197
R6565 w_13193_29093.n1558 w_13193_29093.n1557 0.8197
R6566 w_13193_29093.n1563 w_13193_29093.n1559 0.8197
R6567 w_13193_29093.n1562 w_13193_29093.n511 0.8197
R6568 w_13193_29093.n510 w_13193_29093.n507 0.8197
R6569 w_13193_29093.n1571 w_13193_29093.n1570 0.8197
R6570 w_13193_29093.n508 w_13193_29093.n452 0.8197
R6571 w_13193_29093.n1299 w_13193_29093.n1229 0.8197
R6572 w_13193_29093.n1301 w_13193_29093.n1300 0.8197
R6573 w_13193_29093.n1308 w_13193_29093.n1227 0.8197
R6574 w_13193_29093.n1307 w_13193_29093.n1225 0.8197
R6575 w_13193_29093.n1314 w_13193_29093.n1224 0.8197
R6576 w_13193_29093.n1316 w_13193_29093.n1315 0.8197
R6577 w_13193_29093.n1323 w_13193_29093.n1222 0.8197
R6578 w_13193_29093.n1322 w_13193_29093.n1220 0.8197
R6579 w_13193_29093.n1219 w_13193_29093.n1216 0.8197
R6580 w_13193_29093.n1902 w_13193_29093.n1899 0.8197
R6581 w_13193_29093.n1901 w_13193_29093.n333 0.8197
R6582 w_13193_29093.n332 w_13193_29093.n329 0.8197
R6583 w_13193_29093.n1910 w_13193_29093.n1909 0.8197
R6584 w_13193_29093.n367 w_13193_29093.n330 0.8197
R6585 w_13193_29093.n370 w_13193_29093.n369 0.8197
R6586 w_13193_29093.n375 w_13193_29093.n366 0.8197
R6587 w_13193_29093.n377 w_13193_29093.n376 0.8197
R6588 w_13193_29093.n1845 w_13193_29093.n351 0.8197
R6589 w_13193_29093.n1665 w_13193_29093.n487 0.8197
R6590 w_13193_29093.n1664 w_13193_29093.n485 0.8197
R6591 w_13193_29093.n484 w_13193_29093.n476 0.8197
R6592 w_13193_29093.n1673 w_13193_29093.n1672 0.8197
R6593 w_13193_29093.n482 w_13193_29093.n477 0.8197
R6594 w_13193_29093.n481 w_13193_29093.n479 0.8197
R6595 w_13193_29093.n1687 w_13193_29093.n466 0.8197
R6596 w_13193_29093.n1686 w_13193_29093.n464 0.8197
R6597 w_13193_29093.n463 w_13193_29093.n460 0.8197
R6598 w_13193_29093.n2213 w_13193_29093.n2212 0.799839
R6599 w_13193_29093.n2522 w_13193_29093.n210 0.703977
R6600 w_13193_29093.n771 w_13193_29093.n258 0.65675
R6601 w_13193_29093.n1088 w_13193_29093.n776 0.542167
R6602 w_13193_29093.n90 w_13193_29093.n89 0.492597
R6603 w_13193_29093.n2468 w_13193_29093.n2467 0.215014
R6604 w_13193_29093.n2556 w_13193_29093.n2555 0.206967
R6605 w_13193_29093.n2326 w_13193_29093.n2325 0.206942
R6606 w_13193_29093.n2328 w_13193_29093.n2238 0.206942
R6607 w_13193_29093.n2464 w_13193_29093.n2214 0.199496
R6608 w_13193_29093.n2584 w_13193_29093.n2580 0.196005
R6609 w_13193_29093.n1091 w_13193_29093.n1090 0.188
R6610 w_13193_29093.n1087 w_13193_29093.n1085 0.188
R6611 w_13193_29093.n2210 w_13193_29093.n2209 0.188
R6612 w_13193_29093.n2393 w_13193_29093.n2392 0.185879
R6613 w_13193_29093.n90 w_13193_29093.n85 0.15675
R6614 w_13193_29093.n94 w_13193_29093.n85 0.15675
R6615 w_13193_29093.n95 w_13193_29093.n94 0.15675
R6616 w_13193_29093.n96 w_13193_29093.n95 0.15675
R6617 w_13193_29093.n96 w_13193_29093.n83 0.15675
R6618 w_13193_29093.n100 w_13193_29093.n83 0.15675
R6619 w_13193_29093.n101 w_13193_29093.n100 0.15675
R6620 w_13193_29093.n102 w_13193_29093.n101 0.15675
R6621 w_13193_29093.n102 w_13193_29093.n80 0.15675
R6622 w_13193_29093.n108 w_13193_29093.n80 0.15675
R6623 w_13193_29093.n109 w_13193_29093.n108 0.15675
R6624 w_13193_29093.n110 w_13193_29093.n109 0.15675
R6625 w_13193_29093.n110 w_13193_29093.n78 0.15675
R6626 w_13193_29093.n115 w_13193_29093.n78 0.15675
R6627 w_13193_29093.n116 w_13193_29093.n115 0.15675
R6628 w_13193_29093.n117 w_13193_29093.n116 0.15675
R6629 w_13193_29093.n117 w_13193_29093.n76 0.15675
R6630 w_13193_29093.n121 w_13193_29093.n76 0.15675
R6631 w_13193_29093.n122 w_13193_29093.n121 0.15675
R6632 w_13193_29093.n123 w_13193_29093.n122 0.15675
R6633 w_13193_29093.n123 w_13193_29093.n74 0.15675
R6634 w_13193_29093.n129 w_13193_29093.n74 0.15675
R6635 w_13193_29093.n130 w_13193_29093.n129 0.15675
R6636 w_13193_29093.n131 w_13193_29093.n130 0.15675
R6637 w_13193_29093.n131 w_13193_29093.n71 0.15675
R6638 w_13193_29093.n135 w_13193_29093.n71 0.15675
R6639 w_13193_29093.n136 w_13193_29093.n135 0.15675
R6640 w_13193_29093.n2689 w_13193_29093.n136 0.15675
R6641 w_13193_29093.n2689 w_13193_29093.n2688 0.15675
R6642 w_13193_29093.n2688 w_13193_29093.n2687 0.15675
R6643 w_13193_29093.n2687 w_13193_29093.n137 0.15675
R6644 w_13193_29093.n138 w_13193_29093.n137 0.15675
R6645 w_13193_29093.n2682 w_13193_29093.n138 0.15675
R6646 w_13193_29093.n2682 w_13193_29093.n2681 0.15675
R6647 w_13193_29093.n2681 w_13193_29093.n2680 0.15675
R6648 w_13193_29093.n2680 w_13193_29093.n140 0.15675
R6649 w_13193_29093.n2675 w_13193_29093.n140 0.15675
R6650 w_13193_29093.n2675 w_13193_29093.n2674 0.15675
R6651 w_13193_29093.n2674 w_13193_29093.n2673 0.15675
R6652 w_13193_29093.n2673 w_13193_29093.n143 0.15675
R6653 w_13193_29093.n2668 w_13193_29093.n143 0.15675
R6654 w_13193_29093.n2668 w_13193_29093.n2667 0.15675
R6655 w_13193_29093.n2667 w_13193_29093.n2666 0.15675
R6656 w_13193_29093.n2666 w_13193_29093.n146 0.15675
R6657 w_13193_29093.n2661 w_13193_29093.n146 0.15675
R6658 w_13193_29093.n2661 w_13193_29093.n2660 0.15675
R6659 w_13193_29093.n2660 w_13193_29093.n2659 0.15675
R6660 w_13193_29093.n2659 w_13193_29093.n149 0.15675
R6661 w_13193_29093.n2655 w_13193_29093.n149 0.15675
R6662 w_13193_29093.n2655 w_13193_29093.n2654 0.15675
R6663 w_13193_29093.n2654 w_13193_29093.n2653 0.15675
R6664 w_13193_29093.n2653 w_13193_29093.n152 0.15675
R6665 w_13193_29093.n2648 w_13193_29093.n152 0.15675
R6666 w_13193_29093.n2648 w_13193_29093.n2647 0.15675
R6667 w_13193_29093.n2647 w_13193_29093.n2646 0.15675
R6668 w_13193_29093.n2646 w_13193_29093.n155 0.15675
R6669 w_13193_29093.n2642 w_13193_29093.n155 0.15675
R6670 w_13193_29093.n2642 w_13193_29093.n2641 0.15675
R6671 w_13193_29093.n2641 w_13193_29093.n2640 0.15675
R6672 w_13193_29093.n2640 w_13193_29093.n158 0.15675
R6673 w_13193_29093.n2635 w_13193_29093.n158 0.15675
R6674 w_13193_29093.n2635 w_13193_29093.n2634 0.15675
R6675 w_13193_29093.n2634 w_13193_29093.n2633 0.15675
R6676 w_13193_29093.n2633 w_13193_29093.n161 0.15675
R6677 w_13193_29093.n2629 w_13193_29093.n161 0.15675
R6678 w_13193_29093.n2629 w_13193_29093.n2628 0.15675
R6679 w_13193_29093.n2628 w_13193_29093.n165 0.15675
R6680 w_13193_29093.n2624 w_13193_29093.n165 0.15675
R6681 w_13193_29093.n2624 w_13193_29093.n2623 0.15675
R6682 w_13193_29093.n2623 w_13193_29093.n2622 0.15675
R6683 w_13193_29093.n2622 w_13193_29093.n167 0.15675
R6684 w_13193_29093.n2618 w_13193_29093.n167 0.15675
R6685 w_13193_29093.n2618 w_13193_29093.n2617 0.15675
R6686 w_13193_29093.n2617 w_13193_29093.n2616 0.15675
R6687 w_13193_29093.n2616 w_13193_29093.n170 0.15675
R6688 w_13193_29093.n172 w_13193_29093.n170 0.15675
R6689 w_13193_29093.n2611 w_13193_29093.n172 0.15675
R6690 w_13193_29093.n2611 w_13193_29093.n2610 0.15675
R6691 w_13193_29093.n2610 w_13193_29093.n2609 0.15675
R6692 w_13193_29093.n2609 w_13193_29093.n175 0.15675
R6693 w_13193_29093.n2605 w_13193_29093.n175 0.15675
R6694 w_13193_29093.n2605 w_13193_29093.n2604 0.15675
R6695 w_13193_29093.n2604 w_13193_29093.n2603 0.15675
R6696 w_13193_29093.n2603 w_13193_29093.n179 0.15675
R6697 w_13193_29093.n2599 w_13193_29093.n179 0.15675
R6698 w_13193_29093.n2599 w_13193_29093.n2598 0.15675
R6699 w_13193_29093.n2598 w_13193_29093.n2597 0.15675
R6700 w_13193_29093.n2597 w_13193_29093.n182 0.15675
R6701 w_13193_29093.n184 w_13193_29093.n182 0.15675
R6702 w_13193_29093.n2592 w_13193_29093.n184 0.15675
R6703 w_13193_29093.n2592 w_13193_29093.n2591 0.15675
R6704 w_13193_29093.n2591 w_13193_29093.n2590 0.15675
R6705 w_13193_29093.n2590 w_13193_29093.n187 0.15675
R6706 w_13193_29093.n2586 w_13193_29093.n187 0.15675
R6707 w_13193_29093.n2586 w_13193_29093.n2585 0.15675
R6708 w_13193_29093.n2585 w_13193_29093.n2584 0.15675
R6709 w_13193_29093.n2575 w_13193_29093.n191 0.15675
R6710 w_13193_29093.n2575 w_13193_29093.n2574 0.15675
R6711 w_13193_29093.n2574 w_13193_29093.n2573 0.15675
R6712 w_13193_29093.n2573 w_13193_29093.n194 0.15675
R6713 w_13193_29093.n2569 w_13193_29093.n194 0.15675
R6714 w_13193_29093.n2569 w_13193_29093.n2568 0.15675
R6715 w_13193_29093.n2568 w_13193_29093.n2567 0.15675
R6716 w_13193_29093.n2567 w_13193_29093.n196 0.15675
R6717 w_13193_29093.n2563 w_13193_29093.n196 0.15675
R6718 w_13193_29093.n2563 w_13193_29093.n2562 0.15675
R6719 w_13193_29093.n2562 w_13193_29093.n2561 0.15675
R6720 w_13193_29093.n2561 w_13193_29093.n199 0.15675
R6721 w_13193_29093.n2557 w_13193_29093.n199 0.15675
R6722 w_13193_29093.n2557 w_13193_29093.n2556 0.15675
R6723 w_13193_29093.n2325 w_13193_29093.n2254 0.15675
R6724 w_13193_29093.n2321 w_13193_29093.n2254 0.15675
R6725 w_13193_29093.n2321 w_13193_29093.n2320 0.15675
R6726 w_13193_29093.n2320 w_13193_29093.n2319 0.15675
R6727 w_13193_29093.n2319 w_13193_29093.n2256 0.15675
R6728 w_13193_29093.n2257 w_13193_29093.n2256 0.15675
R6729 w_13193_29093.n2314 w_13193_29093.n2257 0.15675
R6730 w_13193_29093.n2314 w_13193_29093.n2313 0.15675
R6731 w_13193_29093.n2313 w_13193_29093.n2312 0.15675
R6732 w_13193_29093.n2312 w_13193_29093.n2263 0.15675
R6733 w_13193_29093.n2308 w_13193_29093.n2263 0.15675
R6734 w_13193_29093.n2308 w_13193_29093.n2307 0.15675
R6735 w_13193_29093.n2307 w_13193_29093.n2306 0.15675
R6736 w_13193_29093.n2306 w_13193_29093.n2265 0.15675
R6737 w_13193_29093.n2267 w_13193_29093.n2265 0.15675
R6738 w_13193_29093.n2301 w_13193_29093.n2267 0.15675
R6739 w_13193_29093.n2301 w_13193_29093.n2300 0.15675
R6740 w_13193_29093.n2300 w_13193_29093.n2299 0.15675
R6741 w_13193_29093.n2299 w_13193_29093.n2269 0.15675
R6742 w_13193_29093.n2295 w_13193_29093.n2269 0.15675
R6743 w_13193_29093.n2295 w_13193_29093.n2294 0.15675
R6744 w_13193_29093.n2294 w_13193_29093.n2293 0.15675
R6745 w_13193_29093.n2293 w_13193_29093.n2272 0.15675
R6746 w_13193_29093.n2288 w_13193_29093.n2272 0.15675
R6747 w_13193_29093.n2288 w_13193_29093.n2287 0.15675
R6748 w_13193_29093.n2287 w_13193_29093.n2286 0.15675
R6749 w_13193_29093.n2286 w_13193_29093.n2275 0.15675
R6750 w_13193_29093.n2282 w_13193_29093.n2275 0.15675
R6751 w_13193_29093.n2282 w_13193_29093.n2281 0.15675
R6752 w_13193_29093.n2281 w_13193_29093.n2220 0.15675
R6753 w_13193_29093.n2220 w_13193_29093.n2218 0.15675
R6754 w_13193_29093.n2451 w_13193_29093.n2218 0.15675
R6755 w_13193_29093.n2452 w_13193_29093.n2451 0.15675
R6756 w_13193_29093.n2453 w_13193_29093.n2452 0.15675
R6757 w_13193_29093.n2456 w_13193_29093.n2453 0.15675
R6758 w_13193_29093.n2456 w_13193_29093.n2455 0.15675
R6759 w_13193_29093.n2455 w_13193_29093.n2214 0.15675
R6760 w_13193_29093.n2332 w_13193_29093.n2238 0.15675
R6761 w_13193_29093.n2333 w_13193_29093.n2332 0.15675
R6762 w_13193_29093.n2334 w_13193_29093.n2333 0.15675
R6763 w_13193_29093.n2334 w_13193_29093.n2236 0.15675
R6764 w_13193_29093.n2236 w_13193_29093.n2235 0.15675
R6765 w_13193_29093.n2339 w_13193_29093.n2235 0.15675
R6766 w_13193_29093.n2340 w_13193_29093.n2339 0.15675
R6767 w_13193_29093.n2340 w_13193_29093.n2232 0.15675
R6768 w_13193_29093.n2345 w_13193_29093.n2232 0.15675
R6769 w_13193_29093.n2346 w_13193_29093.n2345 0.15675
R6770 w_13193_29093.n2347 w_13193_29093.n2346 0.15675
R6771 w_13193_29093.n2347 w_13193_29093.n2230 0.15675
R6772 w_13193_29093.n2351 w_13193_29093.n2230 0.15675
R6773 w_13193_29093.n2352 w_13193_29093.n2351 0.15675
R6774 w_13193_29093.n2353 w_13193_29093.n2352 0.15675
R6775 w_13193_29093.n2353 w_13193_29093.n2228 0.15675
R6776 w_13193_29093.n2357 w_13193_29093.n2228 0.15675
R6777 w_13193_29093.n2358 w_13193_29093.n2357 0.15675
R6778 w_13193_29093.n2359 w_13193_29093.n2358 0.15675
R6779 w_13193_29093.n2430 w_13193_29093.n2359 0.15675
R6780 w_13193_29093.n2430 w_13193_29093.n2429 0.15675
R6781 w_13193_29093.n2429 w_13193_29093.n2428 0.15675
R6782 w_13193_29093.n2428 w_13193_29093.n2361 0.15675
R6783 w_13193_29093.n2423 w_13193_29093.n2361 0.15675
R6784 w_13193_29093.n2423 w_13193_29093.n2422 0.15675
R6785 w_13193_29093.n2422 w_13193_29093.n2421 0.15675
R6786 w_13193_29093.n2421 w_13193_29093.n2363 0.15675
R6787 w_13193_29093.n2417 w_13193_29093.n2363 0.15675
R6788 w_13193_29093.n2417 w_13193_29093.n2416 0.15675
R6789 w_13193_29093.n2416 w_13193_29093.n2415 0.15675
R6790 w_13193_29093.n2415 w_13193_29093.n2365 0.15675
R6791 w_13193_29093.n2411 w_13193_29093.n2365 0.15675
R6792 w_13193_29093.n2411 w_13193_29093.n2410 0.15675
R6793 w_13193_29093.n2410 w_13193_29093.n2409 0.15675
R6794 w_13193_29093.n2406 w_13193_29093.n2405 0.15675
R6795 w_13193_29093.n2405 w_13193_29093.n2404 0.15675
R6796 w_13193_29093.n2404 w_13193_29093.n2370 0.15675
R6797 w_13193_29093.n2400 w_13193_29093.n2370 0.15675
R6798 w_13193_29093.n2400 w_13193_29093.n2399 0.15675
R6799 w_13193_29093.n2399 w_13193_29093.n2398 0.15675
R6800 w_13193_29093.n2398 w_13193_29093.n2373 0.15675
R6801 w_13193_29093.n2394 w_13193_29093.n2373 0.15675
R6802 w_13193_29093.n2394 w_13193_29093.n2393 0.15675
R6803 w_13193_29093.n2757 w_13193_29093.n35 0.15675
R6804 w_13193_29093.n2753 w_13193_29093.n2752 0.15675
R6805 w_13193_29093.n2752 w_13193_29093.n2751 0.15675
R6806 w_13193_29093.n2751 w_13193_29093.n39 0.15675
R6807 w_13193_29093.n2747 w_13193_29093.n2746 0.15675
R6808 w_13193_29093.n2746 w_13193_29093.n2745 0.15675
R6809 w_13193_29093.n2745 w_13193_29093.n45 0.15675
R6810 w_13193_29093.n2741 w_13193_29093.n2740 0.15675
R6811 w_13193_29093.n2740 w_13193_29093.n2739 0.15675
R6812 w_13193_29093.n2739 w_13193_29093.n49 0.15675
R6813 w_13193_29093.n2735 w_13193_29093.n2734 0.15675
R6814 w_13193_29093.n2734 w_13193_29093.n2733 0.15675
R6815 w_13193_29093.n2733 w_13193_29093.n53 0.15675
R6816 w_13193_29093.n2729 w_13193_29093.n2728 0.15675
R6817 w_13193_29093.n2468 w_13193_29093.n239 0.15675
R6818 w_13193_29093.n2472 w_13193_29093.n239 0.15675
R6819 w_13193_29093.n2473 w_13193_29093.n2472 0.15675
R6820 w_13193_29093.n2474 w_13193_29093.n2473 0.15675
R6821 w_13193_29093.n2474 w_13193_29093.n236 0.15675
R6822 w_13193_29093.n236 w_13193_29093.n235 0.15675
R6823 w_13193_29093.n2479 w_13193_29093.n235 0.15675
R6824 w_13193_29093.n2480 w_13193_29093.n2479 0.15675
R6825 w_13193_29093.n2481 w_13193_29093.n2480 0.15675
R6826 w_13193_29093.n2481 w_13193_29093.n220 0.15675
R6827 w_13193_29093.n2485 w_13193_29093.n220 0.15675
R6828 w_13193_29093.n2486 w_13193_29093.n2485 0.15675
R6829 w_13193_29093.n2487 w_13193_29093.n2486 0.15675
R6830 w_13193_29093.n2487 w_13193_29093.n217 0.15675
R6831 w_13193_29093.n2491 w_13193_29093.n217 0.15675
R6832 w_13193_29093.n2492 w_13193_29093.n2491 0.15675
R6833 w_13193_29093.n2493 w_13193_29093.n2492 0.15675
R6834 w_13193_29093.n2493 w_13193_29093.n214 0.15675
R6835 w_13193_29093.n2508 w_13193_29093.n214 0.15675
R6836 w_13193_29093.n2509 w_13193_29093.n2508 0.15675
R6837 w_13193_29093.n2510 w_13193_29093.n2509 0.15675
R6838 w_13193_29093.n2510 w_13193_29093.n212 0.15675
R6839 w_13193_29093.n2515 w_13193_29093.n212 0.15675
R6840 w_13193_29093.n2516 w_13193_29093.n2515 0.15675
R6841 w_13193_29093.n2517 w_13193_29093.n2516 0.15675
R6842 w_13193_29093.n2517 w_13193_29093.n210 0.15675
R6843 w_13193_29093.n2579 w_13193_29093.n191 0.141125
R6844 w_13193_29093.n2466 w_13193_29093.n192 0.1321
R6845 w_13193_29093.n2727 w_13193_29093.n2726 0.131895
R6846 w_13193_29093.n1093 w_13193_29093.n1092 0.1255
R6847 w_13193_29093.n1083 w_13193_29093.n778 0.1255
R6848 w_13193_29093.n2206 w_13193_29093.n265 0.1255
R6849 w_13193_29093.n2406 w_13193_29093.n2368 0.109875
R6850 w_13193_29093.n2758 w_13193_29093.n34 0.0986461
R6851 w_13193_29093.n2758 w_13193_29093.n2757 0.09425
R6852 w_13193_29093.n2753 w_13193_29093.n38 0.09425
R6853 w_13193_29093.n2747 w_13193_29093.n44 0.09425
R6854 w_13193_29093.n2741 w_13193_29093.n48 0.09425
R6855 w_13193_29093.n2735 w_13193_29093.n52 0.09425
R6856 w_13193_29093.n2729 w_13193_29093.n56 0.09425
R6857 w_13193_29093.n38 w_13193_29093.n35 0.063
R6858 w_13193_29093.n44 w_13193_29093.n39 0.063
R6859 w_13193_29093.n48 w_13193_29093.n45 0.063
R6860 w_13193_29093.n52 w_13193_29093.n49 0.063
R6861 w_13193_29093.n56 w_13193_29093.n53 0.063
R6862 w_13193_29093.n2728 w_13193_29093.n2727 0.063
R6863 w_13193_29093.n1093 w_13193_29093.n747 0.0626438
R6864 w_13193_29093.n1084 w_13193_29093.n1083 0.0626438
R6865 w_13193_29093.n2207 w_13193_29093.n2206 0.0626438
R6866 w_13193_29093.n2409 w_13193_29093.n2368 0.047375
R6867 w_13193_29093.n2579 w_13193_29093.n2578 0.0430057
R6868 w_13193_29093.n1088 w_13193_29093.n751 0.0421667
R6869 w_13193_29093.n1090 w_13193_29093.n1089 0.0217373
R6870 w_13193_29093.n1087 w_13193_29093.n777 0.0217373
R6871 w_13193_29093.n1089 w_13193_29093.n750 0.0217373
R6872 w_13193_29093.n777 w_13193_29093.n750 0.0217373
R6873 w_13193_29093.n770 w_13193_29093.n752 0.0217373
R6874 w_13193_29093.n772 w_13193_29093.n753 0.0217373
R6875 w_13193_29093.n771 w_13193_29093.n752 0.0217373
R6876 w_13193_29093.n1086 w_13193_29093.n749 0.0217373
R6877 w_13193_29093.n775 w_13193_29093.n753 0.0217373
R6878 w_13193_29093.n751 w_13193_29093.n749 0.0217373
R6879 w_13193_29093.n773 w_13193_29093.n770 0.0217373
R6880 w_13193_29093.n774 w_13193_29093.n773 0.0217373
R6881 w_13193_29093.n776 w_13193_29093.n775 0.0217373
R6882 w_13193_29093.n2248 w_13193_29093.n2245 0.01225
R6883 w_13193_29093.n2247 w_13193_29093.n2241 0.0068649
R6884 w_13193_29093.n2243 w_13193_29093.n2239 0.0068649
R6885 w_13193_29093.n2250 w_13193_29093.n2242 0.0068649
R6886 w_13193_29093.n2251 w_13193_29093.n2240 0.0068649
R6887 w_13193_29093.n2249 w_13193_29093.n2248 0.0068649
R6888 w_13193_29093.n2247 w_13193_29093.n2246 0.0068649
R6889 w_13193_29093.n2244 w_13193_29093.n2240 0.0068649
R6890 w_13193_29093.n2243 w_13193_29093.n2241 0.0068649
R6891 w_13193_29093.n2242 w_13193_29093.n2239 0.0068649
R6892 w_13193_29093.n2249 w_13193_29093.n2244 0.0068649
R6893 a_18974_25970.n10 a_18974_25970.t8 1834.89
R6894 a_18974_25970.n0 a_18974_25970.t10 377.567
R6895 a_18974_25970.n5 a_18974_25970.t11 377.567
R6896 a_18974_25970.n1 a_18974_25970.n0 257.067
R6897 a_18974_25970.n4 a_18974_25970.n3 257.067
R6898 a_18974_25970.n6 a_18974_25970.n5 257.067
R6899 a_18974_25970.n9 a_18974_25970.n8 159.12
R6900 a_18974_25970.n11 a_18974_25970.n10 154.319
R6901 a_18974_25970.n9 a_18974_25970.n7 153.601
R6902 a_18974_25970.n10 a_18974_25970.n2 152
R6903 a_18974_25970.n4 a_18974_25970.t0 120.501
R6904 a_18974_25970.n3 a_18974_25970.t6 120.501
R6905 a_18974_25970.n1 a_18974_25970.t2 120.501
R6906 a_18974_25970.n0 a_18974_25970.t12 120.501
R6907 a_18974_25970.n6 a_18974_25970.t4 120.501
R6908 a_18974_25970.n5 a_18974_25970.t9 120.501
R6909 a_18974_25970.n10 a_18974_25970.n9 108.8
R6910 a_18974_25970.n2 a_18974_25970.n1 85.6894
R6911 a_18974_25970.n3 a_18974_25970.n2 85.6894
R6912 a_18974_25970.n7 a_18974_25970.n4 85.6894
R6913 a_18974_25970.n7 a_18974_25970.n6 85.6894
R6914 a_18974_25970.n8 a_18974_25970.t1 19.7005
R6915 a_18974_25970.n8 a_18974_25970.t5 19.7005
R6916 a_18974_25970.n11 a_18974_25970.t3 19.7005
R6917 a_18974_25970.t7 a_18974_25970.n11 19.7005
R6918 a_18974_25060.n6 a_18974_25060.t8 580.49
R6919 a_18974_25060.n2 a_18974_25060.t11 317.317
R6920 a_18974_25060.n4 a_18974_25060.t12 317.317
R6921 a_18974_25060.n3 a_18974_25060.n2 257.067
R6922 a_18974_25060.n9 a_18974_25060.n8 257.067
R6923 a_18974_25060.n5 a_18974_25060.n4 257.067
R6924 a_18974_25060.n11 a_18974_25060.n10 155.201
R6925 a_18974_25060.n7 a_18974_25060.n6 152
R6926 a_18974_25060.n1 a_18974_25060.n0 120.981
R6927 a_18974_25060.n12 a_18974_25060.n11 120.981
R6928 a_18974_25060.n11 a_18974_25060.n1 102.4
R6929 a_18974_25060.n10 a_18974_25060.n3 85.6894
R6930 a_18974_25060.n10 a_18974_25060.n9 85.6894
R6931 a_18974_25060.n8 a_18974_25060.n7 85.6894
R6932 a_18974_25060.n7 a_18974_25060.n5 85.6894
R6933 a_18974_25060.n8 a_18974_25060.t0 60.2505
R6934 a_18974_25060.n9 a_18974_25060.t6 60.2505
R6935 a_18974_25060.n3 a_18974_25060.t2 60.2505
R6936 a_18974_25060.n2 a_18974_25060.t9 60.2505
R6937 a_18974_25060.n5 a_18974_25060.t4 60.2505
R6938 a_18974_25060.n4 a_18974_25060.t10 60.2505
R6939 a_18974_25060.n0 a_18974_25060.t1 24.0005
R6940 a_18974_25060.n0 a_18974_25060.t5 24.0005
R6941 a_18974_25060.n12 a_18974_25060.t3 24.0005
R6942 a_18974_25060.t7 a_18974_25060.n12 24.0005
R6943 a_18974_25060.n6 a_18974_25060.n1 3.2005
R6944 a_18180_33430.n0 a_18180_33430.n3 199.935
R6945 a_18180_33430.n0 a_18180_33430.n1 199.53
R6946 a_18180_33430.n0 a_18180_33430.n2 199.53
R6947 a_18180_33430.n0 a_18180_33430.n4 199.53
R6948 a_18180_33430.n5 a_18180_33430.n0 199.53
R6949 a_18180_33430.n0 a_18180_33430.t8 98.9938
R6950 a_18180_33430.n1 a_18180_33430.t1 48.0005
R6951 a_18180_33430.n1 a_18180_33430.t7 48.0005
R6952 a_18180_33430.n2 a_18180_33430.t6 48.0005
R6953 a_18180_33430.n2 a_18180_33430.t2 48.0005
R6954 a_18180_33430.n4 a_18180_33430.t3 48.0005
R6955 a_18180_33430.n4 a_18180_33430.t4 48.0005
R6956 a_18180_33430.n3 a_18180_33430.t5 48.0005
R6957 a_18180_33430.n3 a_18180_33430.t10 48.0005
R6958 a_18180_33430.t0 a_18180_33430.n5 48.0005
R6959 a_18180_33430.n5 a_18180_33430.t9 48.0005
R6960 a_25860_20180.n1 a_25860_20180.t3 600.206
R6961 a_25860_20180.t0 a_25860_20180.n5 576.192
R6962 a_25860_20180.n2 a_25860_20180.n1 568.072
R6963 a_25860_20180.n4 a_25860_20180.n2 392.486
R6964 a_25860_20180.n0 a_25860_20180.t2 289.791
R6965 a_25860_20180.n5 a_25860_20180.n4 168.067
R6966 a_25860_20180.n3 a_25860_20180.n0 97.9242
R6967 a_25860_20180.n4 a_25860_20180.n3 37.7572
R6968 a_25860_20180.n2 a_25860_20180.t4 32.1338
R6969 a_25860_20180.n1 a_25860_20180.t5 32.1338
R6970 a_25860_20180.n3 a_25860_20180.t1 32.1338
R6971 a_25860_20180.n5 a_25860_20180.n0 28.3357
R6972 a_26640_21760.t1 a_26640_21760.n0 708.125
R6973 a_26640_21760.t1 a_26640_21760.n1 708.125
R6974 a_26640_21760.n1 a_26640_21760.t2 410.519
R6975 a_26640_21760.n0 a_26640_21760.t0 305.649
R6976 a_26640_21760.n1 a_26640_21760.n0 21.3338
R6977 a_24280_30060.t0 a_24280_30060.n2 500.086
R6978 a_24280_30060.n0 a_24280_30060.t2 490.034
R6979 a_24280_30060.t0 a_24280_30060.n2 461.389
R6980 a_24280_30060.n1 a_24280_30060.n0 449.233
R6981 a_24280_30060.n0 a_24280_30060.t3 345.433
R6982 a_24280_30060.n1 a_24280_30060.t1 177.577
R6983 a_24280_30060.n2 a_24280_30060.n1 48.3899
R6984 a_23100_30460.n1 a_23100_30460.t2 586.433
R6985 a_23100_30460.n2 a_23100_30460.n1 456.351
R6986 a_23100_30460.n0 a_23100_30460.t4 441.834
R6987 a_23100_30460.n0 a_23100_30460.t5 393.634
R6988 a_23100_30460.n3 a_23100_30460.n2 328.733
R6989 a_23100_30460.t1 a_23100_30460.n3 288.37
R6990 a_23100_30460.n1 a_23100_30460.t3 249.034
R6991 a_23100_30460.n3 a_23100_30460.t0 177.577
R6992 a_23100_30460.n2 a_23100_30460.n0 152.633
R6993 a_14730_30630.n8 a_14730_30630.n7 314.526
R6994 a_14730_30630.n9 a_14730_30630.t12 287.764
R6995 a_14730_30630.n10 a_14730_30630.t10 287.764
R6996 a_14730_30630.n9 a_14730_30630.t8 287.591
R6997 a_14730_30630.n11 a_14730_30630.t11 287.012
R6998 a_14730_30630.n12 a_14730_30630.t9 287.012
R6999 a_14730_30630.n14 a_14730_30630.t2 158.046
R7000 a_14730_30630.n6 a_14730_30630.n4 107.079
R7001 a_14730_30630.n6 a_14730_30630.n5 104.828
R7002 a_14730_30630.n22 a_14730_30630.n21 83.7933
R7003 a_14730_30630.n1 a_14730_30630.n0 83.5719
R7004 a_14730_30630.n18 a_14730_30630.n17 83.5719
R7005 a_14730_30630.n7 a_14730_30630.t0 39.4005
R7006 a_14730_30630.n7 a_14730_30630.t3 39.4005
R7007 a_14730_30630.t1 a_14730_30630.n16 36.6632
R7008 a_14730_30630.n17 a_14730_30630.n0 26.074
R7009 a_14730_30630.n22 a_14730_30630.n0 26.074
R7010 a_14730_30630.n17 a_14730_30630.t1 25.7843
R7011 a_14730_30630.n15 a_14730_30630.n14 23.9067
R7012 a_14730_30630.n23 a_14730_30630.n22 20.5696
R7013 a_14730_30630.n4 a_14730_30630.t7 13.1338
R7014 a_14730_30630.n4 a_14730_30630.t6 13.1338
R7015 a_14730_30630.n5 a_14730_30630.t4 13.1338
R7016 a_14730_30630.n5 a_14730_30630.t5 13.1338
R7017 a_14730_30630.n14 a_14730_30630.n13 13.0943
R7018 a_14730_30630.n13 a_14730_30630.n8 10.7505
R7019 a_14730_30630.n13 a_14730_30630.n12 6.78086
R7020 a_14730_30630.n8 a_14730_30630.n6 2.0005
R7021 a_14730_30630.n16 a_14730_30630.n3 1.80777
R7022 a_14730_30630.n21 a_14730_30630.n20 1.56836
R7023 a_14730_30630.n20 a_14730_30630.n19 1.5505
R7024 a_14730_30630.n3 a_14730_30630.n2 1.5505
R7025 a_14730_30630.n21 a_14730_30630.n1 1.43912
R7026 a_14730_30630.n19 a_14730_30630.n18 1.25468
R7027 a_14730_30630.n16 a_14730_30630.n15 1.04793
R7028 a_14730_30630.n18 a_14730_30630.n3 0.590702
R7029 a_14730_30630.n11 a_14730_30630.n10 0.579071
R7030 a_14730_30630.n19 a_14730_30630.n1 0.406264
R7031 a_14730_30630.n12 a_14730_30630.n11 0.282643
R7032 a_14730_30630.n10 a_14730_30630.n9 0.2755
R7033 a_14730_30630.n20 a_14730_30630.n2 0.0183571
R7034 a_14730_30630.n15 a_14730_30630.n2 0.0106786
R7035 a_19910_25340.n4 a_19910_25340.n0 427.647
R7036 a_19910_25340.n1 a_19910_25340.t7 297.233
R7037 a_19910_25340.n5 a_19910_25340.n4 210.601
R7038 a_19910_25340.n3 a_19910_25340.t3 174.056
R7039 a_19910_25340.n2 a_19910_25340.n1 160.667
R7040 a_19910_25340.n4 a_19910_25340.n3 152
R7041 a_19910_25340.n1 a_19910_25340.t6 136.567
R7042 a_19910_25340.n2 a_19910_25340.t1 136.567
R7043 a_19910_25340.t4 a_19910_25340.n5 60.0005
R7044 a_19910_25340.n5 a_19910_25340.t2 60.0005
R7045 a_19910_25340.n0 a_19910_25340.t5 49.2505
R7046 a_19910_25340.n0 a_19910_25340.t0 49.2505
R7047 a_19910_25340.n3 a_19910_25340.n2 37.4894
R7048 a_19910_24200.n1 a_19910_24200.t6 377.567
R7049 a_19910_24200.n0 a_19910_24200.t8 297.233
R7050 a_19910_24200.n2 a_19910_24200.n1 233.476
R7051 a_19910_24200.n1 a_19910_24200.t7 216.9
R7052 a_19910_24200.n2 a_19910_24200.n0 213.998
R7053 a_19910_24200.n7 a_19910_24200.n6 205.862
R7054 a_19910_24200.n4 a_19910_24200.n3 178.903
R7055 a_19910_24200.n6 a_19910_24200.n5 178.901
R7056 a_19910_24200.n0 a_19910_24200.t9 136.567
R7057 a_19910_24200.n4 a_19910_24200.n2 66.8859
R7058 a_19910_24200.n6 a_19910_24200.n4 57.6005
R7059 a_19910_24200.n5 a_19910_24200.t3 24.6255
R7060 a_19910_24200.n5 a_19910_24200.t0 24.6255
R7061 a_19910_24200.n3 a_19910_24200.t5 24.6255
R7062 a_19910_24200.n3 a_19910_24200.t4 24.6255
R7063 a_19910_24200.t1 a_19910_24200.n7 15.0005
R7064 a_19910_24200.n7 a_19910_24200.t2 15.0005
R7065 a_19040_22530.t4 a_19040_22530.n6 1128.89
R7066 a_19040_22530.n3 a_19040_22530.n2 459.132
R7067 a_19040_22530.n2 a_19040_22530.n0 386.048
R7068 a_19040_22530.n2 a_19040_22530.n1 265
R7069 a_19040_22530.n3 a_19040_22530.t7 232.968
R7070 a_19040_22530.n4 a_19040_22530.t8 232.968
R7071 a_19040_22530.n5 a_19040_22530.t5 232.968
R7072 a_19040_22530.n6 a_19040_22530.t6 232.968
R7073 a_19040_22530.n4 a_19040_22530.n3 160.667
R7074 a_19040_22530.n5 a_19040_22530.n4 160.667
R7075 a_19040_22530.n6 a_19040_22530.n5 160.667
R7076 a_19040_22530.n1 a_19040_22530.t1 60.0005
R7077 a_19040_22530.n1 a_19040_22530.t0 60.0005
R7078 a_19040_22530.n0 a_19040_22530.t2 49.2505
R7079 a_19040_22530.n0 a_19040_22530.t3 49.2505
R7080 a_20480_25210.n5 a_20480_25210.n3 522.322
R7081 a_20480_25210.n11 a_20480_25210.t7 384.967
R7082 a_20480_25210.n0 a_20480_25210.t4 384.967
R7083 a_20480_25210.n0 a_20480_25210.t6 376.56
R7084 a_20480_25210.t8 a_20480_25210.n11 376.56
R7085 a_20480_25210.n8 a_20480_25210.n7 322.046
R7086 a_20480_25210.n10 a_20480_25210.n9 322.046
R7087 a_20480_25210.n2 a_20480_25210.n1 320.902
R7088 a_20480_25210.n5 a_20480_25210.n4 160.721
R7089 a_20480_25210.n10 a_20480_25210.n8 70.4005
R7090 a_20480_25210.n1 a_20480_25210.t11 49.2505
R7091 a_20480_25210.n1 a_20480_25210.t5 49.2505
R7092 a_20480_25210.n7 a_20480_25210.t10 49.2505
R7093 a_20480_25210.n7 a_20480_25210.t12 49.2505
R7094 a_20480_25210.n9 a_20480_25210.t9 49.2505
R7095 a_20480_25210.n9 a_20480_25210.t13 49.2505
R7096 a_20480_25210.n6 a_20480_25210.n5 37.763
R7097 a_20480_25210.n6 a_20480_25210.n2 36.2672
R7098 a_20480_25210.n4 a_20480_25210.t2 19.7005
R7099 a_20480_25210.n4 a_20480_25210.t0 19.7005
R7100 a_20480_25210.n3 a_20480_25210.t3 19.7005
R7101 a_20480_25210.n3 a_20480_25210.t1 19.7005
R7102 a_20480_25210.n8 a_20480_25210.n6 17.0672
R7103 a_20480_25210.n2 a_20480_25210.n0 9.6005
R7104 a_20480_25210.n11 a_20480_25210.n10 9.6005
R7105 a_26320_28790.n4 a_26320_28790.t0 782.52
R7106 a_26320_28790.t11 a_26320_28790.t2 514.134
R7107 a_26320_28790.t5 a_26320_28790.n5 377.567
R7108 a_26320_28790.n0 a_26320_28790.t3 377.567
R7109 a_26320_28790.n3 a_26320_28790.n2 321.334
R7110 a_26320_28790.n6 a_26320_28790.t5 318.702
R7111 a_26320_28790.n6 a_26320_28790.t11 307.909
R7112 a_26320_28790.n4 a_26320_28790.n3 275.341
R7113 a_26320_28790.n5 a_26320_28790.t7 265.101
R7114 a_26320_28790.t1 a_26320_28790.n7 233
R7115 a_26320_28790.n0 a_26320_28790.t8 168.701
R7116 a_26320_28790.n5 a_26320_28790.t6 136.567
R7117 a_26320_28790.n1 a_26320_28790.t4 136.567
R7118 a_26320_28790.n2 a_26320_28790.t9 136.567
R7119 a_26320_28790.n2 a_26320_28790.n1 128.534
R7120 a_26320_28790.n3 a_26320_28790.t10 126.927
R7121 a_26320_28790.n1 a_26320_28790.n0 48.2005
R7122 a_26320_28790.n7 a_26320_28790.n6 38.2642
R7123 a_26320_28790.n7 a_26320_28790.n4 26.4538
R7124 a_26420_30200.n0 a_26420_30200.t0 691.534
R7125 a_26420_30200.n1 a_26420_30200.t2 691.534
R7126 a_26420_30200.n0 a_26420_30200.t3 527.867
R7127 a_26420_30200.t1 a_26420_30200.n1 343.401
R7128 a_26420_30200.n1 a_26420_30200.n0 92.8005
R7129 a_13532_27710.t0 a_13532_27710.t16 170.145
R7130 a_13532_27710.t17 a_13532_27710.t10 0.1603
R7131 a_13532_27710.t11 a_13532_27710.t17 0.1603
R7132 a_13532_27710.t19 a_13532_27710.t11 0.1603
R7133 a_13532_27710.t3 a_13532_27710.t19 0.1603
R7134 a_13532_27710.t6 a_13532_27710.t3 0.1603
R7135 a_13532_27710.t4 a_13532_27710.t6 0.1603
R7136 a_13532_27710.t8 a_13532_27710.t4 0.1603
R7137 a_13532_27710.t14 a_13532_27710.t8 0.1603
R7138 a_13532_27710.t13 a_13532_27710.t20 0.1603
R7139 a_13532_27710.t7 a_13532_27710.t13 0.1603
R7140 a_13532_27710.t12 a_13532_27710.t7 0.1603
R7141 a_13532_27710.t5 a_13532_27710.t12 0.1603
R7142 a_13532_27710.t2 a_13532_27710.t5 0.1603
R7143 a_13532_27710.t18 a_13532_27710.t2 0.1603
R7144 a_13532_27710.t1 a_13532_27710.t18 0.1603
R7145 a_13532_27710.t16 a_13532_27710.t1 0.1603
R7146 a_13532_27710.t15 a_13532_27710.n0 0.159278
R7147 a_13532_27710.t20 a_13532_27710.t15 0.137822
R7148 a_13532_27710.n0 a_13532_27710.t14 0.1368
R7149 a_13532_27710.n0 a_13532_27710.t9 0.00152174
R7150 a_23100_27770.n0 a_23100_27770.t5 1180.9
R7151 a_23100_27770.n2 a_23100_27770.t3 522.168
R7152 a_23100_27770.t0 a_23100_27770.n4 458.818
R7153 a_23100_27770.t0 a_23100_27770.n4 429.281
R7154 a_23100_27770.n1 a_23100_27770.n0 417.733
R7155 a_23100_27770.n0 a_23100_27770.t2 232.968
R7156 a_23100_27770.n3 a_23100_27770.n2 228.8
R7157 a_23100_27770.n1 a_23100_27770.t4 217.905
R7158 a_23100_27770.n3 a_23100_27770.t1 164.775
R7159 a_23100_27770.n4 a_23100_27770.n3 60.248
R7160 a_23100_27770.n2 a_23100_27770.n1 15.063
R7161 a_23130_27670.t1 a_23130_27670.n8 458.818
R7162 a_23130_27670.t1 a_23130_27670.n8 429.281
R7163 a_23130_27670.n3 a_23130_27670.t6 326.658
R7164 a_23130_27670.t3 a_23130_27670.n5 297.233
R7165 a_23130_27670.n4 a_23130_27670.t7 297.233
R7166 a_23130_27670.n0 a_23130_27670.t2 294.829
R7167 a_23130_27670.n2 a_23130_27670.n1 257.067
R7168 a_23130_27670.n7 a_23130_27670.n6 242.494
R7169 a_23130_27670.n3 a_23130_27670.n2 226.942
R7170 a_23130_27670.n6 a_23130_27670.n1 226.942
R7171 a_23130_27670.n5 a_23130_27670.n4 216.9
R7172 a_23130_27670.n0 a_23130_27670.t0 151.976
R7173 a_23130_27670.n7 a_23130_27670.n0 137.601
R7174 a_23130_27670.n6 a_23130_27670.t3 92.3838
R7175 a_23130_27670.t7 a_23130_27670.n3 92.3838
R7176 a_23130_27670.n2 a_23130_27670.t5 80.3338
R7177 a_23130_27670.n4 a_23130_27670.t5 80.3338
R7178 a_23130_27670.t4 a_23130_27670.n1 80.3338
R7179 a_23130_27670.n5 a_23130_27670.t4 80.3338
R7180 a_23130_27670.n8 a_23130_27670.n7 34.648
R7181 a_19940_23090.n3 a_19940_23090.n1 418.048
R7182 a_19940_23090.n3 a_19940_23090.n2 360.447
R7183 a_19940_23090.n5 a_19940_23090.t8 328.175
R7184 a_19940_23090.n14 a_19940_23090.n0 306.601
R7185 a_19940_23090.t15 a_19940_23090.n9 297.233
R7186 a_19940_23090.n8 a_19940_23090.t14 297.233
R7187 a_19940_23090.t14 a_19940_23090.n7 297.233
R7188 a_19940_23090.n15 a_19940_23090.n14 249
R7189 a_19940_23090.n9 a_19940_23090.n8 216.9
R7190 a_19940_23090.n7 a_19940_23090.n6 216.9
R7191 a_19940_23090.n11 a_19940_23090.n10 210.351
R7192 a_19940_23090.n4 a_19940_23090.n3 208
R7193 a_19940_23090.n14 a_19940_23090.n13 208
R7194 a_19940_23090.n10 a_19940_23090.n6 180.75
R7195 a_19940_23090.n5 a_19940_23090.t6 118.627
R7196 a_19940_23090.n10 a_19940_23090.t15 92.3838
R7197 a_19940_23090.n7 a_19940_23090.t11 80.3338
R7198 a_19940_23090.n8 a_19940_23090.t11 80.3338
R7199 a_19940_23090.t10 a_19940_23090.n6 80.3338
R7200 a_19940_23090.n9 a_19940_23090.t10 80.3338
R7201 a_19940_23090.n13 a_19940_23090.t12 76.4829
R7202 a_19940_23090.n12 a_19940_23090.n11 73.0531
R7203 a_19940_23090.n4 a_19940_23090.t13 70.0829
R7204 a_19940_23090.n11 a_19940_23090.n5 62.8355
R7205 a_19940_23090.n0 a_19940_23090.t2 60.0005
R7206 a_19940_23090.n0 a_19940_23090.t1 60.0005
R7207 a_19940_23090.t4 a_19940_23090.n15 60.0005
R7208 a_19940_23090.n15 a_19940_23090.t3 60.0005
R7209 a_19940_23090.n13 a_19940_23090.n12 57.6005
R7210 a_19940_23090.n12 a_19940_23090.n4 54.4005
R7211 a_19940_23090.n1 a_19940_23090.t5 49.2505
R7212 a_19940_23090.n1 a_19940_23090.t9 49.2505
R7213 a_19940_23090.n2 a_19940_23090.t7 49.2505
R7214 a_19940_23090.n2 a_19940_23090.t0 49.2505
R7215 a_23100_30570.n4 a_23100_30570.n0 1295.28
R7216 a_23100_30570.n0 a_23100_30570.t3 586.433
R7217 a_23100_30570.n1 a_23100_30570.t5 388.813
R7218 a_23100_30570.n1 a_23100_30570.t6 356.68
R7219 a_23100_30570.n0 a_23100_30570.t4 249.034
R7220 a_23100_30570.n3 a_23100_30570.n1 225.601
R7221 a_23100_30570.t2 a_23100_30570.n4 221.411
R7222 a_23100_30570.n3 a_23100_30570.n2 163.677
R7223 a_23100_30570.n4 a_23100_30570.n3 84.24
R7224 a_23100_30570.n2 a_23100_30570.t0 24.0005
R7225 a_23100_30570.n2 a_23100_30570.t1 24.0005
R7226 a_23550_30490.t0 a_23550_30490.t1 39.4005
R7227 a_23100_30980.n0 a_23100_30980.t3 517.347
R7228 a_23100_30980.n2 a_23100_30980.n0 417.574
R7229 a_23100_30980.n2 a_23100_30980.n1 244.715
R7230 a_23100_30980.n0 a_23100_30980.t4 228.148
R7231 a_23100_30980.t1 a_23100_30980.n2 221.411
R7232 a_23100_30980.n1 a_23100_30980.t0 24.0005
R7233 a_23100_30980.n1 a_23100_30980.t2 24.0005
R7234 a_19250_24340.n6 a_19250_24340.n4 482.582
R7235 a_19250_24340.n10 a_19250_24340.t4 304.634
R7236 a_19250_24340.n0 a_19250_24340.t1 304.634
R7237 a_19250_24340.n0 a_19250_24340.t3 276.289
R7238 a_19250_24340.t5 a_19250_24340.n10 276.289
R7239 a_19250_24340.n2 a_19250_24340.n1 210.601
R7240 a_19250_24340.n9 a_19250_24340.n8 210.601
R7241 a_19250_24340.n7 a_19250_24340.n3 207.4
R7242 a_19250_24340.n6 a_19250_24340.n5 120.981
R7243 a_19250_24340.n7 a_19250_24340.n2 64.0005
R7244 a_19250_24340.n9 a_19250_24340.n7 64.0005
R7245 a_19250_24340.n1 a_19250_24340.t12 60.0005
R7246 a_19250_24340.n1 a_19250_24340.t2 60.0005
R7247 a_19250_24340.n3 a_19250_24340.t13 60.0005
R7248 a_19250_24340.n3 a_19250_24340.t11 60.0005
R7249 a_19250_24340.n8 a_19250_24340.t6 60.0005
R7250 a_19250_24340.n8 a_19250_24340.t0 60.0005
R7251 a_19250_24340.n7 a_19250_24340.n6 47.363
R7252 a_19250_24340.n5 a_19250_24340.t9 24.0005
R7253 a_19250_24340.n5 a_19250_24340.t7 24.0005
R7254 a_19250_24340.n4 a_19250_24340.t8 24.0005
R7255 a_19250_24340.n4 a_19250_24340.t10 24.0005
R7256 a_19250_24340.n2 a_19250_24340.n0 9.6005
R7257 a_19250_24340.n10 a_19250_24340.n9 9.6005
R7258 a_19190_29290.n15 a_19190_29290.t18 310.488
R7259 a_19190_29290.n1 a_19190_29290.t21 310.488
R7260 a_19190_29290.n6 a_19190_29290.t17 310.488
R7261 a_19190_29290.n4 a_19190_29290.n0 297.433
R7262 a_19190_29290.n9 a_19190_29290.n5 297.433
R7263 a_19190_29290.n19 a_19190_29290.n18 297.433
R7264 a_19190_29290.n13 a_19190_29290.t13 248.133
R7265 a_19190_29290.n13 a_19190_29290.n12 199.383
R7266 a_19190_29290.n14 a_19190_29290.n11 194.883
R7267 a_19190_29290.n17 a_19190_29290.t10 184.097
R7268 a_19190_29290.n3 a_19190_29290.t6 184.097
R7269 a_19190_29290.n8 a_19190_29290.t4 184.097
R7270 a_19190_29290.n16 a_19190_29290.n15 167.094
R7271 a_19190_29290.n2 a_19190_29290.n1 167.094
R7272 a_19190_29290.n7 a_19190_29290.n6 167.094
R7273 a_19190_29290.n18 a_19190_29290.n17 161.3
R7274 a_19190_29290.n4 a_19190_29290.n3 161.3
R7275 a_19190_29290.n9 a_19190_29290.n8 161.3
R7276 a_19190_29290.n16 a_19190_29290.t8 120.501
R7277 a_19190_29290.n15 a_19190_29290.t19 120.501
R7278 a_19190_29290.n2 a_19190_29290.t0 120.501
R7279 a_19190_29290.n1 a_19190_29290.t20 120.501
R7280 a_19190_29290.n7 a_19190_29290.t2 120.501
R7281 a_19190_29290.n6 a_19190_29290.t22 120.501
R7282 a_19190_29290.n12 a_19190_29290.t16 48.0005
R7283 a_19190_29290.n12 a_19190_29290.t12 48.0005
R7284 a_19190_29290.n11 a_19190_29290.t14 48.0005
R7285 a_19190_29290.n11 a_19190_29290.t15 48.0005
R7286 a_19190_29290.n17 a_19190_29290.n16 40.7027
R7287 a_19190_29290.n3 a_19190_29290.n2 40.7027
R7288 a_19190_29290.n8 a_19190_29290.n7 40.7027
R7289 a_19190_29290.n0 a_19190_29290.t1 39.4005
R7290 a_19190_29290.n0 a_19190_29290.t7 39.4005
R7291 a_19190_29290.n5 a_19190_29290.t3 39.4005
R7292 a_19190_29290.n5 a_19190_29290.t5 39.4005
R7293 a_19190_29290.n19 a_19190_29290.t9 39.4005
R7294 a_19190_29290.t11 a_19190_29290.n19 39.4005
R7295 a_19190_29290.n10 a_19190_29290.n4 6.6255
R7296 a_19190_29290.n10 a_19190_29290.n9 6.6255
R7297 a_19190_29290.n14 a_19190_29290.n13 5.2505
R7298 a_19190_29290.n18 a_19190_29290.n10 4.5005
R7299 a_19190_29290.n18 a_19190_29290.n14 0.78175
R7300 a_17540_31010.n1 a_17540_31010.t7 238.322
R7301 a_17540_31010.n1 a_17540_31010.t6 238.322
R7302 a_17540_31010.n3 a_17540_31010.n1 168.8
R7303 a_17540_31010.n0 a_17540_31010.t1 130
R7304 a_17540_31010.n5 a_17540_31010.n4 105.171
R7305 a_17540_31010.n3 a_17540_31010.n2 105.171
R7306 a_17540_31010.n0 a_17540_31010.t0 83.3658
R7307 a_17540_31010.n4 a_17540_31010.n0 35.4806
R7308 a_17540_31010.n2 a_17540_31010.t3 13.1338
R7309 a_17540_31010.n2 a_17540_31010.t2 13.1338
R7310 a_17540_31010.n5 a_17540_31010.t4 13.1338
R7311 a_17540_31010.t5 a_17540_31010.n5 13.1338
R7312 a_17540_31010.n4 a_17540_31010.n3 3.3755
R7313 a_26390_26310.n9 a_26390_26310.t0 729.933
R7314 a_26390_26310.n8 a_26390_26310.t1 729.933
R7315 a_26390_26310.n3 a_26390_26310.n2 718.41
R7316 a_26390_26310.n2 a_26390_26310.n1 660.706
R7317 a_26390_26310.n0 a_26390_26310.t11 361.5
R7318 a_26390_26310.n7 a_26390_26310.n6 342.757
R7319 a_26390_26310.n0 a_26390_26310.t4 281.168
R7320 a_26390_26310.t2 a_26390_26310.n9 260.733
R7321 a_26390_26310.n4 a_26390_26310.n3 224.934
R7322 a_26390_26310.n7 a_26390_26310.t3 190.123
R7323 a_26390_26310.n8 a_26390_26310.n7 180.8
R7324 a_26390_26310.n3 a_26390_26310.t8 168.701
R7325 a_26390_26310.n0 a_26390_26310.t10 152.633
R7326 a_26390_26310.n1 a_26390_26310.t6 152.633
R7327 a_26390_26310.n4 a_26390_26310.t12 136.567
R7328 a_26390_26310.n5 a_26390_26310.t9 136.567
R7329 a_26390_26310.n6 a_26390_26310.t5 136.567
R7330 a_26390_26310.n2 a_26390_26310.t7 131.976
R7331 a_26390_26310.n1 a_26390_26310.n0 128.534
R7332 a_26390_26310.n5 a_26390_26310.n4 128.534
R7333 a_26390_26310.n6 a_26390_26310.n5 128.534
R7334 a_26390_26310.n9 a_26390_26310.n8 57.6005
R7335 a_26420_26230.t0 a_26420_26230.t1 96.0005
R7336 a_26420_26340.n0 a_26420_26340.t1 713.933
R7337 a_26420_26340.n0 a_26420_26340.t2 314.233
R7338 a_26420_26340.t0 a_26420_26340.n0 308.2
R7339 a_18180_28430.n6 a_18180_28430.n1 199.935
R7340 a_18180_28430.n1 a_18180_28430.n5 199.53
R7341 a_18180_28430.n1 a_18180_28430.n4 199.53
R7342 a_18180_28430.n0 a_18180_28430.n3 199.53
R7343 a_18180_28430.n0 a_18180_28430.n2 199.53
R7344 a_18180_28430.n0 a_18180_28430.t10 55.175
R7345 a_18180_28430.n5 a_18180_28430.t5 48.0005
R7346 a_18180_28430.n5 a_18180_28430.t0 48.0005
R7347 a_18180_28430.n4 a_18180_28430.t2 48.0005
R7348 a_18180_28430.n4 a_18180_28430.t9 48.0005
R7349 a_18180_28430.n3 a_18180_28430.t6 48.0005
R7350 a_18180_28430.n3 a_18180_28430.t1 48.0005
R7351 a_18180_28430.n2 a_18180_28430.t3 48.0005
R7352 a_18180_28430.n2 a_18180_28430.t8 48.0005
R7353 a_18180_28430.t4 a_18180_28430.n6 48.0005
R7354 a_18180_28430.n6 a_18180_28430.t7 48.0005
R7355 a_18180_28430.n1 a_18180_28430.n0 1.09425
R7356 a_14990_33500.n3 a_14990_33500.t6 291.503
R7357 a_14990_33500.n3 a_14990_33500.t10 291.288
R7358 a_14990_33500.n4 a_14990_33500.t8 291.288
R7359 a_14990_33500.n5 a_14990_33500.t9 291.288
R7360 a_14990_33500.n6 a_14990_33500.t7 291.288
R7361 a_14990_33500.t0 a_14990_33500.n8 165.601
R7362 a_14990_33500.n8 a_14990_33500.t5 108.424
R7363 a_14990_33500.n2 a_14990_33500.n0 105.609
R7364 a_14990_33500.n2 a_14990_33500.n1 104.484
R7365 a_14990_33500.n8 a_14990_33500.n7 21.4246
R7366 a_14990_33500.n7 a_14990_33500.n2 14.2349
R7367 a_14990_33500.n0 a_14990_33500.t4 13.1338
R7368 a_14990_33500.n0 a_14990_33500.t3 13.1338
R7369 a_14990_33500.n1 a_14990_33500.t2 13.1338
R7370 a_14990_33500.n1 a_14990_33500.t1 13.1338
R7371 a_14990_33500.n7 a_14990_33500.n6 6.43621
R7372 a_14990_33500.n4 a_14990_33500.n3 0.643357
R7373 a_14990_33500.n6 a_14990_33500.n5 0.643357
R7374 a_14990_33500.n5 a_14990_33500.n4 0.214786
R7375 a_26390_27520.n0 a_26390_27520.t0 663.801
R7376 a_26390_27520.t5 a_26390_27520.t3 514.134
R7377 a_26390_27520.n0 a_26390_27520.t5 479.284
R7378 a_26390_27520.n3 a_26390_27520.n2 320.7
R7379 a_26390_27520.t1 a_26390_27520.n3 275.454
R7380 a_26390_27520.n2 a_26390_27520.t2 265.101
R7381 a_26390_27520.n1 a_26390_27520.t6 265.101
R7382 a_26390_27520.n1 a_26390_27520.t4 136.567
R7383 a_26390_27520.n2 a_26390_27520.n1 112.468
R7384 a_26390_27520.n3 a_26390_27520.n0 97.9205
R7385 a_26310_26200.n8 a_26310_26200.n7 949.764
R7386 a_26310_26200.n3 a_26310_26200.n2 895.144
R7387 a_26310_26200.t10 a_26310_26200.t8 819.4
R7388 a_26310_26200.n10 a_26310_26200.n9 628.734
R7389 a_26310_26200.n2 a_26310_26200.n1 496.262
R7390 a_26310_26200.n0 a_26310_26200.t5 361.5
R7391 a_26310_26200.n8 a_26310_26200.t10 336.25
R7392 a_26310_26200.n7 a_26310_26200.n6 321.334
R7393 a_26310_26200.n0 a_26310_26200.t7 281.168
R7394 a_26310_26200.n9 a_26310_26200.t0 257.534
R7395 a_26310_26200.n4 a_26310_26200.n3 208.868
R7396 a_26310_26200.n4 a_26310_26200.t3 168.701
R7397 a_26310_26200.n3 a_26310_26200.t14 168.701
R7398 a_26310_26200.n0 a_26310_26200.t4 152.633
R7399 a_26310_26200.n1 a_26310_26200.t11 152.633
R7400 a_26310_26200.n5 a_26310_26200.t12 136.567
R7401 a_26310_26200.n6 a_26310_26200.t6 136.567
R7402 a_26310_26200.n2 a_26310_26200.t9 131.976
R7403 a_26310_26200.n1 a_26310_26200.n0 128.534
R7404 a_26310_26200.n6 a_26310_26200.n5 128.534
R7405 a_26310_26200.n7 a_26310_26200.t13 126.927
R7406 a_26310_26200.n10 a_26310_26200.t1 78.8005
R7407 a_26310_26200.t2 a_26310_26200.n10 78.8005
R7408 a_26310_26200.n5 a_26310_26200.n4 48.2005
R7409 a_26310_26200.n9 a_26310_26200.n8 11.2005
R7410 a_24280_30570.n4 a_24280_30570.n3 1295.28
R7411 a_24280_30570.n3 a_24280_30570.t4 586.433
R7412 a_24280_30570.n0 a_24280_30570.t3 388.813
R7413 a_24280_30570.n0 a_24280_30570.t5 356.68
R7414 a_24280_30570.n3 a_24280_30570.t6 249.034
R7415 a_24280_30570.n2 a_24280_30570.n0 225.601
R7416 a_24280_30570.t1 a_24280_30570.n4 221.411
R7417 a_24280_30570.n2 a_24280_30570.n1 163.678
R7418 a_24280_30570.n4 a_24280_30570.n2 84.24
R7419 a_24280_30570.n1 a_24280_30570.t2 24.0005
R7420 a_24280_30570.n1 a_24280_30570.t0 24.0005
R7421 a_24310_31390.t0 a_24310_31390.t1 39.4005
R7422 a_23100_30050.t4 a_23100_30050.t5 835.467
R7423 a_23100_30050.n3 a_23100_30050.t4 564.496
R7424 a_23100_30050.n2 a_23100_30050.t6 538.234
R7425 a_23100_30050.n1 a_23100_30050.t8 517.347
R7426 a_23100_30050.n3 a_23100_30050.n2 431.12
R7427 a_23100_30050.n4 a_23100_30050.n1 369.601
R7428 a_23100_30050.n2 a_23100_30050.t7 297.233
R7429 a_23100_30050.n5 a_23100_30050.n0 244.716
R7430 a_23100_30050.n1 a_23100_30050.t3 228.148
R7431 a_23100_30050.t2 a_23100_30050.n5 221.411
R7432 a_23100_30050.n5 a_23100_30050.n4 47.9734
R7433 a_23100_30050.n4 a_23100_30050.n3 39.5568
R7434 a_23100_30050.n0 a_23100_30050.t1 24.0005
R7435 a_23100_30050.n0 a_23100_30050.t0 24.0005
R7436 a_24280_31090.n2 a_24280_31090.n1 1295.28
R7437 a_24280_31090.t6 a_24280_31090.t4 1188.93
R7438 a_24280_31090.t4 a_24280_31090.t3 835.467
R7439 a_24280_31090.n1 a_24280_31090.t5 586.433
R7440 a_24280_31090.n1 a_24280_31090.t6 249.034
R7441 a_24280_31090.n2 a_24280_31090.n0 247.916
R7442 a_24280_31090.t1 a_24280_31090.n2 221.411
R7443 a_24280_31090.n0 a_24280_31090.t2 24.0005
R7444 a_24280_31090.n0 a_24280_31090.t0 24.0005
R7445 a_24310_31010.t0 a_24310_31010.t1 39.4005
R7446 a_26390_28180.n0 a_26390_28180.t3 729.933
R7447 a_26390_28180.n1 a_26390_28180.t4 547.134
R7448 a_26390_28180.n0 a_26390_28180.t1 260.733
R7449 a_26390_28180.n2 a_26390_28180.n1 212.733
R7450 a_26390_28180.n1 a_26390_28180.n0 57.6005
R7451 a_26390_28180.t2 a_26390_28180.n2 48.0005
R7452 a_26390_28180.n2 a_26390_28180.t0 48.0005
R7453 V_CONT.n0 V_CONT.t8 1132.7
R7454 V_CONT.n1 V_CONT.n0 915.801
R7455 V_CONT.n12 V_CONT.n2 706.639
R7456 V_CONT.n2 V_CONT.n1 385.601
R7457 V_CONT.n4 V_CONT.t11 377.567
R7458 V_CONT.n3 V_CONT.t9 297.233
R7459 V_CONT.n5 V_CONT.n3 237.851
R7460 V_CONT.n9 V_CONT.n7 236.501
R7461 V_CONT.n5 V_CONT.n4 232.809
R7462 V_CONT.n0 V_CONT.t15 216.9
R7463 V_CONT.n1 V_CONT.t12 216.9
R7464 V_CONT.n2 V_CONT.t13 216.9
R7465 V_CONT.n4 V_CONT.t10 216.9
R7466 V_CONT.n9 V_CONT.n8 178.901
R7467 V_CONT.n3 V_CONT.t14 136.567
R7468 V_CONT.t7 V_CONT.n13 126.139
R7469 V_CONT.n11 V_CONT.n10 117.546
R7470 V_CONT.n10 V_CONT.n6 113.061
R7471 V_CONT.n11 V_CONT.n5 51.2088
R7472 V_CONT.n10 V_CONT.n9 35.2005
R7473 V_CONT.n8 V_CONT.t1 24.6255
R7474 V_CONT.n8 V_CONT.t0 24.6255
R7475 V_CONT.n7 V_CONT.t3 24.6255
R7476 V_CONT.n7 V_CONT.t2 24.6255
R7477 V_CONT.n6 V_CONT.t4 15.0005
R7478 V_CONT.n6 V_CONT.t6 15.0005
R7479 V_CONT.n12 V_CONT.n11 11.5239
R7480 V_CONT.n13 V_CONT.t5 3.82928
R7481 V_CONT.n13 V_CONT.n12 0.09475
R7482 a_25860_21760.n0 a_25860_21760.t1 284.2
R7483 a_25860_21760.n0 a_25860_21760.t2 233
R7484 a_25860_21760.t0 a_25860_21760.n0 184.191
R7485 a_19940_24490.n1 a_19940_24490.t7 335.793
R7486 a_19940_24490.n5 a_19940_24490.n4 325.248
R7487 a_19940_24490.n4 a_19940_24490.n0 313
R7488 a_19940_24490.n3 a_19940_24490.t4 252.248
R7489 a_19940_24490.n1 a_19940_24490.t6 216.9
R7490 a_19940_24490.n2 a_19940_24490.t2 216.9
R7491 a_19940_24490.n2 a_19940_24490.n1 160.667
R7492 a_19940_24490.n4 a_19940_24490.n3 152
R7493 a_19940_24490.n0 a_19940_24490.t0 60.0005
R7494 a_19940_24490.n0 a_19940_24490.t1 60.0005
R7495 a_19940_24490.n5 a_19940_24490.t5 49.2505
R7496 a_19940_24490.t3 a_19940_24490.n5 49.2505
R7497 a_19940_24490.n3 a_19940_24490.n2 35.3472
R7498 a_23100_29610.n0 a_23100_29610.t3 490.034
R7499 a_23100_29610.n1 a_23100_29610.n0 457.233
R7500 a_23100_29610.n0 a_23100_29610.t4 345.433
R7501 a_23100_29610.n2 a_23100_29610.n1 226.887
R7502 a_23100_29610.n1 a_23100_29610.t1 172.458
R7503 a_23100_29610.t0 a_23100_29610.n2 19.7005
R7504 a_23100_29610.n2 a_23100_29610.t2 19.7005
R7505 a_23100_29280.t1 a_23100_29280.n2 500.086
R7506 a_23100_29280.n0 a_23100_29280.t2 490.034
R7507 a_23100_29280.t1 a_23100_29280.n2 461.389
R7508 a_23100_29280.n1 a_23100_29280.n0 449.233
R7509 a_23100_29280.n0 a_23100_29280.t3 345.433
R7510 a_23100_29280.n1 a_23100_29280.t0 177.577
R7511 a_23100_29280.n2 a_23100_29280.n1 48.3899
R7512 a_14558_34050.n0 a_14558_34050.t25 403.952
R7513 a_14558_34050.n18 a_14558_34050.t26 403.755
R7514 a_14558_34050.n17 a_14558_34050.t23 403.755
R7515 a_14558_34050.n16 a_14558_34050.t14 403.755
R7516 a_14558_34050.n15 a_14558_34050.t27 403.755
R7517 a_14558_34050.n14 a_14558_34050.t18 403.755
R7518 a_14558_34050.n13 a_14558_34050.t11 403.755
R7519 a_14558_34050.n12 a_14558_34050.t24 403.755
R7520 a_14558_34050.n11 a_14558_34050.t16 403.755
R7521 a_14558_34050.n10 a_14558_34050.t29 403.755
R7522 a_14558_34050.n9 a_14558_34050.t20 403.755
R7523 a_14558_34050.n8 a_14558_34050.t21 403.755
R7524 a_14558_34050.n7 a_14558_34050.t17 403.755
R7525 a_14558_34050.n6 a_14558_34050.t10 403.755
R7526 a_14558_34050.n5 a_14558_34050.t22 403.755
R7527 a_14558_34050.n4 a_14558_34050.t13 403.755
R7528 a_14558_34050.n3 a_14558_34050.t15 403.755
R7529 a_14558_34050.n2 a_14558_34050.t28 403.755
R7530 a_14558_34050.n1 a_14558_34050.t19 403.755
R7531 a_14558_34050.n0 a_14558_34050.t12 403.755
R7532 a_14558_34050.n26 a_14558_34050.n25 301.933
R7533 a_14558_34050.n24 a_14558_34050.n23 301.933
R7534 a_14558_34050.n22 a_14558_34050.n21 301.933
R7535 a_14558_34050.n20 a_14558_34050.n19 301.933
R7536 a_14558_34050.t0 a_14558_34050.n27 157.238
R7537 a_14558_34050.n20 a_14558_34050.t1 103.826
R7538 a_14558_34050.n25 a_14558_34050.t3 39.4005
R7539 a_14558_34050.n25 a_14558_34050.t5 39.4005
R7540 a_14558_34050.n23 a_14558_34050.t6 39.4005
R7541 a_14558_34050.n23 a_14558_34050.t7 39.4005
R7542 a_14558_34050.n21 a_14558_34050.t8 39.4005
R7543 a_14558_34050.n21 a_14558_34050.t9 39.4005
R7544 a_14558_34050.n19 a_14558_34050.t4 39.4005
R7545 a_14558_34050.n19 a_14558_34050.t2 39.4005
R7546 a_14558_34050.n27 a_14558_34050.n18 10.3335
R7547 a_14558_34050.n27 a_14558_34050.n26 5.313
R7548 a_14558_34050.n9 a_14558_34050.n8 1.6255
R7549 a_14558_34050.n26 a_14558_34050.n24 1.1255
R7550 a_14558_34050.n24 a_14558_34050.n22 1.1255
R7551 a_14558_34050.n22 a_14558_34050.n20 1.1255
R7552 a_14558_34050.n18 a_14558_34050.n17 0.196929
R7553 a_14558_34050.n17 a_14558_34050.n16 0.196929
R7554 a_14558_34050.n16 a_14558_34050.n15 0.196929
R7555 a_14558_34050.n15 a_14558_34050.n14 0.196929
R7556 a_14558_34050.n14 a_14558_34050.n13 0.196929
R7557 a_14558_34050.n13 a_14558_34050.n12 0.196929
R7558 a_14558_34050.n12 a_14558_34050.n11 0.196929
R7559 a_14558_34050.n11 a_14558_34050.n10 0.196929
R7560 a_14558_34050.n10 a_14558_34050.n9 0.196929
R7561 a_14558_34050.n8 a_14558_34050.n7 0.196929
R7562 a_14558_34050.n7 a_14558_34050.n6 0.196929
R7563 a_14558_34050.n6 a_14558_34050.n5 0.196929
R7564 a_14558_34050.n5 a_14558_34050.n4 0.196929
R7565 a_14558_34050.n4 a_14558_34050.n3 0.196929
R7566 a_14558_34050.n3 a_14558_34050.n2 0.196929
R7567 a_14558_34050.n2 a_14558_34050.n1 0.196929
R7568 a_14558_34050.n1 a_14558_34050.n0 0.196929
R7569 a_22190_29430.n5 a_22190_29430.n4 1269.42
R7570 a_22190_29430.n11 a_22190_29430.n10 297.663
R7571 a_22190_29430.n21 a_22190_29430.n20 297.663
R7572 a_22190_29430.n19 a_22190_29430.n18 297.663
R7573 a_22190_29430.n17 a_22190_29430.n15 297.663
R7574 a_22190_29430.n14 a_22190_29430.n13 297.663
R7575 a_22190_29430.n25 a_22190_29430.n24 297.663
R7576 a_22190_29430.n5 a_22190_29430.t13 275.325
R7577 a_22190_29430.n7 a_22190_29430.n6 248.4
R7578 a_22190_29430.n2 a_22190_29430.t15 239.3
R7579 a_22190_29430.n2 a_22190_29430.t0 207.504
R7580 a_22190_29430.n8 a_22190_29430.n2 166.232
R7581 a_22190_29430.n4 a_22190_29430.t19 151.792
R7582 a_22190_29430.n6 a_22190_29430.t11 140.583
R7583 a_22190_29430.n6 a_22190_29430.t13 140.583
R7584 a_22190_29430.n7 a_22190_29430.n3 98.6614
R7585 a_22190_29430.t11 a_22190_29430.n5 80.3338
R7586 a_22190_29430.n4 a_22190_29430.t18 44.2902
R7587 a_22190_29430.n10 a_22190_29430.t16 39.4005
R7588 a_22190_29430.n10 a_22190_29430.t4 39.4005
R7589 a_22190_29430.n20 a_22190_29430.t3 39.4005
R7590 a_22190_29430.n20 a_22190_29430.t8 39.4005
R7591 a_22190_29430.n18 a_22190_29430.t7 39.4005
R7592 a_22190_29430.n18 a_22190_29430.t1 39.4005
R7593 a_22190_29430.n15 a_22190_29430.t5 39.4005
R7594 a_22190_29430.n15 a_22190_29430.t9 39.4005
R7595 a_22190_29430.n13 a_22190_29430.t2 39.4005
R7596 a_22190_29430.n13 a_22190_29430.t17 39.4005
R7597 a_22190_29430.n25 a_22190_29430.t6 39.4005
R7598 a_22190_29430.t10 a_22190_29430.n25 39.4005
R7599 a_22190_29430.n8 a_22190_29430.n7 17.0229
R7600 a_22190_29430.n3 a_22190_29430.t14 15.0005
R7601 a_22190_29430.n3 a_22190_29430.t12 15.0005
R7602 a_22190_29430.n23 a_22190_29430.n11 4.84425
R7603 a_22190_29430.n16 a_22190_29430.n14 4.84425
R7604 a_22190_29430.n17 a_22190_29430.n16 4.5005
R7605 a_22190_29430.n19 a_22190_29430.n12 4.5005
R7606 a_22190_29430.n22 a_22190_29430.n21 4.5005
R7607 a_22190_29430.n24 a_22190_29430.n23 4.5005
R7608 a_22190_29430.n9 a_22190_29430.n8 9.35425
R7609 a_22190_29430.n0 a_22190_29430.n14 1.85607
R7610 a_22190_29430.n11 a_22190_29430.n9 1.74185
R7611 a_22190_29430.n21 a_22190_29430.n1 1.74185
R7612 a_22190_29430.n0 a_22190_29430.n19 1.74185
R7613 a_22190_29430.n0 a_22190_29430.n17 1.74185
R7614 a_22190_29430.n24 a_22190_29430.n1 1.74185
R7615 a_22190_29430.n23 a_22190_29430.n22 0.34425
R7616 a_22190_29430.n22 a_22190_29430.n12 0.34425
R7617 a_22190_29430.n16 a_22190_29430.n12 0.34425
R7618 a_22190_29430.n1 a_22190_29430.n0 0.229667
R7619 a_22190_29430.n9 a_22190_29430.n1 0.229667
R7620 a_26300_23070.n2 a_26300_23070.t3 755.889
R7621 a_26300_23070.n1 a_26300_23070.t4 343.034
R7622 a_26300_23070.t0 a_26300_23070.n2 270.334
R7623 a_26300_23070.n1 a_26300_23070.n0 212.733
R7624 a_26300_23070.n0 a_26300_23070.t1 48.0005
R7625 a_26300_23070.n0 a_26300_23070.t2 48.0005
R7626 a_26300_23070.n2 a_26300_23070.n1 35.2005
R7627 a_26300_22300.t4 a_26300_22300.t3 1012.2
R7628 a_26300_22300.n1 a_26300_22300.t1 663.801
R7629 a_26300_22300.t5 a_26300_22300.t6 401.668
R7630 a_26300_22300.n2 a_26300_22300.n0 400.901
R7631 a_26300_22300.n0 a_26300_22300.t2 377.567
R7632 a_26300_22300.n1 a_26300_22300.t4 361.661
R7633 a_26300_22300.t0 a_26300_22300.n2 314.601
R7634 a_26300_22300.n0 a_26300_22300.t5 281.168
R7635 a_26300_22300.n2 a_26300_22300.n1 73.6005
R7636 a_26420_27440.t0 a_26420_27440.t1 96.0005
R7637 a_26390_29930.n0 a_26390_29930.t0 767.801
R7638 a_26390_29930.n1 a_26390_29930.t4 343.949
R7639 a_26390_29930.n0 a_26390_29930.t2 260.733
R7640 a_26390_29930.n2 a_26390_29930.n1 212.733
R7641 a_26390_29930.n1 a_26390_29930.n0 57.6005
R7642 a_26390_29930.t3 a_26390_29930.n2 48.0005
R7643 a_26390_29930.n2 a_26390_29930.t1 48.0005
R7644 a_14140_28370.n2 a_14140_28370.n0 302.507
R7645 a_14140_28370.n10 a_14140_28370.n9 302.163
R7646 a_14140_28370.n8 a_14140_28370.n7 302.163
R7647 a_14140_28370.n6 a_14140_28370.n5 302.163
R7648 a_14140_28370.n4 a_14140_28370.n3 302.163
R7649 a_14140_28370.n2 a_14140_28370.n1 302.163
R7650 a_14140_28370.n11 a_14140_28370.t13 291.503
R7651 a_14140_28370.n14 a_14140_28370.t17 291.288
R7652 a_14140_28370.n13 a_14140_28370.t15 291.288
R7653 a_14140_28370.n12 a_14140_28370.t16 291.288
R7654 a_14140_28370.n11 a_14140_28370.t14 291.288
R7655 a_14140_28370.t0 a_14140_28370.n15 173.233
R7656 a_14140_28370.n9 a_14140_28370.t11 39.4005
R7657 a_14140_28370.n9 a_14140_28370.t3 39.4005
R7658 a_14140_28370.n7 a_14140_28370.t5 39.4005
R7659 a_14140_28370.n7 a_14140_28370.t9 39.4005
R7660 a_14140_28370.n5 a_14140_28370.t2 39.4005
R7661 a_14140_28370.n5 a_14140_28370.t7 39.4005
R7662 a_14140_28370.n3 a_14140_28370.t10 39.4005
R7663 a_14140_28370.n3 a_14140_28370.t4 39.4005
R7664 a_14140_28370.n1 a_14140_28370.t8 39.4005
R7665 a_14140_28370.n1 a_14140_28370.t1 39.4005
R7666 a_14140_28370.n0 a_14140_28370.t6 39.4005
R7667 a_14140_28370.n0 a_14140_28370.t12 39.4005
R7668 a_14140_28370.n15 a_14140_28370.n10 12.0474
R7669 a_14140_28370.n15 a_14140_28370.n14 6.4005
R7670 a_14140_28370.n14 a_14140_28370.n13 0.643357
R7671 a_14140_28370.n12 a_14140_28370.n11 0.643357
R7672 a_14140_28370.n10 a_14140_28370.n8 0.34425
R7673 a_14140_28370.n8 a_14140_28370.n6 0.34425
R7674 a_14140_28370.n6 a_14140_28370.n4 0.34425
R7675 a_14140_28370.n4 a_14140_28370.n2 0.34425
R7676 a_14140_28370.n13 a_14140_28370.n12 0.214786
R7677 a_26390_31270.n0 a_26390_31270.t0 729.933
R7678 a_26390_31270.n1 a_26390_31270.t4 547.134
R7679 a_26390_31270.n0 a_26390_31270.t1 260.733
R7680 a_26390_31270.n2 a_26390_31270.n1 212.733
R7681 a_26390_31270.n1 a_26390_31270.n0 57.6005
R7682 a_26390_31270.n2 a_26390_31270.t2 48.0005
R7683 a_26390_31270.t3 a_26390_31270.n2 48.0005
R7684 a_13370_29270.n134 a_13370_29270.n133 808.569
R7685 a_13370_29270.n81 a_13370_29270.t8 132.74
R7686 a_13370_29270.n133 a_13370_29270.n132 83.7933
R7687 a_13370_29270.n110 a_13370_29270.n11 83.5719
R7688 a_13370_29270.n115 a_13370_29270.n10 83.5719
R7689 a_13370_29270.n122 a_13370_29270.n121 83.5719
R7690 a_13370_29270.n8 a_13370_29270.n5 83.5719
R7691 a_13370_29270.n127 a_13370_29270.n4 83.5719
R7692 a_13370_29270.n103 a_13370_29270.n102 83.5719
R7693 a_13370_29270.n101 a_13370_29270.n100 83.5719
R7694 a_13370_29270.n99 a_13370_29270.n98 83.5719
R7695 a_13370_29270.n93 a_13370_29270.n92 83.5719
R7696 a_13370_29270.n94 a_13370_29270.n25 83.5719
R7697 a_13370_29270.n84 a_13370_29270.n28 83.5719
R7698 a_13370_29270.n76 a_13370_29270.n29 83.5719
R7699 a_13370_29270.n78 a_13370_29270.n77 83.5719
R7700 a_13370_29270.n70 a_13370_29270.n33 83.5719
R7701 a_13370_29270.n60 a_13370_29270.n59 83.5719
R7702 a_13370_29270.n58 a_13370_29270.n57 83.5719
R7703 a_13370_29270.n56 a_13370_29270.n55 83.5719
R7704 a_13370_29270.n1 a_13370_29270.n0 83.5719
R7705 a_13370_29270.n44 a_13370_29270.n43 83.5719
R7706 a_13370_29270.n117 a_13370_29270.n10 73.3165
R7707 a_13370_29270.n129 a_13370_29270.n4 73.3165
R7708 a_13370_29270.n99 a_13370_29270.n17 73.3165
R7709 a_13370_29270.n93 a_13370_29270.n26 73.3165
R7710 a_13370_29270.n77 a_13370_29270.n75 73.3165
R7711 a_13370_29270.n56 a_13370_29270.n40 73.3165
R7712 a_13370_29270.n121 a_13370_29270.n120 73.19
R7713 a_13370_29270.n104 a_13370_29270.n103 73.19
R7714 a_13370_29270.n86 a_13370_29270.n28 73.19
R7715 a_13370_29270.n72 a_13370_29270.n33 73.19
R7716 a_13370_29270.n61 a_13370_29270.n60 73.19
R7717 a_13370_29270.n111 a_13370_29270.t1 65.0331
R7718 a_13370_29270.n95 a_13370_29270.t6 65.0331
R7719 a_13370_29270.n34 a_13370_29270.t3 36.6632
R7720 a_13370_29270.t7 a_13370_29270.n41 36.6632
R7721 a_13370_29270.n110 a_13370_29270.n10 26.074
R7722 a_13370_29270.n8 a_13370_29270.n4 26.074
R7723 a_13370_29270.n101 a_13370_29270.n99 26.074
R7724 a_13370_29270.n94 a_13370_29270.n93 26.074
R7725 a_13370_29270.n77 a_13370_29270.n76 26.074
R7726 a_13370_29270.n58 a_13370_29270.n56 26.074
R7727 a_13370_29270.n43 a_13370_29270.n0 26.074
R7728 a_13370_29270.n133 a_13370_29270.n0 26.074
R7729 a_13370_29270.n121 a_13370_29270.t4 25.7843
R7730 a_13370_29270.n103 a_13370_29270.t5 25.7843
R7731 a_13370_29270.t0 a_13370_29270.n28 25.7843
R7732 a_13370_29270.t3 a_13370_29270.n33 25.7843
R7733 a_13370_29270.n60 a_13370_29270.t2 25.7843
R7734 a_13370_29270.n43 a_13370_29270.t7 25.7843
R7735 a_13370_29270.n50 a_13370_29270.n38 9.3005
R7736 a_13370_29270.n50 a_13370_29270.n36 9.3005
R7737 a_13370_29270.n50 a_13370_29270.n39 9.3005
R7738 a_13370_29270.n65 a_13370_29270.n50 9.3005
R7739 a_13370_29270.n52 a_13370_29270.n38 9.3005
R7740 a_13370_29270.n52 a_13370_29270.n36 9.3005
R7741 a_13370_29270.n52 a_13370_29270.n39 9.3005
R7742 a_13370_29270.n65 a_13370_29270.n52 9.3005
R7743 a_13370_29270.n49 a_13370_29270.n38 9.3005
R7744 a_13370_29270.n49 a_13370_29270.n36 9.3005
R7745 a_13370_29270.n49 a_13370_29270.n39 9.3005
R7746 a_13370_29270.n65 a_13370_29270.n49 9.3005
R7747 a_13370_29270.n64 a_13370_29270.n38 9.3005
R7748 a_13370_29270.n64 a_13370_29270.n36 9.3005
R7749 a_13370_29270.n64 a_13370_29270.n39 9.3005
R7750 a_13370_29270.n65 a_13370_29270.n64 9.3005
R7751 a_13370_29270.n48 a_13370_29270.n38 9.3005
R7752 a_13370_29270.n48 a_13370_29270.n36 9.3005
R7753 a_13370_29270.n48 a_13370_29270.n39 9.3005
R7754 a_13370_29270.n48 a_13370_29270.n35 9.3005
R7755 a_13370_29270.n65 a_13370_29270.n48 9.3005
R7756 a_13370_29270.n66 a_13370_29270.n38 9.3005
R7757 a_13370_29270.n66 a_13370_29270.n36 9.3005
R7758 a_13370_29270.n66 a_13370_29270.n39 9.3005
R7759 a_13370_29270.n66 a_13370_29270.n35 9.3005
R7760 a_13370_29270.n66 a_13370_29270.n65 9.3005
R7761 a_13370_29270.n19 a_13370_29270.n15 9.3005
R7762 a_13370_29270.n19 a_13370_29270.n14 9.3005
R7763 a_13370_29270.n19 a_13370_29270.n16 9.3005
R7764 a_13370_29270.n108 a_13370_29270.n19 9.3005
R7765 a_13370_29270.n21 a_13370_29270.n15 9.3005
R7766 a_13370_29270.n21 a_13370_29270.n14 9.3005
R7767 a_13370_29270.n21 a_13370_29270.n16 9.3005
R7768 a_13370_29270.n108 a_13370_29270.n21 9.3005
R7769 a_13370_29270.n18 a_13370_29270.n15 9.3005
R7770 a_13370_29270.n18 a_13370_29270.n14 9.3005
R7771 a_13370_29270.n18 a_13370_29270.n16 9.3005
R7772 a_13370_29270.n108 a_13370_29270.n18 9.3005
R7773 a_13370_29270.n23 a_13370_29270.n15 9.3005
R7774 a_13370_29270.n23 a_13370_29270.n14 9.3005
R7775 a_13370_29270.n23 a_13370_29270.n16 9.3005
R7776 a_13370_29270.n108 a_13370_29270.n23 9.3005
R7777 a_13370_29270.n109 a_13370_29270.n15 9.3005
R7778 a_13370_29270.n109 a_13370_29270.n14 9.3005
R7779 a_13370_29270.n109 a_13370_29270.n16 9.3005
R7780 a_13370_29270.n109 a_13370_29270.n13 9.3005
R7781 a_13370_29270.n109 a_13370_29270.n108 9.3005
R7782 a_13370_29270.n107 a_13370_29270.n15 9.3005
R7783 a_13370_29270.n107 a_13370_29270.n14 9.3005
R7784 a_13370_29270.n107 a_13370_29270.n16 9.3005
R7785 a_13370_29270.n107 a_13370_29270.n13 9.3005
R7786 a_13370_29270.n108 a_13370_29270.n107 9.3005
R7787 a_13370_29270.n51 a_13370_29270.n35 4.64654
R7788 a_13370_29270.n62 a_13370_29270.n54 4.64654
R7789 a_13370_29270.n53 a_13370_29270.n35 4.64654
R7790 a_13370_29270.n63 a_13370_29270.n62 4.64654
R7791 a_13370_29270.n62 a_13370_29270.n37 4.64654
R7792 a_13370_29270.n20 a_13370_29270.n13 4.64654
R7793 a_13370_29270.n105 a_13370_29270.n97 4.64654
R7794 a_13370_29270.n22 a_13370_29270.n13 4.64654
R7795 a_13370_29270.n105 a_13370_29270.n12 4.64654
R7796 a_13370_29270.n106 a_13370_29270.n105 4.64654
R7797 a_13370_29270.n120 a_13370_29270.n119 2.36206
R7798 a_13370_29270.n87 a_13370_29270.n86 2.36206
R7799 a_13370_29270.n73 a_13370_29270.n72 2.36206
R7800 a_13370_29270.n118 a_13370_29270.n117 2.19742
R7801 a_13370_29270.n130 a_13370_29270.n129 2.19742
R7802 a_13370_29270.n88 a_13370_29270.n26 2.19742
R7803 a_13370_29270.n75 a_13370_29270.n74 2.19742
R7804 a_13370_29270.n69 a_13370_29270.n34 1.80777
R7805 a_13370_29270.n45 a_13370_29270.n41 1.80777
R7806 a_13370_29270.n111 a_13370_29270.n11 1.56484
R7807 a_13370_29270.n95 a_13370_29270.n25 1.56484
R7808 a_13370_29270.n71 a_13370_29270.n32 1.5505
R7809 a_13370_29270.n69 a_13370_29270.n68 1.5505
R7810 a_13370_29270.n85 a_13370_29270.n27 1.5505
R7811 a_13370_29270.n83 a_13370_29270.n82 1.5505
R7812 a_13370_29270.n80 a_13370_29270.n79 1.5505
R7813 a_13370_29270.n31 a_13370_29270.n30 1.5505
R7814 a_13370_29270.n91 a_13370_29270.n24 1.5505
R7815 a_13370_29270.n90 a_13370_29270.n89 1.5505
R7816 a_13370_29270.n7 a_13370_29270.n6 1.5505
R7817 a_13370_29270.n124 a_13370_29270.n123 1.5505
R7818 a_13370_29270.n126 a_13370_29270.n125 1.5505
R7819 a_13370_29270.n128 a_13370_29270.n3 1.5505
R7820 a_13370_29270.n114 a_13370_29270.n113 1.5505
R7821 a_13370_29270.n116 a_13370_29270.n9 1.5505
R7822 a_13370_29270.n132 a_13370_29270.n131 1.5505
R7823 a_13370_29270.n42 a_13370_29270.n2 1.5505
R7824 a_13370_29270.n46 a_13370_29270.n45 1.5505
R7825 a_13370_29270.n132 a_13370_29270.n1 1.43912
R7826 a_13370_29270.n122 a_13370_29270.n7 1.25468
R7827 a_13370_29270.n102 a_13370_29270.n15 1.25468
R7828 a_13370_29270.n85 a_13370_29270.n84 1.25468
R7829 a_13370_29270.n71 a_13370_29270.n70 1.25468
R7830 a_13370_29270.n59 a_13370_29270.n38 1.25468
R7831 a_13370_29270.n44 a_13370_29270.n42 1.25468
R7832 a_13370_29270.n117 a_13370_29270.n116 1.19225
R7833 a_13370_29270.n129 a_13370_29270.n128 1.19225
R7834 a_13370_29270.n17 a_13370_29270.n13 1.19225
R7835 a_13370_29270.n90 a_13370_29270.n26 1.19225
R7836 a_13370_29270.n75 a_13370_29270.n31 1.19225
R7837 a_13370_29270.n40 a_13370_29270.n35 1.19225
R7838 a_13370_29270.n123 a_13370_29270.n5 1.07024
R7839 a_13370_29270.n100 a_13370_29270.n14 1.07024
R7840 a_13370_29270.n83 a_13370_29270.n29 1.07024
R7841 a_13370_29270.n57 a_13370_29270.n36 1.07024
R7842 a_13370_29270.n67 a_13370_29270.n34 1.04793
R7843 a_13370_29270.n47 a_13370_29270.n41 1.04793
R7844 a_13370_29270.n120 a_13370_29270.n7 1.0237
R7845 a_13370_29270.n104 a_13370_29270.n15 1.0237
R7846 a_13370_29270.n86 a_13370_29270.n85 1.0237
R7847 a_13370_29270.n72 a_13370_29270.n71 1.0237
R7848 a_13370_29270.n61 a_13370_29270.n38 1.0237
R7849 a_13370_29270.n116 a_13370_29270.n115 0.959578
R7850 a_13370_29270.n128 a_13370_29270.n127 0.959578
R7851 a_13370_29270.n98 a_13370_29270.n13 0.959578
R7852 a_13370_29270.n92 a_13370_29270.n90 0.959578
R7853 a_13370_29270.n78 a_13370_29270.n31 0.959578
R7854 a_13370_29270.n55 a_13370_29270.n35 0.959578
R7855 a_13370_29270.n115 a_13370_29270.n114 0.885803
R7856 a_13370_29270.n127 a_13370_29270.n126 0.885803
R7857 a_13370_29270.n98 a_13370_29270.n16 0.885803
R7858 a_13370_29270.n92 a_13370_29270.n91 0.885803
R7859 a_13370_29270.n79 a_13370_29270.n78 0.885803
R7860 a_13370_29270.n55 a_13370_29270.n39 0.885803
R7861 a_13370_29270.n105 a_13370_29270.n104 0.812055
R7862 a_13370_29270.n62 a_13370_29270.n61 0.812055
R7863 a_13370_29270.n114 a_13370_29270.n11 0.77514
R7864 a_13370_29270.n126 a_13370_29270.n5 0.77514
R7865 a_13370_29270.n100 a_13370_29270.n16 0.77514
R7866 a_13370_29270.n91 a_13370_29270.n25 0.77514
R7867 a_13370_29270.n79 a_13370_29270.n29 0.77514
R7868 a_13370_29270.n57 a_13370_29270.n39 0.77514
R7869 a_13370_29270.n108 a_13370_29270.n17 0.647417
R7870 a_13370_29270.n65 a_13370_29270.n40 0.647417
R7871 a_13370_29270.n123 a_13370_29270.n122 0.590702
R7872 a_13370_29270.n102 a_13370_29270.n14 0.590702
R7873 a_13370_29270.n84 a_13370_29270.n83 0.590702
R7874 a_13370_29270.n70 a_13370_29270.n69 0.590702
R7875 a_13370_29270.n59 a_13370_29270.n36 0.590702
R7876 a_13370_29270.n45 a_13370_29270.n44 0.590702
R7877 a_13370_29270.n96 a_13370_29270.n95 0.531214
R7878 a_13370_29270.n112 a_13370_29270.n111 0.531214
R7879 a_13370_29270.n42 a_13370_29270.n1 0.406264
R7880 a_13370_29270.t1 a_13370_29270.n110 0.290206
R7881 a_13370_29270.t4 a_13370_29270.n8 0.290206
R7882 a_13370_29270.t5 a_13370_29270.n101 0.290206
R7883 a_13370_29270.t6 a_13370_29270.n94 0.290206
R7884 a_13370_29270.n76 a_13370_29270.t0 0.290206
R7885 a_13370_29270.t2 a_13370_29270.n58 0.290206
R7886 a_13370_29270.n74 a_13370_29270.n73 0.154071
R7887 a_13370_29270.n88 a_13370_29270.n87 0.154071
R7888 a_13370_29270.n131 a_13370_29270.n130 0.154071
R7889 a_13370_29270.n119 a_13370_29270.n118 0.154071
R7890 a_13370_29270.n67 a_13370_29270.n66 0.137464
R7891 a_13370_29270.n107 a_13370_29270.n96 0.137464
R7892 a_13370_29270.n48 a_13370_29270.n47 0.134964
R7893 a_13370_29270.n112 a_13370_29270.n109 0.134964
R7894 a_13370_29270.n68 a_13370_29270.n32 0.0183571
R7895 a_13370_29270.n73 a_13370_29270.n32 0.0183571
R7896 a_13370_29270.n74 a_13370_29270.n30 0.0183571
R7897 a_13370_29270.n80 a_13370_29270.n30 0.0183571
R7898 a_13370_29270.n82 a_13370_29270.n27 0.0183571
R7899 a_13370_29270.n87 a_13370_29270.n27 0.0183571
R7900 a_13370_29270.n89 a_13370_29270.n88 0.0183571
R7901 a_13370_29270.n89 a_13370_29270.n24 0.0183571
R7902 a_13370_29270.n46 a_13370_29270.n2 0.0183571
R7903 a_13370_29270.n131 a_13370_29270.n2 0.0183571
R7904 a_13370_29270.n130 a_13370_29270.n3 0.0183571
R7905 a_13370_29270.n125 a_13370_29270.n3 0.0183571
R7906 a_13370_29270.n125 a_13370_29270.n124 0.0183571
R7907 a_13370_29270.n124 a_13370_29270.n6 0.0183571
R7908 a_13370_29270.n119 a_13370_29270.n6 0.0183571
R7909 a_13370_29270.n118 a_13370_29270.n9 0.0183571
R7910 a_13370_29270.n113 a_13370_29270.n9 0.0183571
R7911 a_13370_29270.n68 a_13370_29270.n67 0.0106786
R7912 a_13370_29270.n82 a_13370_29270.n81 0.0106786
R7913 a_13370_29270.n47 a_13370_29270.n46 0.0106786
R7914 a_13370_29270.n66 a_13370_29270.n37 0.00992001
R7915 a_13370_29270.n52 a_13370_29270.n51 0.00992001
R7916 a_13370_29270.n54 a_13370_29270.n49 0.00992001
R7917 a_13370_29270.n64 a_13370_29270.n53 0.00992001
R7918 a_13370_29270.n63 a_13370_29270.n48 0.00992001
R7919 a_13370_29270.n50 a_13370_29270.n37 0.00992001
R7920 a_13370_29270.n51 a_13370_29270.n50 0.00992001
R7921 a_13370_29270.n54 a_13370_29270.n52 0.00992001
R7922 a_13370_29270.n53 a_13370_29270.n49 0.00992001
R7923 a_13370_29270.n64 a_13370_29270.n63 0.00992001
R7924 a_13370_29270.n107 a_13370_29270.n106 0.00992001
R7925 a_13370_29270.n21 a_13370_29270.n20 0.00992001
R7926 a_13370_29270.n97 a_13370_29270.n18 0.00992001
R7927 a_13370_29270.n23 a_13370_29270.n22 0.00992001
R7928 a_13370_29270.n109 a_13370_29270.n12 0.00992001
R7929 a_13370_29270.n106 a_13370_29270.n19 0.00992001
R7930 a_13370_29270.n20 a_13370_29270.n19 0.00992001
R7931 a_13370_29270.n97 a_13370_29270.n21 0.00992001
R7932 a_13370_29270.n22 a_13370_29270.n18 0.00992001
R7933 a_13370_29270.n23 a_13370_29270.n12 0.00992001
R7934 a_13370_29270.n81 a_13370_29270.n80 0.00817857
R7935 a_13370_29270.n96 a_13370_29270.n24 0.00817857
R7936 a_13370_29270.n113 a_13370_29270.n112 0.00817857
R7937 a_24280_31990.n3 a_24280_31990.t7 796.295
R7938 a_24280_31990.n1 a_24280_31990.t0 761.4
R7939 a_24280_31990.n4 a_24280_31990.n3 631.564
R7940 a_24280_31990.n0 a_24280_31990.t2 538.234
R7941 a_24280_31990.t7 a_24280_31990.t5 514.134
R7942 a_24280_31990.n1 a_24280_31990.n0 435.952
R7943 a_24280_31990.n2 a_24280_31990.t4 313.3
R7944 a_24280_31990.n0 a_24280_31990.t3 297.233
R7945 a_24280_31990.t1 a_24280_31990.n4 233
R7946 a_24280_31990.n2 a_24280_31990.t6 200.833
R7947 a_24280_31990.n3 a_24280_31990.n2 160.667
R7948 a_24280_31990.n4 a_24280_31990.n1 46.7205
R7949 a_26640_21160.t1 a_26640_21160.n0 708.125
R7950 a_26640_21160.t1 a_26640_21160.n1 708.125
R7951 a_26640_21160.n1 a_26640_21160.t2 410.519
R7952 a_26640_21160.n0 a_26640_21160.t0 305.649
R7953 a_26640_21160.n1 a_26640_21160.n0 21.3338
R7954 a_24280_27770.n0 a_24280_27770.t3 1004.17
R7955 a_24280_27770.n2 a_24280_27770.n1 545.634
R7956 a_24280_27770.t0 a_24280_27770.n3 458.818
R7957 a_24280_27770.t0 a_24280_27770.n3 429.281
R7958 a_24280_27770.n1 a_24280_27770.t5 425.767
R7959 a_24280_27770.n1 a_24280_27770.n0 417.733
R7960 a_24280_27770.n0 a_24280_27770.t2 409.7
R7961 a_24280_27770.n1 a_24280_27770.t4 409.7
R7962 a_24280_27770.n2 a_24280_27770.t1 173.095
R7963 a_24280_27770.n3 a_24280_27770.n2 36.568
R7964 a_24310_27670.t2 a_24310_27670.n4 458.818
R7965 a_24310_27670.t2 a_24310_27670.n4 429.281
R7966 a_24310_27670.t5 a_24310_27670.t3 377.567
R7967 a_24310_27670.n0 a_24310_27670.t4 326.658
R7968 a_24310_27670.n2 a_24310_27670.n1 252.345
R7969 a_24310_27670.n1 a_24310_27670.n0 196.817
R7970 a_24310_27670.n3 a_24310_27670.t0 164.775
R7971 a_24310_27670.n2 a_24310_27670.t1 164.775
R7972 a_24310_27670.n3 a_24310_27670.n2 112.001
R7973 a_24310_27670.n1 a_24310_27670.t5 92.3838
R7974 a_24310_27670.t3 a_24310_27670.n0 92.3838
R7975 a_24310_27670.n4 a_24310_27670.n3 60.248
R7976 a_23130_29200.t1 a_23130_29200.n2 500.086
R7977 a_23130_29200.n0 a_23130_29200.t2 490.034
R7978 a_23130_29200.t1 a_23130_29200.n2 461.389
R7979 a_23130_29200.n1 a_23130_29200.n0 368.524
R7980 a_23130_29200.n0 a_23130_29200.t3 345.433
R7981 a_23130_29200.n1 a_23130_29200.t0 177.577
R7982 a_23130_29200.n2 a_23130_29200.n1 48.3899
R7983 a_24280_29730.t1 a_24280_29730.n2 500.086
R7984 a_24280_29730.n0 a_24280_29730.t2 490.034
R7985 a_24280_29730.t1 a_24280_29730.n2 461.389
R7986 a_24280_29730.n1 a_24280_29730.n0 449.233
R7987 a_24280_29730.n0 a_24280_29730.t3 345.433
R7988 a_24280_29730.n1 a_24280_29730.t0 177.577
R7989 a_24280_29730.n2 a_24280_29730.n1 48.3899
R7990 a_26300_24370.n0 a_26300_24370.t1 755.889
R7991 a_26300_24370.n1 a_26300_24370.t4 343.034
R7992 a_26300_24370.n0 a_26300_24370.t2 270.334
R7993 a_26300_24370.n2 a_26300_24370.n1 212.733
R7994 a_26300_24370.n2 a_26300_24370.t3 48.0005
R7995 a_26300_24370.t0 a_26300_24370.n2 48.0005
R7996 a_26300_24370.n1 a_26300_24370.n0 35.2005
R7997 a_26300_23600.t4 a_26300_23600.t3 1012.2
R7998 a_26300_23600.n1 a_26300_23600.t0 663.801
R7999 a_26300_23600.t5 a_26300_23600.t6 401.668
R8000 a_26300_23600.n2 a_26300_23600.n0 400.901
R8001 a_26300_23600.n0 a_26300_23600.t2 377.567
R8002 a_26300_23600.n1 a_26300_23600.t4 361.661
R8003 a_26300_23600.t1 a_26300_23600.n2 314.601
R8004 a_26300_23600.n0 a_26300_23600.t5 281.168
R8005 a_26300_23600.n2 a_26300_23600.n1 73.6005
R8006 a_26390_30500.n0 a_26390_30500.t1 719.801
R8007 a_26390_30500.t3 a_26390_30500.t2 514.134
R8008 a_26390_30500.n0 a_26390_30500.t3 332.783
R8009 a_26390_30500.t0 a_26390_30500.n0 330.601
R8010 a_26420_30420.t0 a_26420_30420.n0 531.067
R8011 a_26420_30420.n0 a_26420_30420.t1 48.0005
R8012 a_26420_30420.n0 a_26420_30420.t2 48.0005
R8013 ua[1].n3 ua[1].n1 409.7
R8014 ua[1].t4 ua[1].t6 401.668
R8015 ua[1].n1 ua[1].t3 377.567
R8016 ua[1].n0 ua[1].t1 372.118
R8017 ua[1].n1 ua[1].t4 281.168
R8018 ua[1].n2 ua[1].t5 249.034
R8019 ua[1].n0 ua[1].t0 247.934
R8020 ua[1].n3 ua[1].n2 200.833
R8021 ua[1].n4 ua[1].n3 171.457
R8022 ua[1].n2 ua[1].t2 168.701
R8023 ua[1].n4 ua[1].n0 65.3005
R8024 ua[1] ua[1].n4 18.0284
R8025 a_26400_21130.n1 a_26400_21130.n0 413.634
R8026 a_26400_21130.t0 a_26400_21130.n1 372.118
R8027 a_26400_21130.n0 a_26400_21130.t2 249.034
R8028 a_26400_21130.n1 a_26400_21130.t1 247.934
R8029 a_26400_21130.n0 a_26400_21130.t3 168.701
R8030 a_26420_27220.n0 a_26420_27220.t1 691.534
R8031 a_26420_27220.n1 a_26420_27220.t2 663.801
R8032 a_26420_27220.n0 a_26420_27220.t3 527.867
R8033 a_26420_27220.t0 a_26420_27220.n1 372.2
R8034 a_26420_27220.n1 a_26420_27220.n0 85.3338
R8035 a_26390_32300.n0 a_26390_32300.t0 767.801
R8036 a_26390_32300.n1 a_26390_32300.t4 343.034
R8037 a_26390_32300.n0 a_26390_32300.t1 260.733
R8038 a_26390_32300.n2 a_26390_32300.n1 212.733
R8039 a_26390_32300.n1 a_26390_32300.n0 57.6005
R8040 a_26390_32300.n2 a_26390_32300.t2 48.0005
R8041 a_26390_32300.t3 a_26390_32300.n2 48.0005
R8042 ua[0] ua[0].n0 546.412
R8043 ua[0].n0 ua[0].t0 538.234
R8044 ua[0].n0 ua[0].t1 297.233
R8045 a_23550_31910.t0 a_23550_31910.t1 39.4005
R8046 a_26300_24900.t4 a_26300_24900.t2 1012.2
R8047 a_26300_24900.n1 a_26300_24900.t1 663.801
R8048 a_26300_24900.t5 a_26300_24900.t6 401.668
R8049 a_26300_24900.n2 a_26300_24900.n0 400.901
R8050 a_26300_24900.n1 a_26300_24900.t4 361.661
R8051 a_26300_24900.t0 a_26300_24900.n2 314.601
R8052 a_26300_24900.n0 a_26300_24900.t5 281.168
R8053 a_26300_24900.n0 a_26300_24900.t3 232.968
R8054 a_26300_24900.n2 a_26300_24900.n1 73.6005
R8055 a_24310_30490.t0 a_24310_30490.t1 39.4005
R8056 a_24280_30980.n1 a_24280_30980.t3 517.347
R8057 a_24280_30980.n2 a_24280_30980.n1 417.574
R8058 a_24280_30980.n2 a_24280_30980.n0 244.716
R8059 a_24280_30980.n1 a_24280_30980.t4 228.148
R8060 a_24280_30980.t1 a_24280_30980.n2 221.411
R8061 a_24280_30980.n0 a_24280_30980.t0 24.0005
R8062 a_24280_30980.n0 a_24280_30980.t2 24.0005
R8063 a_26400_20530.n1 a_26400_20530.n0 413.634
R8064 a_26400_20530.t1 a_26400_20530.n1 372.118
R8065 a_26400_20530.n0 a_26400_20530.t2 249.034
R8066 a_26400_20530.n1 a_26400_20530.t0 247.934
R8067 a_26400_20530.n0 a_26400_20530.t3 168.701
R8068 a_26640_20560.t1 a_26640_20560.n0 708.125
R8069 a_26640_20560.t1 a_26640_20560.n1 708.125
R8070 a_26640_20560.n1 a_26640_20560.t2 410.519
R8071 a_26640_20560.n0 a_26640_20560.t0 305.649
R8072 a_26640_20560.n1 a_26640_20560.n0 21.3338
R8073 a_26740_30530.t0 a_26740_30530.t1 157.601
R8074 a_23020_31090.n2 a_23020_31090.n0 1295.28
R8075 a_23020_31090.t4 a_23020_31090.t6 1188.93
R8076 a_23020_31090.t6 a_23020_31090.t5 835.467
R8077 a_23020_31090.n0 a_23020_31090.t3 586.433
R8078 a_23020_31090.n0 a_23020_31090.t4 249.034
R8079 a_23020_31090.n2 a_23020_31090.n1 247.917
R8080 a_23020_31090.t2 a_23020_31090.n2 221.411
R8081 a_23020_31090.n1 a_23020_31090.t0 24.0005
R8082 a_23020_31090.n1 a_23020_31090.t1 24.0005
R8083 a_26300_22410.n4 a_26300_22410.t1 758.734
R8084 a_26300_22410.t2 a_26300_22410.n5 758.734
R8085 a_26300_22410.n0 a_26300_22410.t4 538.234
R8086 a_26300_22410.n3 a_26300_22410.n2 342.757
R8087 a_26300_22410.n5 a_26300_22410.t0 260.733
R8088 a_26300_22410.n3 a_26300_22410.t6 190.123
R8089 a_26300_22410.n4 a_26300_22410.n3 180.8
R8090 a_26300_22410.n0 a_26300_22410.t5 136.567
R8091 a_26300_22410.n1 a_26300_22410.t3 136.567
R8092 a_26300_22410.n2 a_26300_22410.t7 136.567
R8093 a_26300_22410.n1 a_26300_22410.n0 128.534
R8094 a_26300_22410.n2 a_26300_22410.n1 128.534
R8095 a_26300_22410.n5 a_26300_22410.n4 57.6005
R8096 a_26390_26970.n2 a_26390_26970.t3 727.09
R8097 a_26390_26970.n1 a_26390_26970.t4 343.949
R8098 a_26390_26970.t2 a_26390_26970.n2 270.334
R8099 a_26390_26970.n1 a_26390_26970.n0 212.733
R8100 a_26390_26970.n0 a_26390_26970.t0 48.0005
R8101 a_26390_26970.n0 a_26390_26970.t1 48.0005
R8102 a_26390_26970.n2 a_26390_26970.n1 35.2005
R8103 a_25350_8708.t1 a_25350_8708.t0 127.201
R8104 a_13742_34050.t0 a_13742_34050.t12 178.589
R8105 a_13742_34050.t13 a_13742_34050.t6 0.1603
R8106 a_13742_34050.t7 a_13742_34050.t13 0.1603
R8107 a_13742_34050.t15 a_13742_34050.t7 0.1603
R8108 a_13742_34050.t19 a_13742_34050.t15 0.1603
R8109 a_13742_34050.t2 a_13742_34050.t19 0.1603
R8110 a_13742_34050.t20 a_13742_34050.t2 0.1603
R8111 a_13742_34050.t4 a_13742_34050.t20 0.1603
R8112 a_13742_34050.t10 a_13742_34050.t4 0.1603
R8113 a_13742_34050.t9 a_13742_34050.t16 0.1603
R8114 a_13742_34050.t3 a_13742_34050.t9 0.1603
R8115 a_13742_34050.t8 a_13742_34050.t3 0.1603
R8116 a_13742_34050.t1 a_13742_34050.t8 0.1603
R8117 a_13742_34050.t18 a_13742_34050.t1 0.1603
R8118 a_13742_34050.t14 a_13742_34050.t18 0.1603
R8119 a_13742_34050.t17 a_13742_34050.t14 0.1603
R8120 a_13742_34050.t12 a_13742_34050.t17 0.1603
R8121 a_13742_34050.t11 a_13742_34050.n0 0.159278
R8122 a_13742_34050.t16 a_13742_34050.t11 0.137822
R8123 a_13742_34050.n0 a_13742_34050.t10 0.1368
R8124 a_13742_34050.n0 a_13742_34050.t5 0.00152174
R8125 a_23020_29890.t4 a_23020_29890.t3 835.467
R8126 a_23020_29890.n0 a_23020_29890.t7 517.347
R8127 a_23020_29890.n1 a_23020_29890.t5 490.034
R8128 a_23020_29890.n2 a_23020_29890.n1 429.932
R8129 a_23020_29890.n2 a_23020_29890.t4 394.267
R8130 a_23020_29890.n1 a_23020_29890.t6 345.433
R8131 a_23020_29890.n5 a_23020_29890.n4 244.715
R8132 a_23020_29890.n0 a_23020_29890.t8 228.148
R8133 a_23020_29890.t2 a_23020_29890.n5 221.411
R8134 a_23020_29890.n3 a_23020_29890.n0 209.601
R8135 a_23020_29890.n5 a_23020_29890.n3 207.974
R8136 a_23020_29890.n3 a_23020_29890.n2 123.35
R8137 a_23020_29890.n4 a_23020_29890.t1 24.0005
R8138 a_23020_29890.n4 a_23020_29890.t0 24.0005
R8139 a_23130_29970.t0 a_23130_29970.t1 48.0005
R8140 a_26300_23710.n4 a_26300_23710.t1 758.734
R8141 a_26300_23710.t2 a_26300_23710.n5 758.734
R8142 a_26300_23710.n0 a_26300_23710.t4 538.234
R8143 a_26300_23710.n3 a_26300_23710.n2 342.757
R8144 a_26300_23710.n5 a_26300_23710.t0 260.733
R8145 a_26300_23710.n3 a_26300_23710.t6 190.123
R8146 a_26300_23710.n4 a_26300_23710.n3 180.8
R8147 a_26300_23710.n0 a_26300_23710.t5 136.567
R8148 a_26300_23710.n1 a_26300_23710.t3 136.567
R8149 a_26300_23710.n2 a_26300_23710.t7 136.567
R8150 a_26300_23710.n1 a_26300_23710.n0 128.534
R8151 a_26300_23710.n2 a_26300_23710.n1 128.534
R8152 a_26300_23710.n5 a_26300_23710.n4 57.6005
R8153 a_13532_33810.t0 a_13532_33810.t1 258.591
R8154 a_14610_33690.t0 a_14610_33690.t1 258.591
R8155 a_24310_31910.t0 a_24310_31910.t1 39.4005
R8156 a_24310_27960.n0 a_24310_27960.t3 605.311
R8157 a_24310_27960.t1 a_24310_27960.n1 458.818
R8158 a_24310_27960.t1 a_24310_27960.n1 429.281
R8159 a_24310_27960.t3 a_24310_27960.t2 423.983
R8160 a_24310_27960.n0 a_24310_27960.t0 148.775
R8161 a_24310_27960.n1 a_24310_27960.n0 65.048
R8162 a_26390_29240.t2 a_26390_29240.n2 749.134
R8163 a_26390_29240.n2 a_26390_29240.t1 691.534
R8164 a_26390_29240.n1 a_26390_29240.n0 359.233
R8165 a_26390_29240.n1 a_26390_29240.t0 346.601
R8166 a_26390_29240.n0 a_26390_29240.t3 345.433
R8167 a_26390_29240.n0 a_26390_29240.t4 168.701
R8168 a_26390_29240.n2 a_26390_29240.n1 6.4005
R8169 a_19940_24230.t2 a_19940_24230.n6 1026.49
R8170 a_19940_24230.n3 a_19940_24230.n2 398.401
R8171 a_19940_24230.n2 a_19940_24230.n0 328.447
R8172 a_19940_24230.n2 a_19940_24230.n1 322.601
R8173 a_19940_24230.n4 a_19940_24230.t8 313.3
R8174 a_19940_24230.n5 a_19940_24230.t5 313.3
R8175 a_19940_24230.n6 a_19940_24230.t6 313.3
R8176 a_19940_24230.n3 a_19940_24230.t7 232.968
R8177 a_19940_24230.n4 a_19940_24230.n3 175.73
R8178 a_19940_24230.n5 a_19940_24230.n4 160.667
R8179 a_19940_24230.n6 a_19940_24230.n5 160.667
R8180 a_19940_24230.n1 a_19940_24230.t4 60.0005
R8181 a_19940_24230.n1 a_19940_24230.t3 60.0005
R8182 a_19940_24230.n0 a_19940_24230.t1 49.2505
R8183 a_19940_24230.n0 a_19940_24230.t0 49.2505
R8184 a_23550_31390.t0 a_23550_31390.t1 39.4005
R8185 a_26420_27330.t0 a_26420_27330.t1 96.0005
R8186 a_14610_33930.n6 a_14610_33930.t10 287.764
R8187 a_14610_33930.n5 a_14610_33930.t8 287.764
R8188 a_14610_33930.n5 a_14610_33930.t7 287.591
R8189 a_14610_33930.n8 a_14610_33930.t11 287.012
R8190 a_14610_33930.n7 a_14610_33930.t9 287.012
R8191 a_14610_33930.t0 a_14610_33930.n9 155.326
R8192 a_14610_33930.n2 a_14610_33930.n0 107.266
R8193 a_14610_33930.n4 a_14610_33930.n3 105.016
R8194 a_14610_33930.n2 a_14610_33930.n1 105.016
R8195 a_14610_33930.n3 a_14610_33930.t6 13.1338
R8196 a_14610_33930.n3 a_14610_33930.t4 13.1338
R8197 a_14610_33930.n1 a_14610_33930.t2 13.1338
R8198 a_14610_33930.n1 a_14610_33930.t3 13.1338
R8199 a_14610_33930.n0 a_14610_33930.t1 13.1338
R8200 a_14610_33930.n0 a_14610_33930.t5 13.1338
R8201 a_14610_33930.n9 a_14610_33930.n4 9.0005
R8202 a_14610_33930.n9 a_14610_33930.n8 6.78086
R8203 a_14610_33930.n4 a_14610_33930.n2 2.2505
R8204 a_14610_33930.n7 a_14610_33930.n6 0.579071
R8205 a_14610_33930.n8 a_14610_33930.n7 0.282643
R8206 a_14610_33930.n6 a_14610_33930.n5 0.2755
R8207 a_26420_29270.t0 a_26420_29270.t1 96.0005
R8208 a_26330_22330.t0 a_26330_22330.t1 96.0005
R8209 a_26390_27410.n1 a_26390_27410.t0 691
R8210 a_26390_27410.n1 a_26390_27410.n0 674.168
R8211 a_26390_27410.n0 a_26390_27410.t2 345.433
R8212 a_26390_27410.t1 a_26390_27410.n1 330.601
R8213 a_26390_27410.n0 a_26390_27410.t3 168.701
R8214 a_26420_29380.n0 a_26420_29380.t0 663.801
R8215 a_26420_29380.t1 a_26420_29380.n0 406.334
R8216 a_26420_29380.n0 a_26420_29380.t2 348.851
R8217 a_26330_23630.t0 a_26330_23630.t1 96.0005
R8218 a_26330_22440.n0 a_26330_22440.t1 713.933
R8219 a_26330_22440.t0 a_26330_22440.n0 337
R8220 a_26330_22440.n0 a_26330_22440.t2 314.233
R8221 a_23130_27960.n0 a_23130_27960.t0 496.889
R8222 a_23130_27960.t2 a_23130_27960.n2 458.818
R8223 a_23130_27960.t2 a_23130_27960.n2 429.281
R8224 a_23130_27960.n0 a_23130_27960.t3 393.634
R8225 a_23130_27960.n1 a_23130_27960.n0 384.967
R8226 a_23130_27960.n1 a_23130_27960.t1 177.576
R8227 a_23130_27960.n2 a_23130_27960.n1 34.648
R8228 a_26330_24930.t0 a_26330_24930.t1 96.0005
R8229 a_26330_23740.n0 a_26330_23740.t1 713.933
R8230 a_26330_23740.t0 a_26330_23740.n0 337
R8231 a_26330_23740.n0 a_26330_23740.t2 314.233
R8232 a_18460_22530.t1 a_18460_22530.t0 286.111
R8233 a_21386_22530.t0 a_21386_22530.t1 364.192
R8234 a_26420_31640.t0 a_26420_31640.t1 96.0005
R8235 a_23100_28450.t1 a_23100_28450.n2 458.818
R8236 a_23100_28450.n0 a_23100_28450.t2 441.834
R8237 a_23100_28450.t1 a_23100_28450.n2 429.281
R8238 a_23100_28450.n0 a_23100_28450.t3 313.3
R8239 a_23100_28450.n1 a_23100_28450.n0 228.8
R8240 a_23100_28450.n1 a_23100_28450.t0 174.375
R8241 a_23100_28450.n2 a_23100_28450.n1 50.648
R8242 a_23550_31010.t0 a_23550_31010.t1 39.4005
R8243 a_26330_25040.n0 a_26330_25040.t0 713.933
R8244 a_26330_25040.t1 a_26330_25040.n0 337
R8245 a_26330_25040.n0 a_26330_25040.t2 314.233
R8246 a_26420_31750.n0 a_26420_31750.t0 663.801
R8247 a_26420_31750.t1 a_26420_31750.n0 406.334
R8248 a_26420_31750.n0 a_26420_31750.t2 355.378
R8249 a_26420_30310.t0 a_26420_30310.t1 96.0005
R8250 a_25860_20560.n0 a_25860_20560.t1 284.2
R8251 a_25860_20560.n0 a_25860_20560.t2 233
R8252 a_25860_20560.t0 a_25860_20560.n0 184.191
R8253 a_24310_28480.t1 a_24310_28480.n2 458.818
R8254 a_24310_28480.t1 a_24310_28480.n2 429.281
R8255 a_24310_28480.n0 a_24310_28480.t2 256.428
R8256 a_24310_28480.n1 a_24310_28480.t0 190.375
R8257 a_24310_28480.n0 a_24310_28480.t3 190.375
R8258 a_24310_28480.n1 a_24310_28480.n0 70.4005
R8259 a_24310_28480.n2 a_24310_28480.n1 34.648
R8260 a_13382_33380.t0 a_13382_33380.t1 258.591
R8261 a_17540_28930.t0 a_17540_28930.t1 178.194
R8262 a_25860_21160.n0 a_25860_21160.t2 284.2
R8263 a_25860_21160.n0 a_25860_21160.t1 233
R8264 a_25860_21160.t0 a_25860_21160.n0 184.191
R8265 a_13382_28490.t0 a_13382_28490.t1 258.591
R8266 a_14990_28610.t0 a_14990_28610.t1 258.591
R8267 a_14990_33260.t0 a_14990_33260.t1 258.591
C0 ua[1] VDPWR 0.708002f
C1 VDPWR ua[0] 0.410436f
C2 VGND VDPWR 10.4345f
C3 VGND 0 20.36459f
C4 ua[1] 0 11.0531f
C5 ua[0] 0 17.6488f
C6 VDPWR 0 0.146274p
C7 a_23130_27960.t1 0 0.026996f
C8 a_23130_27960.t0 0 2.01377f
C9 a_23130_27960.t3 0 0.010471f
C10 a_23130_27960.n0 0 0.029667f
C11 a_23130_27960.n1 0 0.037413f
C12 a_23130_27960.n2 0 0.046542f
C13 a_23130_27960.t2 0 0.03514f
C14 a_14610_33930.t1 0 0.10095f
C15 a_14610_33930.t5 0 0.10095f
C16 a_14610_33930.n0 0 0.2816f
C17 a_14610_33930.t2 0 0.10095f
C18 a_14610_33930.t3 0 0.10095f
C19 a_14610_33930.n1 0 0.253459f
C20 a_14610_33930.n2 0 3.1126f
C21 a_14610_33930.t6 0 0.10095f
C22 a_14610_33930.t4 0 0.10095f
C23 a_14610_33930.n3 0 0.253459f
C24 a_14610_33930.n4 0 2.34993f
C25 a_14610_33930.t7 0 0.055705f
C26 a_14610_33930.t8 0 0.05457f
C27 a_14610_33930.n5 0 0.425181f
C28 a_14610_33930.t10 0 0.05457f
C29 a_14610_33930.n6 0 0.226996f
C30 a_14610_33930.t9 0 0.055305f
C31 a_14610_33930.n7 0 0.228617f
C32 a_14610_33930.t11 0 0.055305f
C33 a_14610_33930.n8 0 0.780841f
C34 a_14610_33930.n9 0 4.14023f
C35 a_14610_33930.t0 0 0.365925f
C36 a_13742_34050.t6 0 0.293845f
C37 a_13742_34050.t13 0 0.309615f
C38 a_13742_34050.t7 0 0.309615f
C39 a_13742_34050.t15 0 0.309615f
C40 a_13742_34050.t19 0 0.309615f
C41 a_13742_34050.t2 0 0.309615f
C42 a_13742_34050.t20 0 0.309615f
C43 a_13742_34050.t4 0 0.309615f
C44 a_13742_34050.t10 0 0.29491f
C45 a_13742_34050.t5 0 0.14206f
C46 a_13742_34050.n0 0 0.183237f
C47 a_13742_34050.t11 0 0.322105f
C48 a_13742_34050.t16 0 0.296149f
C49 a_13742_34050.t9 0 0.309615f
C50 a_13742_34050.t3 0 0.309615f
C51 a_13742_34050.t8 0 0.309615f
C52 a_13742_34050.t1 0 0.309615f
C53 a_13742_34050.t18 0 0.309615f
C54 a_13742_34050.t14 0 0.309615f
C55 a_13742_34050.t17 0 0.309615f
C56 a_13742_34050.t12 0 1.1782f
C57 a_13742_34050.t0 0 0.154879f
C58 a_25350_8708.t0 0 2.39855f
C59 a_14140_28370.t6 0 0.021628f
C60 a_14140_28370.t12 0 0.021628f
C61 a_14140_28370.n0 0 0.047663f
C62 a_14140_28370.t8 0 0.021628f
C63 a_14140_28370.t1 0 0.021628f
C64 a_14140_28370.n1 0 0.047367f
C65 a_14140_28370.n2 0 0.55165f
C66 a_14140_28370.t10 0 0.021628f
C67 a_14140_28370.t4 0 0.021628f
C68 a_14140_28370.n3 0 0.047367f
C69 a_14140_28370.n4 0 0.291113f
C70 a_14140_28370.t2 0 0.021628f
C71 a_14140_28370.t7 0 0.021628f
C72 a_14140_28370.n5 0 0.047367f
C73 a_14140_28370.n6 0 0.291113f
C74 a_14140_28370.t5 0 0.021628f
C75 a_14140_28370.t9 0 0.021628f
C76 a_14140_28370.n7 0 0.047367f
C77 a_14140_28370.n8 0 0.291113f
C78 a_14140_28370.t11 0 0.021628f
C79 a_14140_28370.t3 0 0.021628f
C80 a_14140_28370.n9 0 0.047367f
C81 a_14140_28370.n10 0 1.14445f
C82 a_14140_28370.t13 0 0.033253f
C83 a_14140_28370.t14 0 0.033188f
C84 a_14140_28370.n11 0 0.233433f
C85 a_14140_28370.t16 0 0.033188f
C86 a_14140_28370.n12 0 0.145136f
C87 a_14140_28370.t15 0 0.033188f
C88 a_14140_28370.n13 0 0.145136f
C89 a_14140_28370.t17 0 0.033188f
C90 a_14140_28370.n14 0 0.4804f
C91 a_14140_28370.n15 0 5.4833f
C92 a_14140_28370.t0 0 0.533116f
C93 a_22190_29430.n0 0 0.156934f
C94 a_22190_29430.n1 0 0.118238f
C95 a_22190_29430.t0 0 0.029882f
C96 a_22190_29430.t15 0 0.031397f
C97 a_22190_29430.n2 0 0.067221f
C98 a_22190_29430.t14 0 0.010639f
C99 a_22190_29430.t12 0 0.010639f
C100 a_22190_29430.n3 0 0.041426f
C101 a_22190_29430.t13 0 0.049455f
C102 a_22190_29430.t19 0 0.062085f
C103 a_22190_29430.t18 0 0.04628f
C104 a_22190_29430.n4 0 0.046455f
C105 a_22190_29430.n5 0 0.048543f
C106 a_22190_29430.t11 0 0.03365f
C107 a_22190_29430.n6 0 0.040235f
C108 a_22190_29430.n7 0 0.04416f
C109 a_22190_29430.n8 0 1.61807f
C110 a_22190_29430.n9 0 1.98317f
C111 a_22190_29430.n11 0 0.060082f
C112 a_22190_29430.n12 0 0.018725f
C113 a_22190_29430.n14 0 0.062631f
C114 a_22190_29430.n16 0 0.030586f
C115 a_22190_29430.n17 0 0.059176f
C116 a_22190_29430.n19 0 0.059176f
C117 a_22190_29430.n21 0 0.059176f
C118 a_22190_29430.n22 0 0.018725f
C119 a_22190_29430.n23 0 0.030586f
C120 a_22190_29430.n24 0 0.059176f
C121 a_14558_34050.t25 0 0.049701f
C122 a_14558_34050.t12 0 0.049641f
C123 a_14558_34050.n0 0 0.259633f
C124 a_14558_34050.t19 0 0.049641f
C125 a_14558_34050.n1 0 0.136128f
C126 a_14558_34050.t28 0 0.049641f
C127 a_14558_34050.n2 0 0.136128f
C128 a_14558_34050.t15 0 0.049641f
C129 a_14558_34050.n3 0 0.136128f
C130 a_14558_34050.t13 0 0.049641f
C131 a_14558_34050.n4 0 0.136128f
C132 a_14558_34050.t22 0 0.049641f
C133 a_14558_34050.n5 0 0.136128f
C134 a_14558_34050.t10 0 0.049641f
C135 a_14558_34050.n6 0 0.136128f
C136 a_14558_34050.t17 0 0.049641f
C137 a_14558_34050.n7 0 0.136128f
C138 a_14558_34050.t21 0 0.049641f
C139 a_14558_34050.n8 0 0.337114f
C140 a_14558_34050.t20 0 0.049641f
C141 a_14558_34050.n9 0 0.337114f
C142 a_14558_34050.t29 0 0.049641f
C143 a_14558_34050.n10 0 0.136128f
C144 a_14558_34050.t16 0 0.049641f
C145 a_14558_34050.n11 0 0.136128f
C146 a_14558_34050.t24 0 0.049641f
C147 a_14558_34050.n12 0 0.136128f
C148 a_14558_34050.t11 0 0.049641f
C149 a_14558_34050.n13 0 0.136128f
C150 a_14558_34050.t18 0 0.049641f
C151 a_14558_34050.n14 0 0.136128f
C152 a_14558_34050.t27 0 0.049641f
C153 a_14558_34050.n15 0 0.136128f
C154 a_14558_34050.t14 0 0.049641f
C155 a_14558_34050.n16 0 0.136128f
C156 a_14558_34050.t23 0 0.049641f
C157 a_14558_34050.n17 0 0.136128f
C158 a_14558_34050.t26 0 0.049641f
C159 a_14558_34050.n18 0 0.992373f
C160 a_14558_34050.t1 0 0.434311f
C161 a_14558_34050.t4 0 0.028712f
C162 a_14558_34050.t2 0 0.028712f
C163 a_14558_34050.n19 0 0.062021f
C164 a_14558_34050.n20 0 1.41734f
C165 a_14558_34050.t8 0 0.028712f
C166 a_14558_34050.t9 0 0.028712f
C167 a_14558_34050.n21 0 0.062021f
C168 a_14558_34050.n22 0 0.627074f
C169 a_14558_34050.t6 0 0.028712f
C170 a_14558_34050.t7 0 0.028712f
C171 a_14558_34050.n23 0 0.062021f
C172 a_14558_34050.n24 0 0.614154f
C173 a_14558_34050.t3 0 0.028712f
C174 a_14558_34050.t5 0 0.028712f
C175 a_14558_34050.n25 0 0.062021f
C176 a_14558_34050.n26 0 0.715576f
C177 a_14558_34050.n27 0 4.21165f
C178 a_14558_34050.t0 0 0.341077f
C179 V_CONT.n5 0 0.058699f
C180 V_CONT.n9 0 0.017948f
C181 V_CONT.n10 0 0.014992f
C182 V_CONT.n11 0 0.082943f
C183 V_CONT.n12 0 0.02022f
C184 V_CONT.t5 0 6.66862f
C185 V_CONT.n13 0 0.162298f
C186 V_CONT.t7 0 0.019038f
C187 a_23100_30050.t1 0 0.027951f
C188 a_23100_30050.t0 0 0.027951f
C189 a_23100_30050.n0 0 0.149246f
C190 a_23100_30050.t3 0 0.030633f
C191 a_23100_30050.t8 0 0.069862f
C192 a_23100_30050.n1 0 0.179221f
C193 a_23100_30050.t7 0 0.034065f
C194 a_23100_30050.t6 0 0.070751f
C195 a_23100_30050.n2 0 0.099239f
C196 a_23100_30050.t5 0 0.069179f
C197 a_23100_30050.t4 0 0.104293f
C198 a_23100_30050.n3 0 1.26639f
C199 a_23100_30050.n4 0 0.267564f
C200 a_23100_30050.n5 0 0.256539f
C201 a_23100_30050.t2 0 0.147114f
C202 a_14990_33500.t4 0 0.051177f
C203 a_14990_33500.t3 0 0.051177f
C204 a_14990_33500.n0 0 0.127305f
C205 a_14990_33500.t2 0 0.051177f
C206 a_14990_33500.t1 0 0.051177f
C207 a_14990_33500.n1 0 0.122339f
C208 a_14990_33500.n2 0 1.74488f
C209 a_14990_33500.t6 0 0.026228f
C210 a_14990_33500.t10 0 0.026177f
C211 a_14990_33500.n3 0 0.184117f
C212 a_14990_33500.t8 0 0.026177f
C213 a_14990_33500.n4 0 0.114474f
C214 a_14990_33500.t9 0 0.026177f
C215 a_14990_33500.n5 0 0.114474f
C216 a_14990_33500.t7 0 0.026177f
C217 a_14990_33500.n6 0 0.383297f
C218 a_14990_33500.n7 0 0.903315f
C219 a_14990_33500.t5 0 0.191955f
C220 a_14990_33500.n8 0 2.2109f
C221 a_14990_33500.t0 0 0.267299f
C222 a_17540_31010.t4 0 0.04324f
C223 a_17540_31010.t0 0 1.74484f
C224 a_17540_31010.t1 0 0.045667f
C225 a_17540_31010.n0 0 1.57161f
C226 a_17540_31010.t7 0 0.016248f
C227 a_17540_31010.t6 0 0.016248f
C228 a_17540_31010.n1 0 0.053414f
C229 a_17540_31010.t3 0 0.04324f
C230 a_17540_31010.t2 0 0.04324f
C231 a_17540_31010.n2 0 0.106515f
C232 a_17540_31010.n3 0 1.2172f
C233 a_17540_31010.n4 0 2.04879f
C234 a_17540_31010.n5 0 0.106515f
C235 a_17540_31010.t5 0 0.04324f
C236 a_19190_29290.t9 0 0.018056f
C237 a_19190_29290.t1 0 0.018056f
C238 a_19190_29290.t7 0 0.018056f
C239 a_19190_29290.n0 0 0.036969f
C240 a_19190_29290.t0 0 0.021667f
C241 a_19190_29290.t20 0 0.021667f
C242 a_19190_29290.t21 0 0.034973f
C243 a_19190_29290.n1 0 0.039055f
C244 a_19190_29290.n2 0 0.02668f
C245 a_19190_29290.t6 0 0.027505f
C246 a_19190_29290.n3 0 0.043175f
C247 a_19190_29290.n4 0 0.191386f
C248 a_19190_29290.t3 0 0.018056f
C249 a_19190_29290.t5 0 0.018056f
C250 a_19190_29290.n5 0 0.036969f
C251 a_19190_29290.t2 0 0.021667f
C252 a_19190_29290.t22 0 0.021667f
C253 a_19190_29290.t17 0 0.034973f
C254 a_19190_29290.n6 0 0.039055f
C255 a_19190_29290.n7 0 0.02668f
C256 a_19190_29290.t4 0 0.027505f
C257 a_19190_29290.n8 0 0.043175f
C258 a_19190_29290.n9 0 0.191386f
C259 a_19190_29290.n10 0 0.26218f
C260 a_19190_29290.n11 0 0.019256f
C261 a_19190_29290.t13 0 0.034183f
C262 a_19190_29290.n12 0 0.021429f
C263 a_19190_29290.n13 0 0.554666f
C264 a_19190_29290.n14 0 0.186578f
C265 a_19190_29290.t8 0 0.021667f
C266 a_19190_29290.t19 0 0.021667f
C267 a_19190_29290.t18 0 0.034973f
C268 a_19190_29290.n15 0 0.039055f
C269 a_19190_29290.n16 0 0.02668f
C270 a_19190_29290.t10 0 0.027505f
C271 a_19190_29290.n17 0 0.043175f
C272 a_19190_29290.n18 0 0.239421f
C273 a_19190_29290.n19 0 0.036969f
C274 a_19190_29290.t11 0 0.018056f
C275 a_19940_23090.n3 0 0.026407f
C276 a_19940_23090.t13 0 1.95068f
C277 a_19940_23090.n4 0 0.016771f
C278 a_19940_23090.t8 0 0.021093f
C279 a_19940_23090.n5 0 0.036166f
C280 a_19940_23090.n6 0 0.010682f
C281 a_19940_23090.t10 0 0.011451f
C282 a_19940_23090.t11 0 0.011451f
C283 a_19940_23090.n7 0 0.013804f
C284 a_19940_23090.t14 0 0.026214f
C285 a_19940_23090.n8 0 0.013804f
C286 a_19940_23090.n9 0 0.013804f
C287 a_19940_23090.t15 0 0.019692f
C288 a_19940_23090.n10 0 0.012571f
C289 a_19940_23090.n11 0 0.186702f
C290 a_19940_23090.n12 0 0.09631f
C291 a_19940_23090.t12 0 1.95141f
C292 a_19940_23090.n13 0 0.016583f
C293 a_19940_23090.n14 0 0.01966f
C294 a_13532_27710.t10 0 0.31433f
C295 a_13532_27710.t17 0 0.331199f
C296 a_13532_27710.t11 0 0.331199f
C297 a_13532_27710.t19 0 0.331199f
C298 a_13532_27710.t3 0 0.331199f
C299 a_13532_27710.t6 0 0.331199f
C300 a_13532_27710.t4 0 0.331199f
C301 a_13532_27710.t8 0 0.331199f
C302 a_13532_27710.t14 0 0.315469f
C303 a_13532_27710.t9 0 0.151964f
C304 a_13532_27710.n0 0 0.19601f
C305 a_13532_27710.t15 0 0.344559f
C306 a_13532_27710.t20 0 0.316794f
C307 a_13532_27710.t13 0 0.331199f
C308 a_13532_27710.t7 0 0.331199f
C309 a_13532_27710.t12 0 0.331199f
C310 a_13532_27710.t5 0 0.331199f
C311 a_13532_27710.t2 0 0.331199f
C312 a_13532_27710.t18 0 0.331199f
C313 a_13532_27710.t1 0 0.331199f
C314 a_13532_27710.t16 0 0.743991f
C315 a_13532_27710.t0 0 0.080098f
C316 a_20480_25210.t6 0 0.078785f
C317 a_20480_25210.t4 0 0.030346f
C318 a_20480_25210.n0 0 0.120193f
C319 a_20480_25210.t11 0 0.020046f
C320 a_20480_25210.t5 0 0.020046f
C321 a_20480_25210.n1 0 0.046f
C322 a_20480_25210.n2 0 0.087576f
C323 a_20480_25210.t3 0 0.050114f
C324 a_20480_25210.t1 0 0.050114f
C325 a_20480_25210.n3 0 0.291421f
C326 a_20480_25210.t2 0 0.050114f
C327 a_20480_25210.t0 0 0.050114f
C328 a_20480_25210.n4 0 0.1426f
C329 a_20480_25210.n5 0 0.355827f
C330 a_20480_25210.n6 0 0.128581f
C331 a_20480_25210.t10 0 0.020046f
C332 a_20480_25210.t12 0 0.020046f
C333 a_20480_25210.n7 0 0.045548f
C334 a_20480_25210.n8 0 0.08916f
C335 a_20480_25210.t9 0 0.020046f
C336 a_20480_25210.t13 0 0.020046f
C337 a_20480_25210.n9 0 0.045548f
C338 a_20480_25210.n10 0 0.088358f
C339 a_20480_25210.t7 0 0.030346f
C340 a_20480_25210.n11 0 0.120193f
C341 a_20480_25210.t8 0 0.078785f
C342 a_14730_30630.n0 0 0.226228f
C343 a_14730_30630.n1 0 0.12827f
C344 a_14730_30630.n2 0 0.203125f
C345 a_14730_30630.n3 0 0.200529f
C346 a_14730_30630.t7 0 0.044358f
C347 a_14730_30630.t6 0 0.044358f
C348 a_14730_30630.n4 0 0.118669f
C349 a_14730_30630.t4 0 0.044358f
C350 a_14730_30630.t5 0 0.044358f
C351 a_14730_30630.n5 0 0.107634f
C352 a_14730_30630.n6 0 1.21683f
C353 a_14730_30630.t0 0 0.014786f
C354 a_14730_30630.t3 0 0.014786f
C355 a_14730_30630.n7 0 0.041682f
C356 a_14730_30630.n8 0 0.860437f
C357 a_14730_30630.t8 0 0.024477f
C358 a_14730_30630.t12 0 0.023979f
C359 a_14730_30630.n9 0 0.186829f
C360 a_14730_30630.t10 0 0.023979f
C361 a_14730_30630.n10 0 0.099745f
C362 a_14730_30630.t11 0 0.024302f
C363 a_14730_30630.n11 0 0.100457f
C364 a_14730_30630.t9 0 0.024302f
C365 a_14730_30630.n12 0 0.34311f
C366 a_14730_30630.n13 0 0.545948f
C367 a_14730_30630.t2 0 0.146843f
C368 a_14730_30630.n14 0 1.00301f
C369 a_14730_30630.n15 0 2.40266f
C370 a_14730_30630.n16 0 0.481345f
C371 a_14730_30630.t1 0 0.538618f
C372 a_14730_30630.n17 0 0.224971f
C373 a_14730_30630.n18 0 0.12827f
C374 a_14730_30630.n19 0 0.115443f
C375 a_14730_30630.n20 0 0.624567f
C376 a_14730_30630.n21 0 0.334582f
C377 a_14730_30630.n22 0 0.202918f
C378 a_14730_30630.n23 0 0.089235f
C379 a_25860_20180.t2 0 0.104706f
C380 a_25860_20180.n0 0 0.184398f
C381 a_25860_20180.t4 0 0.298444f
C382 a_25860_20180.t5 0 0.298444f
C383 a_25860_20180.t3 0 0.497217f
C384 a_25860_20180.n1 0 0.243367f
C385 a_25860_20180.n2 0 0.217957f
C386 a_25860_20180.t1 0 0.298444f
C387 a_25860_20180.n3 0 0.169192f
C388 a_25860_20180.n4 0 0.045341f
C389 a_25860_20180.n5 0 0.177419f
C390 a_25860_20180.t0 0 0.165068f
C391 a_18974_25970.t3 0 0.042383f
C392 a_18974_25970.t8 0 0.314286f
C393 a_18974_25970.t2 0 0.116977f
C394 a_18974_25970.t12 0 0.116977f
C395 a_18974_25970.t10 0 0.160839f
C396 a_18974_25970.n0 0 0.090068f
C397 a_18974_25970.n1 0 0.063914f
C398 a_18974_25970.n2 0 0.027464f
C399 a_18974_25970.t0 0 0.116977f
C400 a_18974_25970.t6 0 0.116977f
C401 a_18974_25970.n3 0 0.063914f
C402 a_18974_25970.n4 0 0.063914f
C403 a_18974_25970.t4 0 0.116977f
C404 a_18974_25970.t9 0 0.116977f
C405 a_18974_25970.t11 0 0.160839f
C406 a_18974_25970.n5 0 0.090068f
C407 a_18974_25970.n6 0 0.063914f
C408 a_18974_25970.n7 0 0.027591f
C409 a_18974_25970.t1 0 0.042383f
C410 a_18974_25970.t5 0 0.042383f
C411 a_18974_25970.n8 0 0.119624f
C412 a_18974_25970.n9 0 0.145636f
C413 a_18974_25970.n10 0 0.520173f
C414 a_18974_25970.n11 0 0.116362f
C415 a_18974_25970.t7 0 0.042383f
C416 a_19190_31850.n0 0 0.454298f
C417 a_19190_31850.n1 0 0.360667f
C418 a_19190_31850.n2 0 0.360667f
C419 a_19190_31850.n3 0 0.541f
C420 a_19190_31850.n4 0 0.360667f
C421 a_19190_31850.n5 0 0.360667f
C422 a_19190_31850.n6 0 0.360667f
C423 a_19190_31850.n7 0 0.360667f
C424 a_19190_31850.n8 0 1.23776f
C425 a_19190_31850.t9 0 0.010305f
C426 a_19190_31850.t25 0 0.0244f
C427 a_19190_31850.t31 0 0.41219f
C428 a_19190_31850.t23 0 0.419031f
C429 a_19190_31850.t16 0 0.41219f
C430 a_19190_31850.t21 0 0.41219f
C431 a_19190_31850.t15 0 0.41219f
C432 a_19190_31850.t36 0 0.41219f
C433 a_19190_31850.t28 0 0.41219f
C434 a_19190_31850.t34 0 0.41219f
C435 a_19190_31850.t27 0 0.41219f
C436 a_19190_31850.t18 0 0.41219f
C437 a_19190_31850.t24 0 0.41219f
C438 a_19190_31850.t26 0 0.41219f
C439 a_19190_31850.t33 0 0.41219f
C440 a_19190_31850.t13 0 0.41219f
C441 a_19190_31850.t35 0 0.41219f
C442 a_19190_31850.t14 0 0.41219f
C443 a_19190_31850.t20 0 0.41219f
C444 a_19190_31850.t29 0 0.41219f
C445 a_19190_31850.t22 0 0.41219f
C446 a_19190_31850.t30 0 0.41219f
C447 a_19190_31850.n9 0 0.949842f
C448 a_19190_31850.t5 0 0.010305f
C449 a_19190_31850.t6 0 0.010305f
C450 a_19190_31850.n10 0 0.022597f
C451 a_19190_31850.n11 0 0.215358f
C452 a_19190_31850.t19 0 0.015954f
C453 a_19190_31850.t17 0 0.015954f
C454 a_19190_31850.n12 0 0.029642f
C455 a_19190_31850.t1 0 0.018148f
C456 a_19190_31850.n13 0 0.013021f
C457 a_19190_31850.n14 0 0.012563f
C458 a_19190_31850.n15 0 0.335083f
C459 a_19190_31850.n16 0 0.110146f
C460 a_19190_31850.n17 0 0.06623f
C461 a_19190_31850.n18 0 0.074194f
C462 a_19190_31850.t8 0 0.010305f
C463 a_19190_31850.t7 0 0.010305f
C464 a_19190_31850.n19 0 0.022597f
C465 a_19190_31850.n20 0 0.169072f
C466 a_19190_31850.t12 0 0.015954f
C467 a_19190_31850.t11 0 0.015954f
C468 a_19190_31850.n21 0 0.030906f
C469 a_19190_31850.n22 0 0.119581f
C470 a_19190_31850.t32 0 0.024727f
C471 a_19190_31850.n23 0 0.245331f
C472 a_19190_31850.n24 0 0.022597f
C473 a_19190_31850.t10 0 0.010305f
C474 a_19190_31610.t12 0 0.016667f
C475 a_19190_31610.t8 0 0.016667f
C476 a_19190_31610.t10 0 0.016667f
C477 a_19190_31610.n0 0 0.034125f
C478 a_19190_31610.t7 0 0.025389f
C479 a_19190_31610.t9 0 0.02f
C480 a_19190_31610.t22 0 0.02f
C481 a_19190_31610.t21 0 0.032283f
C482 a_19190_31610.n1 0 0.036051f
C483 a_19190_31610.n2 0 0.024627f
C484 a_19190_31610.n3 0 0.039854f
C485 a_19190_31610.n4 0 0.176664f
C486 a_19190_31610.t4 0 0.016667f
C487 a_19190_31610.t6 0 0.016667f
C488 a_19190_31610.n5 0 0.034125f
C489 a_19190_31610.t3 0 0.025389f
C490 a_19190_31610.t5 0 0.02f
C491 a_19190_31610.t18 0 0.02f
C492 a_19190_31610.t17 0 0.032283f
C493 a_19190_31610.n6 0 0.036051f
C494 a_19190_31610.n7 0 0.024627f
C495 a_19190_31610.n8 0 0.039854f
C496 a_19190_31610.n9 0 0.176664f
C497 a_19190_31610.n10 0 0.242013f
C498 a_19190_31610.n11 0 0.017774f
C499 a_19190_31610.t16 0 0.031554f
C500 a_19190_31610.n12 0 0.019781f
C501 a_19190_31610.n13 0 0.511999f
C502 a_19190_31610.n14 0 0.172226f
C503 a_19190_31610.t11 0 0.025389f
C504 a_19190_31610.t13 0 0.02f
C505 a_19190_31610.t19 0 0.02f
C506 a_19190_31610.t20 0 0.032283f
C507 a_19190_31610.n15 0 0.036051f
C508 a_19190_31610.n16 0 0.024627f
C509 a_19190_31610.n17 0 0.039854f
C510 a_19190_31610.n18 0 0.221004f
C511 a_19190_31610.n19 0 0.034125f
C512 a_19190_31610.t14 0 0.016667f
C513 a_14348_27710.t37 0 0.176337f
C514 a_14348_27710.n0 0 0.064494f
C515 a_14348_27710.t38 0 0.1754f
C516 a_14348_27710.n1 0 0.073075f
C517 a_14348_27710.t27 0 0.177279f
C518 a_14348_27710.t28 0 0.176515f
C519 a_14348_27710.n2 0 0.219612f
C520 a_14348_27710.t15 0 0.176515f
C521 a_14348_27710.n3 0 0.121656f
C522 a_14348_27710.t16 0 0.176515f
C523 a_14348_27710.n4 0 0.121656f
C524 a_14348_27710.t18 0 0.176515f
C525 a_14348_27710.n5 0 0.121656f
C526 a_14348_27710.t19 0 0.176515f
C527 a_14348_27710.n6 0 0.121656f
C528 a_14348_27710.t20 0 0.176515f
C529 a_14348_27710.n7 0 0.121656f
C530 a_14348_27710.t42 0 0.177201f
C531 a_14348_27710.n8 0 0.113324f
C532 a_14348_27710.n9 0 0.034404f
C533 a_14348_27710.t48 0 0.177779f
C534 a_14348_27710.t47 0 0.176515f
C535 a_14348_27710.n10 0 0.220068f
C536 a_14348_27710.t46 0 0.176515f
C537 a_14348_27710.n11 0 0.121656f
C538 a_14348_27710.t33 0 0.176515f
C539 a_14348_27710.n12 0 0.121656f
C540 a_14348_27710.t40 0 0.176515f
C541 a_14348_27710.n13 0 0.121656f
C542 a_14348_27710.t39 0 0.176515f
C543 a_14348_27710.n14 0 0.121656f
C544 a_14348_27710.n15 0 0.034404f
C545 a_14348_27710.n16 0 0.022936f
C546 a_14348_27710.n17 0 0.127424f
C547 a_14348_27710.t9 0 0.174413f
C548 a_14348_27710.n18 0 0.48222f
C549 a_14348_27710.t13 0 0.012742f
C550 a_14348_27710.t3 0 0.012742f
C551 a_14348_27710.n19 0 0.027525f
C552 a_14348_27710.n20 0 0.259414f
C553 a_14348_27710.t6 0 0.012742f
C554 a_14348_27710.t7 0 0.012742f
C555 a_14348_27710.n21 0 0.027525f
C556 a_14348_27710.n22 0 0.278292f
C557 a_14348_27710.t8 0 0.012742f
C558 a_14348_27710.t4 0 0.012742f
C559 a_14348_27710.n23 0 0.027525f
C560 a_14348_27710.n24 0 0.270646f
C561 a_14348_27710.t2 0 0.012742f
C562 a_14348_27710.t10 0 0.012742f
C563 a_14348_27710.n25 0 0.02609f
C564 a_14348_27710.t12 0 0.012742f
C565 a_14348_27710.t1 0 0.012742f
C566 a_14348_27710.n26 0 0.029654f
C567 a_14348_27710.n27 0 0.349463f
C568 a_14348_27710.t5 0 0.012742f
C569 a_14348_27710.t11 0 0.012742f
C570 a_14348_27710.n28 0 0.02609f
C571 a_14348_27710.n29 0 0.216014f
C572 a_14348_27710.n30 0 0.654381f
C573 a_14348_27710.t14 0 0.509694f
C574 a_14348_27710.t23 0 0.518153f
C575 a_14348_27710.t43 0 0.509694f
C576 a_14348_27710.n31 0 0.338771f
C577 a_14348_27710.t22 0 0.509694f
C578 a_14348_27710.n32 0 0.222991f
C579 a_14348_27710.t41 0 0.509694f
C580 a_14348_27710.n33 0 0.222991f
C581 a_14348_27710.t32 0 0.509694f
C582 a_14348_27710.n34 0 0.222991f
C583 a_14348_27710.t26 0 0.509694f
C584 a_14348_27710.n35 0 0.222991f
C585 a_14348_27710.t31 0 0.509694f
C586 a_14348_27710.n36 0 0.222991f
C587 a_14348_27710.t25 0 0.509694f
C588 a_14348_27710.n37 0 0.222991f
C589 a_14348_27710.t44 0 0.509694f
C590 a_14348_27710.n38 0 0.215027f
C591 a_14348_27710.t24 0 0.509694f
C592 a_14348_27710.n39 0 0.230955f
C593 a_14348_27710.n40 0 0.230955f
C594 a_14348_27710.t36 0 0.509694f
C595 a_14348_27710.n41 0 0.215027f
C596 a_14348_27710.t17 0 0.509694f
C597 a_14348_27710.n42 0 0.222991f
C598 a_14348_27710.t29 0 0.509694f
C599 a_14348_27710.n43 0 0.222991f
C600 a_14348_27710.t21 0 0.509694f
C601 a_14348_27710.n44 0 0.222991f
C602 a_14348_27710.t30 0 0.509694f
C603 a_14348_27710.n45 0 0.222991f
C604 a_14348_27710.t34 0 0.509694f
C605 a_14348_27710.n46 0 0.222991f
C606 a_14348_27710.t45 0 0.509694f
C607 a_14348_27710.n47 0 0.222991f
C608 a_14348_27710.t35 0 0.509694f
C609 a_14348_27710.n48 0 0.221398f
C610 a_14348_27710.t49 0 0.509694f
C611 a_14348_27710.n49 0 0.391094f
C612 a_14348_27710.n50 0 1.23441f
C613 a_14348_27710.t0 0 0.111663f
C614 a_19190_29050.n0 0 1.02458f
C615 a_19190_29050.n1 0 1.10014f
C616 a_19190_29050.n2 0 1.33269f
C617 a_19190_29050.n3 0 0.153679f
C618 a_19190_29050.n4 0 3.88852f
C619 a_19190_29050.t36 0 0.021247f
C620 a_19190_29050.n5 0 0.019024f
C621 a_19190_29050.t17 0 0.013904f
C622 a_19190_29050.t13 0 0.013904f
C623 a_19190_29050.n6 0 0.026482f
C624 a_19190_29050.t25 0 0.359229f
C625 a_19190_29050.t18 0 0.36519f
C626 a_19190_29050.t35 0 0.359229f
C627 a_19190_29050.t15 0 0.359229f
C628 a_19190_29050.t33 0 0.359229f
C629 a_19190_29050.t29 0 0.359229f
C630 a_19190_29050.t22 0 0.359229f
C631 a_19190_29050.t27 0 0.359229f
C632 a_19190_29050.t21 0 0.359229f
C633 a_19190_29050.t12 0 0.359229f
C634 a_19190_29050.t19 0 0.359229f
C635 a_19190_29050.t20 0 0.359229f
C636 a_19190_29050.t26 0 0.359229f
C637 a_19190_29050.t31 0 0.359229f
C638 a_19190_29050.t28 0 0.359229f
C639 a_19190_29050.t32 0 0.359229f
C640 a_19190_29050.t14 0 0.359229f
C641 a_19190_29050.t23 0 0.359229f
C642 a_19190_29050.t16 0 0.359229f
C643 a_19190_29050.t24 0 0.359229f
C644 a_19190_29050.t30 0 0.021589f
C645 a_19190_29050.n7 0 0.019024f
C646 a_19190_29050.t6 0 0.015816f
C647 a_19190_29050.n8 0 0.011348f
C648 a_19190_29050.n9 0 0.010949f
C649 a_19190_29050.n10 0 0.292028f
C650 a_19190_29050.t11 0 0.013904f
C651 a_19190_29050.t34 0 0.013904f
C652 a_19190_29050.n11 0 0.025867f
C653 a_19190_29050.n12 0 0.019024f
C654 VDPWR.n7 0 0.011667f
C655 VDPWR.n11 0 0.011667f
C656 VDPWR.t258 0 0.078178f
C657 VDPWR.n21 0 0.010035f
C658 VDPWR.n22 0 0.034562f
C659 VDPWR.t84 0 0.0357f
C660 VDPWR.t51 0 0.060554f
C661 VDPWR.t82 0 0.060554f
C662 VDPWR.t193 0 0.039767f
C663 VDPWR.t12 0 0.039767f
C664 VDPWR.t211 0 0.019883f
C665 VDPWR.t262 0 0.065977f
C666 VDPWR.t93 0 0.068236f
C667 VDPWR.t102 0 0.028469f
C668 VDPWR.n47 0 0.011667f
C669 VDPWR.n54 0 0.013388f
C670 VDPWR.n56 0 0.0123f
C671 VDPWR.n62 0 0.0123f
C672 VDPWR.n70 0 0.011667f
C673 VDPWR.n77 0 0.011667f
C674 VDPWR.n97 0 0.011667f
C675 VDPWR.n100 0 0.013388f
C676 VDPWR.t260 0 0.032536f
C677 VDPWR.t34 0 0.032536f
C678 VDPWR.t17 0 0.054227f
C679 VDPWR.t390 0 0.056487f
C680 VDPWR.n105 0 0.010035f
C681 VDPWR.n106 0 0.027332f
C682 VDPWR.t114 0 0.028469f
C683 VDPWR.t56 0 0.032536f
C684 VDPWR.t209 0 0.032536f
C685 VDPWR.t89 0 0.054227f
C686 VDPWR.t110 0 0.056487f
C687 VDPWR.t201 0 0.028469f
C688 VDPWR.n117 0 0.011667f
C689 VDPWR.n125 0 0.013388f
C690 VDPWR.n140 0 0.12177f
C691 VDPWR.t404 0 0.407866f
C692 VDPWR.n142 0 0.271911f
C693 VDPWR.t60 0 0.012176f
C694 VDPWR.n144 0 0.010011f
C695 VDPWR.n146 0 0.010011f
C696 VDPWR.n148 0 0.029299f
C697 VDPWR.t405 0 0.018164f
C698 VDPWR.n150 0 0.018936f
C699 VDPWR.n151 0 0.018936f
C700 VDPWR.n154 0 0.033832f
C701 VDPWR.n155 0 0.091555f
C702 VDPWR.t98 0 0.210819f
C703 VDPWR.t59 0 0.166168f
C704 VDPWR.n156 0 0.234146f
C705 VDPWR.t67 0 0.012176f
C706 VDPWR.t61 0 0.032536f
C707 VDPWR.t417 0 0.032536f
C708 VDPWR.t374 0 0.050323f
C709 VDPWR.t68 0 0.236759f
C710 VDPWR.t122 0 0.210819f
C711 VDPWR.t69 0 0.012176f
C712 VDPWR.n160 0 0.089828f
C713 VDPWR.t123 0 0.018155f
C714 VDPWR.n162 0 0.016279f
C715 VDPWR.n164 0 0.01205f
C716 VDPWR.n165 0 0.01205f
C717 VDPWR.n167 0 0.02319f
C718 VDPWR.n169 0 0.234146f
C719 VDPWR.t66 0 0.166168f
C720 VDPWR.t100 0 0.210819f
C721 VDPWR.n170 0 0.089828f
C722 VDPWR.n172 0 0.02319f
C723 VDPWR.t101 0 0.018155f
C724 VDPWR.n174 0 0.01205f
C725 VDPWR.n175 0 0.01205f
C726 VDPWR.n178 0 0.016279f
C727 VDPWR.n188 0 0.124902f
C728 VDPWR.n189 0 0.09212f
C729 VDPWR.n191 0 0.014578f
C730 VDPWR.n197 0 0.011667f
C731 VDPWR.n204 0 0.010035f
C732 VDPWR.n205 0 0.027332f
C733 VDPWR.t73 0 0.056487f
C734 VDPWR.t70 0 0.054227f
C735 VDPWR.t87 0 0.032536f
C736 VDPWR.t95 0 0.032536f
C737 VDPWR.t77 0 0.028469f
C738 VDPWR.n206 0 0.027332f
C739 VDPWR.n207 0 0.010035f
C740 VDPWR.n237 0 0.013388f
C741 VDPWR.n243 0 0.011667f
C742 VDPWR.n250 0 0.010035f
C743 VDPWR.n251 0 0.027332f
C744 VDPWR.t21 0 0.058294f
C745 VDPWR.t384 0 0.056035f
C746 VDPWR.t256 0 0.039767f
C747 VDPWR.t394 0 0.039767f
C748 VDPWR.t153 0 0.05242f
C749 VDPWR.t351 0 0.05242f
C750 VDPWR.t125 0 0.032536f
C751 VDPWR.t162 0 0.032536f
C752 VDPWR.t10 0 0.04067f
C753 VDPWR.t423 0 0.04067f
C754 VDPWR.t75 0 0.0357f
C755 VDPWR.n252 0 0.034562f
C756 VDPWR.n253 0 0.010035f
C757 VDPWR.n265 0 0.014011f
C758 VDPWR.n291 0 0.082532f
C759 VDPWR.n292 0 0.011462f
C760 VDPWR.n298 0 0.010329f
C761 VDPWR.n300 0 0.010011f
C762 VDPWR.n305 0 0.01205f
C763 VDPWR.n307 0 0.01205f
C764 VDPWR.n308 0 0.016766f
C765 VDPWR.t416 0 0.018155f
C766 VDPWR.n310 0 0.017375f
C767 VDPWR.n314 0 0.01205f
C768 VDPWR.n315 0 0.017375f
C769 VDPWR.n317 0 0.01205f
C770 VDPWR.t119 0 0.018155f
C771 VDPWR.n319 0 0.016766f
C772 VDPWR.n321 0 0.157431f
C773 VDPWR.t118 0 0.130748f
C774 VDPWR.t174 0 0.277506f
C775 VDPWR.t124 0 0.277506f
C776 VDPWR.t178 0 0.130748f
C777 VDPWR.n325 0 0.010011f
C778 VDPWR.n326 0 0.022664f
C779 VDPWR.t350 0 0.018164f
C780 VDPWR.n329 0 0.018936f
C781 VDPWR.n330 0 0.018936f
C782 VDPWR.n331 0 0.010011f
C783 VDPWR.n332 0 0.018877f
C784 VDPWR.t246 0 0.018164f
C785 VDPWR.n336 0 0.018936f
C786 VDPWR.n337 0 0.018936f
C787 VDPWR.n338 0 0.010011f
C788 VDPWR.n339 0 0.022664f
C789 VDPWR.n369 0 0.015494f
C790 VDPWR.n380 0 0.01205f
C791 VDPWR.n383 0 0.01205f
C792 VDPWR.n384 0 0.016766f
C793 VDPWR.t141 0 0.018155f
C794 VDPWR.n386 0 0.017017f
C795 VDPWR.n387 0 0.01205f
C796 VDPWR.n390 0 0.01205f
C797 VDPWR.n391 0 0.016766f
C798 VDPWR.t208 0 0.018155f
C799 VDPWR.n393 0 0.017017f
C800 VDPWR.n396 0 0.01205f
C801 VDPWR.n399 0 0.01205f
C802 VDPWR.n400 0 0.016766f
C803 VDPWR.t128 0 0.018155f
C804 VDPWR.n402 0 0.017017f
C805 VDPWR.n403 0 0.01205f
C806 VDPWR.n406 0 0.01205f
C807 VDPWR.n407 0 0.016766f
C808 VDPWR.t393 0 0.018155f
C809 VDPWR.n409 0 0.017017f
C810 VDPWR.t397 0 0.02667f
C811 VDPWR.n410 0 0.028763f
C812 VDPWR.n428 0 0.01205f
C813 VDPWR.n431 0 0.01205f
C814 VDPWR.n432 0 0.016766f
C815 VDPWR.t224 0 0.018155f
C816 VDPWR.n434 0 0.017375f
C817 VDPWR.n435 0 0.01205f
C818 VDPWR.n438 0 0.01205f
C819 VDPWR.n439 0 0.016766f
C820 VDPWR.t425 0 0.018155f
C821 VDPWR.n441 0 0.017375f
C822 VDPWR.n447 0 0.01205f
C823 VDPWR.n450 0 0.01205f
C824 VDPWR.n451 0 0.016766f
C825 VDPWR.t369 0 0.018066f
C826 VDPWR.n453 0 0.017055f
C827 VDPWR.n455 0 0.01205f
C828 VDPWR.n458 0 0.01205f
C829 VDPWR.n459 0 0.016766f
C830 VDPWR.t235 0 0.018155f
C831 VDPWR.n461 0 0.017375f
C832 VDPWR.n483 0 0.015494f
C833 VDPWR.n486 0 0.015494f
C834 VDPWR.n487 0 0.020442f
C835 VDPWR.t367 0 0.024205f
C836 VDPWR.n489 0 0.020792f
C837 VDPWR.n490 0 0.015494f
C838 VDPWR.n493 0 0.015494f
C839 VDPWR.n494 0 0.020442f
C840 VDPWR.t148 0 0.024205f
C841 VDPWR.n496 0 0.020792f
C842 VDPWR.n503 0 0.015494f
C843 VDPWR.n506 0 0.015494f
C844 VDPWR.n507 0 0.020442f
C845 VDPWR.t144 0 0.024205f
C846 VDPWR.n509 0 0.020792f
C847 VDPWR.n513 0 0.066292f
C848 VDPWR.n517 0 0.015494f
C849 VDPWR.n520 0 0.015494f
C850 VDPWR.n521 0 0.020442f
C851 VDPWR.t33 0 0.024205f
C852 VDPWR.n523 0 0.020792f
C853 VDPWR.n524 0 0.015494f
C854 VDPWR.n527 0 0.015494f
C855 VDPWR.n528 0 0.020442f
C856 VDPWR.t155 0 0.024205f
C857 VDPWR.n530 0 0.020792f
C858 VDPWR.t428 0 0.386412f
C859 VDPWR.t430 0 0.40673f
C860 VDPWR.n541 0 0.748f
C861 VDPWR.t429 0 0.40673f
C862 VDPWR.n542 0 0.394833f
C863 VDPWR.t434 0 0.381702f
C864 VDPWR.n543 0 0.468568f
C865 VDPWR.t55 0 0.192464f
C866 VDPWR.t117 0 0.202793f
C867 VDPWR.t373 0 0.202793f
C868 VDPWR.t116 0 0.202793f
C869 VDPWR.t376 0 0.202793f
C870 VDPWR.t65 0 0.202793f
C871 VDPWR.t233 0 0.202793f
C872 VDPWR.t38 0 0.202793f
C873 VDPWR.t182 0 0.193161f
C874 VDPWR.t185 0 0.093047f
C875 VDPWR.n544 0 0.120017f
C876 VDPWR.t120 0 0.210973f
C877 VDPWR.t372 0 0.193973f
C878 VDPWR.t121 0 0.202793f
C879 VDPWR.t377 0 0.202793f
C880 VDPWR.t188 0 0.202793f
C881 VDPWR.t131 0 0.202793f
C882 VDPWR.t215 0 0.202793f
C883 VDPWR.t134 0 0.202793f
C884 VDPWR.t31 0 0.202793f
C885 VDPWR.t135 0 0.313233f
C886 VDPWR.n545 0 0.476642f
C887 VDPWR.n547 0 0.092042f
C888 VDPWR.n548 0 0.013387f
C889 VDPWR.t279 0 0.011976f
C890 VDPWR.n549 0 0.013285f
C891 VDPWR.n551 0 0.092042f
C892 VDPWR.n552 0 0.013387f
C893 VDPWR.t286 0 0.011976f
C894 VDPWR.n553 0 0.013387f
C895 VDPWR.t309 0 0.011976f
C896 VDPWR.n555 0 0.092042f
C897 VDPWR.n557 0 0.092042f
C898 VDPWR.n559 0 0.092042f
C899 VDPWR.n561 0 0.092042f
C900 VDPWR.n563 0 0.092042f
C901 VDPWR.n565 0 0.092042f
C902 VDPWR.n567 0 0.092042f
C903 VDPWR.n569 0 0.12542f
C904 VDPWR.n570 0 0.040251f
C905 VDPWR.n572 0 0.013285f
C906 VDPWR.n573 0 0.042441f
C907 VDPWR.t308 0 0.035731f
C908 VDPWR.t400 0 0.028921f
C909 VDPWR.t180 0 0.028921f
C910 VDPWR.t156 0 0.028921f
C911 VDPWR.t357 0 0.028921f
C912 VDPWR.t355 0 0.028921f
C913 VDPWR.t363 0 0.028921f
C914 VDPWR.t43 0 0.028921f
C915 VDPWR.t229 0 0.028921f
C916 VDPWR.t27 0 0.028921f
C917 VDPWR.t39 0 0.028921f
C918 VDPWR.t41 0 0.028921f
C919 VDPWR.t191 0 0.028921f
C920 VDPWR.t203 0 0.028921f
C921 VDPWR.t158 0 0.028921f
C922 VDPWR.t370 0 0.028921f
C923 VDPWR.t104 0 0.028921f
C924 VDPWR.t221 0 0.028921f
C925 VDPWR.t199 0 0.028921f
C926 VDPWR.t285 0 0.043946f
C927 VDPWR.n574 0 0.036636f
C928 VDPWR.n575 0 0.013285f
C929 VDPWR.n576 0 0.010227f
C930 VDPWR.n577 0 0.028426f
C931 VDPWR.n578 0 0.093567f
C932 VDPWR.n580 0 0.092042f
C933 VDPWR.n582 0 0.092042f
C934 VDPWR.n584 0 0.092042f
C935 VDPWR.n586 0 0.092042f
C936 VDPWR.n588 0 0.092042f
C937 VDPWR.n590 0 0.092042f
C938 VDPWR.n592 0 0.092042f
C939 VDPWR.n594 0 0.092042f
C940 VDPWR.n595 0 0.093567f
C941 VDPWR.n596 0 0.037905f
C942 VDPWR.t339 0 0.011976f
C943 VDPWR.n598 0 0.013387f
C944 VDPWR.n599 0 0.044557f
C945 VDPWR.t338 0 0.036024f
C946 VDPWR.t388 0 0.028921f
C947 VDPWR.t406 0 0.028921f
C948 VDPWR.t225 0 0.028921f
C949 VDPWR.t4 0 0.028921f
C950 VDPWR.t2 0 0.028921f
C951 VDPWR.t49 0 0.028921f
C952 VDPWR.t398 0 0.028921f
C953 VDPWR.t386 0 0.028921f
C954 VDPWR.t151 0 0.028921f
C955 VDPWR.t205 0 0.028921f
C956 VDPWR.t108 0 0.028921f
C957 VDPWR.t378 0 0.028921f
C958 VDPWR.t414 0 0.028921f
C959 VDPWR.t408 0 0.028921f
C960 VDPWR.t227 0 0.028921f
C961 VDPWR.t106 0 0.028921f
C962 VDPWR.t410 0 0.028921f
C963 VDPWR.t129 0 0.028921f
C964 VDPWR.t278 0 0.043276f
C965 VDPWR.n600 0 0.034895f
C966 VDPWR.n601 0 0.013285f
C967 VDPWR.n602 0 0.010227f
C968 VDPWR.n603 0 0.02133f
C969 VDPWR.n604 0 0.257688f
C970 VDPWR.n605 0 0.184855f
C971 VDPWR.n606 0 0.013475f
C972 VDPWR.t294 0 0.010759f
C973 VDPWR.t46 0 0.010759f
C974 VDPWR.n608 0 0.022533f
C975 VDPWR.t80 0 0.010759f
C976 VDPWR.t146 0 0.010759f
C977 VDPWR.n611 0 0.022533f
C978 VDPWR.t161 0 0.010759f
C979 VDPWR.t403 0 0.010759f
C980 VDPWR.n614 0 0.022533f
C981 VDPWR.t150 0 0.010759f
C982 VDPWR.t366 0 0.010759f
C983 VDPWR.n617 0 0.022533f
C984 VDPWR.n620 0 0.02379f
C985 VDPWR.t48 0 0.010759f
C986 VDPWR.t325 0 0.010759f
C987 VDPWR.n622 0 0.022533f
C988 VDPWR.n624 0 0.01897f
C989 VDPWR.n630 0 0.015494f
C990 VDPWR.n631 0 0.015401f
C991 VDPWR.n632 0 0.015494f
C992 VDPWR.n635 0 0.015494f
C993 VDPWR.t293 0 0.010759f
C994 VDPWR.n637 0 0.032278f
C995 VDPWR.t291 0 0.042636f
C996 VDPWR.n638 0 0.015043f
C997 VDPWR.n639 0 0.014744f
C998 VDPWR.n641 0 0.233973f
C999 VDPWR.t247 0 0.112758f
C1000 VDPWR.t292 0 0.073293f
C1001 VDPWR.t250 0 0.087388f
C1002 VDPWR.t81 0 0.098663f
C1003 VDPWR.t45 0 0.073293f
C1004 VDPWR.t251 0 0.112758f
C1005 VDPWR.t79 0 0.073293f
C1006 VDPWR.t177 0 0.08175f
C1007 VDPWR.t249 0 0.104301f
C1008 VDPWR.t145 0 0.143767f
C1009 VDPWR.t160 0 0.152224f
C1010 VDPWR.t297 0 0.015439f
C1011 VDPWR.n643 0 0.01897f
C1012 VDPWR.n644 0 0.011276f
C1013 VDPWR.n645 0 0.038401f
C1014 VDPWR.n646 0 0.121522f
C1015 VDPWR.t402 0 0.093026f
C1016 VDPWR.t296 0 0.093026f
C1017 VDPWR.t91 0 0.093026f
C1018 VDPWR.t149 0 0.073293f
C1019 VDPWR.t19 0 0.112758f
C1020 VDPWR.t365 0 0.073293f
C1021 VDPWR.t175 0 0.087388f
C1022 VDPWR.t136 0 0.098663f
C1023 VDPWR.t47 0 0.073293f
C1024 VDPWR.t317 0 0.112758f
C1025 VDPWR.t324 0 0.093026f
C1026 VDPWR.t319 0 0.015439f
C1027 VDPWR.n648 0 0.01897f
C1028 VDPWR.n649 0 0.011276f
C1029 VDPWR.n650 0 0.038401f
C1030 VDPWR.n651 0 0.109902f
C1031 VDPWR.n655 0 0.015494f
C1032 VDPWR.t326 0 0.010759f
C1033 VDPWR.n657 0 0.015494f
C1034 VDPWR.n660 0 0.015494f
C1035 VDPWR.t323 0 0.043509f
C1036 VDPWR.n661 0 0.030401f
C1037 VDPWR.n662 0 0.032278f
C1038 VDPWR.n663 0 0.013683f
C1039 VDPWR.n665 0 0.088915f
C1040 VDPWR.t305 0 0.015439f
C1041 VDPWR.n666 0 0.011276f
C1042 VDPWR.n667 0 0.038401f
C1043 VDPWR.n668 0 0.107427f
C1044 VDPWR.t304 0 0.166318f
C1045 VDPWR.t112 0 0.146586f
C1046 VDPWR.t239 0 0.146586f
C1047 VDPWR.t197 0 0.146586f
C1048 VDPWR.t8 0 0.146586f
C1049 VDPWR.t288 0 0.293278f
C1050 VDPWR.t290 0 0.015427f
C1051 VDPWR.n669 0 0.108517f
C1052 VDPWR.n670 0 0.011286f
C1053 VDPWR.n671 0 0.01897f
C1054 VDPWR.n672 0 0.025883f
C1055 VDPWR.n673 0 0.077897f
C1056 VDPWR.n674 0 0.077772f
C1057 VDPWR.n681 0 0.075421f
C1058 VDPWR.n688 0 0.075421f
C1059 VDPWR.n695 0 0.075421f
C1060 VDPWR.n702 0 0.075421f
C1061 VDPWR.n706 0 0.071875f
C1062 VDPWR.n707 0 0.119858f
C1063 VDPWR.t16 0 0.010329f
C1064 VDPWR.t54 0 0.010329f
C1065 VDPWR.n708 0 0.040189f
C1066 VDPWR.n709 0 0.138159f
C1067 VDPWR.t274 0 0.049253f
C1068 VDPWR.n713 0 0.01205f
C1069 VDPWR.n720 0 0.01205f
C1070 VDPWR.t133 0 0.010329f
C1071 VDPWR.t14 0 0.010329f
C1072 VDPWR.n721 0 0.040189f
C1073 VDPWR.n722 0 0.138159f
C1074 VDPWR.t422 0 0.010329f
C1075 VDPWR.t214 0 0.010329f
C1076 VDPWR.n723 0 0.040189f
C1077 VDPWR.n724 0 0.138159f
C1078 VDPWR.t184 0 0.010329f
C1079 VDPWR.t420 0 0.010329f
C1080 VDPWR.n725 0 0.040189f
C1081 VDPWR.n726 0 0.138159f
C1082 VDPWR.t64 0 0.010329f
C1083 VDPWR.t30 0 0.010329f
C1084 VDPWR.n727 0 0.040189f
C1085 VDPWR.n728 0 0.138159f
C1086 VDPWR.t381 0 0.010329f
C1087 VDPWR.t383 0 0.010329f
C1088 VDPWR.n729 0 0.040189f
C1089 VDPWR.n730 0 0.138159f
C1090 VDPWR.t187 0 0.010329f
C1091 VDPWR.t37 0 0.010329f
C1092 VDPWR.n731 0 0.040189f
C1093 VDPWR.n732 0 0.138159f
C1094 VDPWR.t190 0 0.010329f
C1095 VDPWR.t232 0 0.010329f
C1096 VDPWR.n733 0 0.040189f
C1097 VDPWR.n734 0 0.196839f
C1098 VDPWR.t313 0 0.049253f
C1099 VDPWR.n735 0 0.019892f
C1100 VDPWR.n736 0 0.0153f
C1101 VDPWR.n741 0 0.01205f
C1102 VDPWR.n743 0 0.011978f
C1103 VDPWR.n744 0 0.011978f
C1104 VDPWR.n746 0 0.01205f
C1105 VDPWR.n747 0 0.01205f
C1106 VDPWR.n749 0 0.014529f
C1107 VDPWR.n751 0 0.096576f
C1108 VDPWR.t314 0 0.102429f
C1109 VDPWR.t189 0 0.105356f
C1110 VDPWR.t231 0 0.105356f
C1111 VDPWR.t186 0 0.105356f
C1112 VDPWR.t36 0 0.105356f
C1113 VDPWR.t380 0 0.105356f
C1114 VDPWR.t382 0 0.105356f
C1115 VDPWR.t63 0 0.105356f
C1116 VDPWR.t29 0 0.105356f
C1117 VDPWR.t183 0 0.105356f
C1118 VDPWR.t419 0 0.105356f
C1119 VDPWR.t421 0 0.105356f
C1120 VDPWR.t213 0 0.105356f
C1121 VDPWR.t132 0 0.105356f
C1122 VDPWR.t13 0 0.105356f
C1123 VDPWR.t15 0 0.105356f
C1124 VDPWR.t53 0 0.105356f
C1125 VDPWR.t275 0 0.102429f
C1126 VDPWR.n755 0 0.011978f
C1127 VDPWR.n756 0 0.011978f
C1128 VDPWR.n757 0 0.01205f
C1129 VDPWR.n758 0 0.01205f
C1130 VDPWR.n760 0 0.014529f
C1131 VDPWR.n762 0 0.096576f
C1132 VDPWR.n766 0 0.01205f
C1133 VDPWR.n768 0 0.0153f
C1134 VDPWR.n769 0 0.018879f
C1135 VDPWR.n770 0 0.116502f
C1136 VDPWR.n771 0 0.114884f
C1137 VDPWR.n772 0 0.013387f
C1138 VDPWR.t273 0 0.011976f
C1139 VDPWR.n773 0 0.014077f
C1140 VDPWR.n774 0 0.043839f
C1141 VDPWR.t336 0 0.013662f
C1142 VDPWR.n776 0 0.014179f
C1143 VDPWR.n777 0 0.043106f
C1144 VDPWR.t335 0 0.035066f
C1145 VDPWR.t72 0 0.026511f
C1146 VDPWR.t236 0 0.026511f
C1147 VDPWR.t272 0 0.041613f
C1148 VDPWR.n778 0 0.034148f
C1149 VDPWR.n779 0 0.013285f
C1150 VDPWR.n780 0 0.010227f
C1151 VDPWR.n781 0 0.023591f
C1152 VDPWR.n782 0 0.28418f
C1153 VDPWR.n783 0 0.106679f
C1154 VDPWR.n785 0 0.040765f
C1155 VDPWR.n786 0 0.013489f
C1156 VDPWR.n787 0 0.013285f
C1157 VDPWR.t270 0 0.011976f
C1158 VDPWR.n790 0 0.040765f
C1159 VDPWR.n791 0 0.013489f
C1160 VDPWR.n792 0 0.013285f
C1161 VDPWR.t322 0 0.011976f
C1162 VDPWR.n795 0 0.040765f
C1163 VDPWR.n797 0 0.040765f
C1164 VDPWR.n799 0 0.040765f
C1165 VDPWR.n801 0 0.050361f
C1166 VDPWR.n802 0 0.017072f
C1167 VDPWR.n803 0 0.022672f
C1168 VDPWR.n804 0 0.013489f
C1169 VDPWR.n805 0 0.041771f
C1170 VDPWR.t321 0 0.03399f
C1171 VDPWR.t348 0 0.026511f
C1172 VDPWR.t166 0 0.026511f
C1173 VDPWR.t142 0 0.026511f
C1174 VDPWR.t168 0 0.026511f
C1175 VDPWR.t164 0 0.026511f
C1176 VDPWR.t219 0 0.026511f
C1177 VDPWR.t346 0 0.026511f
C1178 VDPWR.t266 0 0.026511f
C1179 VDPWR.t138 0 0.026511f
C1180 VDPWR.t170 0 0.026511f
C1181 VDPWR.t332 0 0.041613f
C1182 VDPWR.n806 0 0.034148f
C1183 VDPWR.t333 0 0.011976f
C1184 VDPWR.n807 0 0.013285f
C1185 VDPWR.n808 0 0.022672f
C1186 VDPWR.n809 0 0.016339f
C1187 VDPWR.n810 0 0.027544f
C1188 VDPWR.n812 0 0.040765f
C1189 VDPWR.n814 0 0.040765f
C1190 VDPWR.n816 0 0.040765f
C1191 VDPWR.n818 0 0.040765f
C1192 VDPWR.n819 0 0.027544f
C1193 VDPWR.n820 0 0.016339f
C1194 VDPWR.n821 0 0.022672f
C1195 VDPWR.n822 0 0.013489f
C1196 VDPWR.n823 0 0.041771f
C1197 VDPWR.t269 0 0.03399f
C1198 VDPWR.t217 0 0.026511f
C1199 VDPWR.t243 0 0.026511f
C1200 VDPWR.t344 0 0.026511f
C1201 VDPWR.t254 0 0.026511f
C1202 VDPWR.t264 0 0.026511f
C1203 VDPWR.t241 0 0.026511f
C1204 VDPWR.t252 0 0.026511f
C1205 VDPWR.t426 0 0.026511f
C1206 VDPWR.t353 0 0.026511f
C1207 VDPWR.t172 0 0.026511f
C1208 VDPWR.t311 0 0.041613f
C1209 VDPWR.n824 0 0.034148f
C1210 VDPWR.t312 0 0.011976f
C1211 VDPWR.n825 0 0.013285f
C1212 VDPWR.n826 0 0.022672f
C1213 VDPWR.n827 0 0.016339f
C1214 VDPWR.n828 0 0.130687f
C1215 VDPWR.n829 0 0.10531f
C1216 VDPWR.t299 0 0.042905f
C1217 VDPWR.n831 0 0.014883f
C1218 VDPWR.n833 0 0.024888f
C1219 VDPWR.n836 0 0.024888f
C1220 VDPWR.n838 0 0.024888f
C1221 VDPWR.n839 0 0.035021f
C1222 VDPWR.n842 0 0.033618f
C1223 VDPWR.n847 0 0.02214f
C1224 VDPWR.n852 0 0.015494f
C1225 VDPWR.n854 0 0.015494f
C1226 VDPWR.n855 0 0.020442f
C1227 VDPWR.t301 0 0.024205f
C1228 VDPWR.n857 0 0.019496f
C1229 VDPWR.n859 0 0.097351f
C1230 VDPWR.t300 0 0.107336f
C1231 VDPWR.t412 0 0.109832f
C1232 VDPWR.t361 0 0.109832f
C1233 VDPWR.t237 0 0.109832f
C1234 VDPWR.t0 0 0.109832f
C1235 VDPWR.t341 0 0.107336f
C1236 VDPWR.n862 0 0.024101f
C1237 VDPWR.t340 0 0.040485f
C1238 VDPWR.t280 0 0.040485f
C1239 VDPWR.n864 0 0.018239f
C1240 VDPWR.t282 0 0.024213f
C1241 VDPWR.n866 0 0.035417f
C1242 VDPWR.n867 0 0.012895f
C1243 VDPWR.n868 0 0.012895f
C1244 VDPWR.n869 0 0.024101f
C1245 VDPWR.n872 0 0.104839f
C1246 VDPWR.t281 0 0.107336f
C1247 VDPWR.t359 0 0.109832f
C1248 VDPWR.t6 0 0.109832f
C1249 VDPWR.t23 0 0.109832f
C1250 VDPWR.t195 0 0.109832f
C1251 VDPWR.t328 0 0.107336f
C1252 VDPWR.t330 0 0.024205f
C1253 VDPWR.n873 0 0.020442f
C1254 VDPWR.n874 0 0.015494f
C1255 VDPWR.n875 0 0.015494f
C1256 VDPWR.n878 0 0.097351f
C1257 VDPWR.n880 0 0.019496f
C1258 VDPWR.t327 0 0.042905f
C1259 VDPWR.n881 0 0.016874f
C1260 VDPWR.n882 0 0.011749f
C1261 VDPWR.n883 0 0.024888f
C1262 VDPWR.n884 0 0.035465f
C1263 VDPWR.n891 0 0.024888f
C1264 VDPWR.n892 0 0.033299f
C1265 VDPWR.n899 0 0.024888f
C1266 VDPWR.n900 0 0.035021f
C1267 VDPWR.n905 0 0.010629f
C1268 VDPWR.n917 0 0.035021f
C1269 VDPWR.n923 0 0.035021f
C1270 VDPWR.n926 0 0.065056f
C1271 VDPWR.n927 0 0.167187f
C1272 VDPWR.n928 0 0.060534f
C1273 VDPWR.n930 0 0.020792f
C1274 VDPWR.n932 0 0.015494f
C1275 VDPWR.t26 0 0.024205f
C1276 VDPWR.n934 0 0.020442f
C1277 VDPWR.t25 0 0.253491f
C1278 VDPWR.n936 0 0.208129f
C1279 VDPWR.t97 0 0.274837f
C1280 VDPWR.t32 0 0.242818f
C1281 VDPWR.n937 0 0.208129f
C1282 VDPWR.t58 0 0.208129f
C1283 VDPWR.n938 0 0.208129f
C1284 VDPWR.t147 0 0.208129f
C1285 VDPWR.n939 0 0.226808f
C1286 VDPWR.n940 0 0.146758f
C1287 VDPWR.t140 0 0.072045f
C1288 VDPWR.t207 0 0.072045f
C1289 VDPWR.n941 0 0.104065f
C1290 VDPWR.n942 0 0.104065f
C1291 VDPWR.t127 0 0.072045f
C1292 VDPWR.t392 0 0.072045f
C1293 VDPWR.n943 0 0.104065f
C1294 VDPWR.n944 0 0.104065f
C1295 VDPWR.t396 0 0.066708f
C1296 VDPWR.t368 0 0.06404f
C1297 VDPWR.t234 0 0.072045f
C1298 VDPWR.n945 0 0.141421f
C1299 VDPWR.n946 0 0.146758f
C1300 VDPWR.t223 0 0.130748f
C1301 VDPWR.t86 0 0.277506f
C1302 VDPWR.t216 0 0.277506f
C1303 VDPWR.t245 0 0.130748f
C1304 VDPWR.n947 0 0.14409f
C1305 VDPWR.n949 0 0.018877f
C1306 VDPWR.n950 0 0.010329f
C1307 VDPWR.n961 0 0.054638f
C1308 VDPWR.n962 0 2.86136f
C1309 VDPWR.n963 0 0.03443f
C1310 VDPWR.n964 0 2.97888f
C1311 VDPWR.n965 0 0.03443f
C1312 VDPWR.n967 0 0.03443f
C1313 VDPWR.n969 0 0.03443f
C1314 VDPWR.n970 0 0.03443f
C1315 VDPWR.n971 0 5.835f
C1316 VDPWR.n972 0 5.91335f
.ends

