** sch_path: /foss/designs/TTSKY25a-PLL/mag/tb_project_magic.sch
**.subckt tb_project_magic
V1 VDD GND 1.8
V2 ua[0] GND pulse(0 1.8 12ns 1ns 1ns 24ns 50ns)
x1 ua[1] VDD GND ua[0] project_3
**** begin user architecture code
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt



* .include /foss/designs/TTSKY25a-PLL/mag/project_magic.spice
.include /foss/designs/TTSKY25a-PLL/mag/project_3.spice

.option method=gear
* .option method=trap
.option wnflag=1
* .option savecurrents
* .options RSHUNT=1e15
* .options RSHUNT

.save
+v(ua[0])
+v(ua[1])
+v(x1.v_cont.n0)
+v(x1.v_cont.t0)
+v(x1.ua[0].n0)
+v(x1.ua[0].t0)
+v(x1.ua[1].n0)
+v(x1.ua[1].t0)
+@m.x1.x12.msky130_fd_pr__pfet_01v8[id]
+@m.x1.x47.msky130_fd_pr__pfet_01v8[id]
+@m.x1.x93.msky130_fd_pr__pfet_01v8[id]
+@m.x1.x110.msky130_fd_pr__pfet_01v8[id]
+@m.x1.x220.msky130_fd_pr__pfet_01v8[id]
+@m.x1.x252.msky130_fd_pr__pfet_01v8[id]
+@m.x1.x296.msky130_fd_pr__pfet_01v8[id]
+@m.x1.x343.msky130_fd_pr__pfet_01v8[id]
+@m.x1.x364.msky130_fd_pr__pfet_01v8[id]
+@m.x1.x428.msky130_fd_pr__pfet_01v8[id]

* V_out initial voltage

.ic v(x1.v_cont.n0) = 0.0


.control
  * save v(v_osc)

  * timestep for exact simulation results
  tran 5ps 5us


  remzerovec
  * write tb_project_magic_2.raw
  * write tb_project_magic_3.raw
  * write tb_project_magic_4.raw
  * write tb_project_magic_5.raw
  * write tb_project_magic_6.raw
  * write tb_project_magic_7.raw
  * write tb_project_magic_8.raw
  * write tb_project_magic_9.raw
  * write tb_project_magic_10.raw
  * write tb_project_magic_11.raw
  * write tb_project_magic_12.raw
  * write tb_project_magic_13.raw
  * write tb_project_magic_14.raw
  * write tb_project_magic_15.raw
  * write tb_project_magic_16.raw
  * write tb_project_magic_17.raw
  * write tb_project_magic_18.raw
  write tb_project_magic_19.raw
  wrdata /foss/designs/TTSKY25a-PLL/mag/tb_project_magic_v_osc.txt v(x1.ua[1].n0)

  set appendwrite

.endc



**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
