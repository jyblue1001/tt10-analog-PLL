* NGSPICE file created from project_magic.ext - technology: sky130A

.subckt pll_bgr_magic_flat a_8430_7380# a_1930_4410# w_390_7590# a_11910_970# w_1393_10913#
X0 a_3740_7860# a_6460_13890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1 a_700_7870# a_120_13680# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2 w_1393_10913# a_8430_7380# a_13000_1330# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X3 a_2510_6070# a_1870_6040# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X4 a_2850_2700# a_2250_2730# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X5 w_390_7590# w_390_7590# a_1870_6040# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X6 w_1393_10913# a_3230_3880# a_2850_3880# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X7 w_390_7590# a_3870_7600# a_3870_7600# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X8 a_700_7870# a_120_13680# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9 a_6030_1200# a_6140_1280# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X10 w_1393_10913# a_8770_7150# a_6340_3910# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X11 a_3150_3150# a_2250_2730# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X12 w_1393_10913# a_4150_2700# a_3750_2700# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X13 w_390_7590# a_8930_1150# a_8520_1320# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X14 a_3740_7860# a_6460_13890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X15 a_3740_7860# a_670_12430# a_4030_8570# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X16 w_390_7590# a_4150_2700# a_3750_2700# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X17 a_3740_7860# a_6460_13890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X18 w_390_7590# a_830_7600# a_700_7870# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X19 a_9910_990# a_10610_970# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X20 a_8250_7150# a_8250_7150# a_8250_7150# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=5 ps=27 w=1 l=0.15
X21 a_1870_6040# w_390_7590# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X22 w_390_7590# w_390_7590# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=78.005 ps=467.7 w=2 l=0.6
X23 a_1150_10090# a_1870_6040# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X24 a_8610_990# a_9310_970# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X25 a_2330_2700# a_2250_2730# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X26 w_1393_10913# w_1393_10913# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=100.167 ps=594.6 w=2 l=0.6
X27 w_1393_10913# a_2850_3880# a_2330_3880# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X28 a_240_12810# a_1870_6040# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X29 a_2770_3150# a_2250_2730# a_2330_2700# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X30 w_390_7590# a_3870_7600# a_3870_7600# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X31 a_6360_990# a_6140_1280# a_6830_1340# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X32 a_9910_7150# a_11640_6034# w_1393_10913# sky130_fd_pr__res_xhigh_po_0p35 l=1.14
X33 w_1393_10913# a_3050_1280# a_7930_1340# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X34 w_1393_10913# w_1393_10913# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X35 a_240_13888# a_360_12810# w_1393_10913# sky130_fd_pr__res_xhigh_po_0p35 l=3.35
X36 w_1393_10913# a_2020_1290# a_4970_990# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X37 w_390_7590# a_9910_7150# a_6340_3910# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X38 a_1870_6040# w_390_7590# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 w_390_7590# w_390_7590# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0 ps=0 w=2.5 l=0.5
X40 a_4630_3910# a_4190_3910# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X41 a_9620_7120# a_8430_7380# a_8600_8360# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X42 a_700_7870# a_120_13680# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X43 a_1870_6040# w_390_7590# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X44 a_2250_4530# a_2330_3880# a_2250_3910# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X45 a_6340_3910# a_11640_8960# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X46 a_120_13680# a_120_12862# w_1393_10913# sky130_fd_pr__res_high_po_0p35 l=2.05
X47 a_3870_7600# a_2510_6070# a_4030_8570# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X48 a_2510_6070# a_1150_10090# a_1870_6040# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X49 w_390_7590# a_700_7870# a_120_12862# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X50 a_700_7870# a_120_13680# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X51 a_6030_1200# a_6140_1280# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X52 a_9620_7120# a_9620_7120# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X53 a_670_14038# a_670_12430# w_1393_10913# sky130_fd_pr__res_xhigh_po_0p35 l=6
X54 a_700_7870# a_120_13680# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X55 w_390_7590# w_390_7590# a_1870_6040# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X56 w_390_7590# a_3050_1280# a_2020_1290# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X57 w_1393_10913# a_9820_1320# a_9310_970# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X58 w_1393_10913# a_8430_7380# a_12400_1330# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X59 w_1393_10913# w_1393_10913# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X60 w_390_7590# a_9910_990# a_9310_970# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X61 w_1393_10913# w_1393_10913# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X62 a_1870_6040# w_390_7590# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X63 w_390_7590# a_700_7870# a_120_12862# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X64 a_7220_1240# a_6140_1280# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X65 w_1393_10913# a_3630_5470# a_8580_3960# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X66 a_4030_8570# a_2510_6070# a_3870_7600# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X67 w_390_7590# a_2020_1290# a_1760_1030# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X68 a_8430_7380# a_25092_2440# w_1393_10913# sky130_fd_pr__res_xhigh_po_0p35 l=7.52
X69 w_390_7590# a_1870_6040# a_1150_10090# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X70 a_3870_7600# a_3870_7600# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X71 a_6340_3910# a_8770_7150# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X72 w_390_7590# a_3680_910# a_3630_1020# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X73 w_390_7590# w_390_7590# a_240_12810# w_390_7590# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X74 a_3740_7860# a_6460_13890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X75 w_1393_10913# a_8500_8330# a_8500_8330# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X76 w_390_7590# a_120_12862# a_3630_5470# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X77 a_11910_970# a_13110_1020# a_13600_1330# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X78 a_8250_7150# a_8250_7150# a_8250_7150# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X79 a_700_7870# a_120_13680# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X80 a_5790_2730# w_390_7590# a_5400_2730# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X81 a_6470_3910# a_6180_3910# a_6340_3910# w_390_7590# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X82 w_1393_10913# a_8480_7770# a_8770_7150# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X83 a_5790_2730# w_1393_10913# a_5400_2730# w_390_7590# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X84 w_390_7590# a_120_12862# a_1421_8700# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X85 w_390_7590# a_120_12862# a_1421_8700# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X86 w_1393_10913# a_8500_8330# a_8500_8330# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X87 w_1393_10913# a_9910_990# a_9820_1320# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X88 a_1870_6040# w_390_7590# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X89 a_3230_2700# a_2850_2700# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X90 w_1393_10913# a_3750_2700# a_3230_3880# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X91 a_6340_3910# a_9910_7150# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X92 a_3670_3150# a_2850_2700# a_3230_2700# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X93 a_11210_990# a_11910_970# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X94 a_11910_970# a_13110_1020# a_13600_130# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X95 w_1393_10913# a_8770_7150# a_6340_3910# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X96 a_1870_6040# a_3740_7860# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X97 w_1393_10913# a_8500_8330# a_8600_8360# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X98 w_1393_10913# a_6470_2730# a_8430_7380# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X99 a_830_7600# a_240_12810# a_730_9180# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X100 a_1890_1230# a_2020_1290# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X101 a_4810_2700# a_4630_3910# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X102 w_1393_10913# a_8430_7380# sky130_fd_pr__cap_mim_m3_1 l=60 w=13.8
X103 a_8250_7150# a_8580_3960# a_8770_7150# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X104 w_1393_10913# w_1393_10913# a_1570_11090# sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X105 a_7220_1240# a_6140_1280# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X106 a_4030_8570# w_390_7590# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1.01 ps=6.15 w=2.5 l=5
X107 w_1393_10913# a_9310_970# a_10530_1430# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X108 a_8580_3960# a_3630_5470# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X109 a_700_7870# a_120_13680# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X110 a_2940_1200# a_3050_1280# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X111 a_2850_3880# a_3230_3880# a_3150_3910# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X112 a_1870_6040# w_390_7590# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X113 w_1393_10913# a_8010_970# a_9230_1430# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X114 a_2520_1340# a_2020_1290# a_2410_1340# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X115 w_390_7590# a_120_12862# a_3630_5470# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X116 w_390_7590# a_120_12862# a_3630_5470# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X117 w_1393_10913# a_1421_8700# w_1393_10913# sky130_fd_pr__res_xhigh_po_0p35 l=1
X118 a_4030_8570# a_2510_6070# a_3870_7600# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X119 w_1393_10913# w_390_7590# a_1870_6040# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=1.01 pd=6.15 as=1 ps=5.8 w=2.5 l=5
X120 w_390_7590# a_9910_7150# a_6340_3910# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X121 a_830_7600# a_830_7600# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X122 a_5560_14038# a_5440_12430# w_1393_10913# sky130_fd_pr__res_xhigh_po_0p35 l=6
X123 a_7930_1340# a_6140_1280# a_7630_1150# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X124 a_2510_6070# a_1870_6040# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X125 w_390_7590# a_2850_3880# a_2770_3910# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X126 a_4190_4530# a_2330_2700# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X127 a_12480_100# a_12480_100# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X128 a_3850_1340# a_2020_1290# a_3520_1340# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X129 a_700_7870# a_120_13680# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X130 a_3740_7860# a_6460_13890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X131 w_390_7590# a_120_12862# a_1421_8700# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X132 a_8600_8360# a_8500_8330# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X133 a_3740_7860# a_6460_13890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X134 a_830_7600# a_830_7600# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X135 a_7630_1150# a_3050_1280# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X136 w_1393_10913# a_790_12430# w_1393_10913# sky130_fd_pr__res_xhigh_po_0p35 l=6
X137 a_4260_1240# a_3050_1280# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X138 a_8430_7380# a_6470_2730# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X139 a_1890_1230# a_2020_1290# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X140 a_240_12810# a_1870_6040# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X141 a_8500_8330# a_8500_8330# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X142 a_1870_6040# w_390_7590# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X143 w_1393_10913# w_1393_10913# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X144 w_390_7590# a_3870_7600# a_3870_7600# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X145 w_1393_10913# w_390_7590# a_730_9180# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X146 w_1393_10913# a_2330_2700# a_2250_2730# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X147 a_8520_1320# a_8610_990# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X148 a_2940_1200# a_3050_1280# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X149 a_8770_7150# a_8480_7770# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X150 a_2250_2730# a_2330_2700# a_2250_3150# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X151 a_1870_6040# w_390_7590# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X152 w_1393_10913# w_390_7590# a_13600_1330# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X153 w_390_7590# a_4780_1340# a_4260_1240# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X154 w_390_7590# a_120_12862# a_3630_5470# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X155 a_730_9180# a_1421_8700# a_700_7870# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X156 a_700_7870# a_120_13680# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X157 w_390_7590# a_7840_8820# a_7840_8820# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X158 a_6340_3910# a_8770_7150# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X159 w_390_7590# a_10230_1150# a_9820_1320# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X160 a_1870_6040# w_390_7590# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X161 w_1393_10913# a_1760_1030# a_3520_1340# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X162 w_390_7590# a_120_12862# a_1421_8700# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X163 a_700_7870# a_120_13680# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X164 a_6030_1200# a_6360_990# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X165 a_700_7870# a_830_7600# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X166 a_8770_7150# a_8580_3960# a_8250_7150# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X167 w_1393_10913# a_11210_990# a_11120_1320# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X168 w_390_7590# a_7840_8820# a_7840_8820# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X169 a_730_9180# a_240_12810# a_830_7600# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X170 a_6180_3910# a_5790_3910# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X171 a_700_7870# a_120_13680# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X172 w_1393_10913# w_1393_10913# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X173 a_6720_1340# a_5670_990# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X174 a_5400_3910# a_2330_3880# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X175 a_3740_7860# a_670_12430# a_4030_8570# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X176 w_1393_10913# a_4480_2700# a_4150_2700# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X177 a_1421_8700# a_120_12862# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X178 a_6340_3910# a_9910_7150# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X179 a_3740_7860# a_6460_13890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X180 a_8520_1320# a_8610_990# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X181 w_390_7590# a_4480_2700# a_4150_2700# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X182 a_2250_4530# a_1930_4410# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X183 w_390_7590# a_8010_970# a_6140_1280# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X184 a_8600_8360# a_8600_8360# a_8600_8360# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=2.5 ps=17 w=0.5 l=0.15
X185 a_7840_8820# a_8500_8330# sky130_fd_pr__res_generic_po w=0.33 l=2.4
X186 a_4970_990# a_2020_1290# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X187 a_3740_7860# a_6460_13890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X188 w_1393_10913# a_10610_970# a_11830_1430# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X189 a_6470_2730# a_6180_2730# a_3630_5470# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X190 a_3230_10090# a_1150_10090# a_1150_10090# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X191 w_390_7590# a_830_7600# a_830_7600# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X192 a_6470_2730# a_5790_2730# a_3630_5470# w_390_7590# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X193 w_390_7590# a_120_12862# a_3630_5470# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X194 w_390_7590# a_1870_6040# a_240_12810# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X195 w_390_7590# a_3750_2700# a_3670_3910# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X196 a_3050_1280# a_5670_990# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X197 w_390_7590# a_700_7870# a_120_12862# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X198 w_1393_10913# w_1393_10913# a_1570_11090# sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X199 a_1870_6040# w_390_7590# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X200 w_1393_10913# a_4970_990# a_4890_1340# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X201 a_8580_3960# a_6340_3910# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X202 a_4810_2700# a_4630_3910# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X203 w_390_7590# a_120_12862# a_1421_8700# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X204 w_1393_10913# a_1760_1030# a_2520_1340# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X205 w_390_7590# w_390_7590# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X206 w_1393_10913# a_11120_1320# a_10610_970# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X207 a_3630_5470# a_120_12862# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X208 w_390_7590# a_830_7600# a_830_7600# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X209 w_390_7590# a_11210_990# a_10610_970# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X210 w_390_7590# a_1870_6040# a_2510_6070# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X211 w_1393_10913# a_8480_7770# a_8480_7770# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X212 a_8600_8360# a_8600_8360# a_8600_8360# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X213 w_1393_10913# a_3230_2700# a_2850_2700# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X214 a_8250_7150# a_7840_8820# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X215 a_1870_6040# a_3740_7860# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X216 w_1393_10913# w_1393_10913# a_2510_6070# sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X217 a_2850_2700# a_3230_2700# a_3150_3150# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X218 a_240_12810# w_390_7590# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X219 a_1870_6040# w_390_7590# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X220 w_1393_10913# a_360_12810# w_1393_10913# sky130_fd_pr__res_xhigh_po_0p35 l=3.35
X221 w_390_7590# a_830_7600# a_700_7870# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X222 a_4190_3910# a_2330_2700# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.805 ps=5 w=2 l=0.15
X223 w_1393_10913# w_1393_10913# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X224 a_830_7600# a_240_12810# a_730_9180# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X225 w_390_7590# w_1393_10913# a_13000_130# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X226 w_1393_10913# a_2850_2700# a_2330_2700# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X227 a_6470_3910# a_5790_3910# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X228 a_8250_7150# a_8430_7380# a_8480_7770# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X229 w_390_7590# w_390_7590# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X230 w_1393_10913# a_3050_1280# a_4260_1240# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X231 a_3740_7860# a_6460_13890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X232 w_1393_10913# a_1890_1230# a_1760_1030# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X233 w_390_7590# a_2850_2700# a_2770_3150# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X234 a_1870_6040# a_3740_7860# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X235 a_120_12862# w_390_7590# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X236 w_1393_10913# a_4810_2700# a_4480_2700# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X237 a_120_12862# w_390_7590# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X238 a_700_7870# a_120_13680# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X239 a_6140_1280# a_8010_970# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X240 w_390_7590# w_390_7590# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X241 w_390_7590# a_830_7600# a_700_7870# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X242 w_1393_10913# a_2940_1200# a_2020_1290# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X243 w_390_7590# a_4810_2700# a_4480_2700# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X244 w_390_7590# a_11530_1150# a_11120_1320# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X245 w_390_7590# w_390_7590# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X246 a_670_14038# a_790_12430# w_1393_10913# sky130_fd_pr__res_xhigh_po_0p35 l=6
X247 a_700_7870# a_1421_8700# a_730_9180# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X248 w_1393_10913# a_5670_990# a_3050_1280# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X249 w_1393_10913# w_1393_10913# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X250 a_3740_7860# a_6460_13890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X251 a_8600_8360# a_8580_3960# a_9910_7150# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X252 w_390_7590# w_1393_10913# a_12400_130# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X253 w_1393_10913# a_8430_7380# a_13600_1330# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X254 a_4030_8570# a_670_12430# a_3740_7860# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X255 a_11210_990# a_11910_970# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X256 w_390_7590# a_7840_8820# a_8250_7150# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X257 a_1870_6040# a_1150_10090# a_2510_6070# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X258 a_2850_3880# a_2250_4530# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X259 w_1393_10913# a_6140_1280# a_6030_1200# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X260 a_3740_7860# a_6460_13890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X261 a_1150_10090# a_1870_6040# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X262 a_700_7870# a_830_7600# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X263 w_390_7590# a_10610_970# a_9910_990# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X264 a_3740_7860# a_3870_7600# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X265 w_390_7590# a_12480_100# a_13000_130# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X266 a_2940_1200# a_3270_990# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X267 a_1870_6040# w_390_7590# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X268 a_9820_1320# a_9910_990# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X269 a_830_7600# a_830_7600# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X270 w_390_7590# a_9310_970# a_8610_990# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X271 w_390_7590# a_2410_1340# a_1890_1230# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X272 a_2330_3880# a_2250_4530# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X273 w_390_7590# a_1870_6040# a_240_12810# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X274 w_390_7590# a_3740_7860# a_1870_6040# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X275 w_390_7590# a_9620_7120# a_9910_7150# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X276 a_1870_6040# w_390_7590# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X277 a_6830_1340# a_6800_990# a_6720_1340# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X278 a_6470_2730# a_6180_2730# sky130_fd_pr__cap_mim_m3_1 l=3.8 w=2.7
X279 a_830_7600# a_240_12810# a_730_9180# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X280 w_390_7590# a_6470_3910# a_8430_7380# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X281 a_6180_3910# a_5790_3910# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X282 w_390_7590# w_390_7590# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X283 a_5400_3910# a_2330_3880# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X284 a_700_7870# a_120_13680# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X285 a_6340_3910# a_11640_6034# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X286 a_3270_990# a_2020_1290# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X287 w_390_7590# a_12480_100# a_12400_130# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X288 a_2250_3910# a_1930_4410# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X289 a_13110_1020# a_12510_1020# a_13000_1330# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X290 w_390_7590# a_1870_6040# a_2510_6070# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X291 w_390_7590# a_3740_7860# a_1870_6040# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X292 a_700_7870# a_120_13680# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X293 a_240_13888# a_240_12810# w_1393_10913# sky130_fd_pr__res_xhigh_po_0p35 l=3.35
X294 a_1870_6040# w_390_7590# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.45 ps=2.9 w=1 l=0.15
X295 w_1393_10913# w_1393_10913# a_1570_11090# sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X296 w_1393_10913# a_6030_1200# a_5670_990# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X297 a_1421_8700# a_120_12862# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X298 a_3740_7860# a_6460_13890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X299 a_9820_1320# a_9910_990# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X300 w_1393_10913# a_3750_2700# a_3230_2700# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X301 a_730_9180# a_240_12810# a_830_7600# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X302 a_3740_7860# a_6460_13890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X303 w_390_7590# a_3750_2700# a_3670_3150# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X304 a_13110_1020# a_12510_1020# a_13000_130# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X305 a_3740_7860# a_6460_13890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X306 w_390_7590# a_3740_7860# a_1870_6040# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X307 a_8500_8330# a_8500_8330# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X308 a_120_12862# a_700_7870# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X309 a_1870_6040# w_390_7590# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X310 w_1393_10913# a_6140_1280# a_7220_1240# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X311 a_5560_14038# a_2510_6070# w_1393_10913# sky130_fd_pr__res_xhigh_po_0p35 l=6
X312 a_9910_990# a_10610_970# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X313 a_8430_7380# a_6470_3910# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X314 a_1870_6040# w_390_7590# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X315 a_730_9180# a_1421_8700# a_700_7870# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X316 a_8610_990# a_9310_970# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X317 w_390_7590# a_6340_3910# a_8580_3960# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X318 w_390_7590# a_3870_7600# a_3740_7860# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X319 w_1393_10913# w_1393_10913# a_1570_11090# sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X320 a_3630_1020# a_1760_1030# a_3270_990# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X321 a_8600_8360# a_8500_8330# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X322 w_390_7590# w_1393_10913# a_13600_130# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X323 a_3630_5470# a_120_12862# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X324 a_6460_13890# a_1870_6040# w_1393_10913# sky130_fd_pr__res_high_po_0p35 l=2.05
X325 a_3870_7600# a_2510_6070# a_4030_8570# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X326 a_12480_100# a_8430_7380# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X327 a_700_7870# a_120_13680# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 a_5790_3910# a_5400_3910# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X329 a_730_9180# a_1421_8700# a_700_7870# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X330 a_4190_3910# a_2330_3880# a_4190_4530# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X331 a_3270_990# a_3050_1280# a_3850_1340# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X332 a_1421_8700# w_390_7590# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X333 a_700_7870# a_120_13680# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X334 a_1421_8700# a_120_12862# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X335 w_390_7590# a_5670_990# a_6360_990# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X336 a_6470_2730# a_5790_2730# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X337 w_390_7590# a_3870_7600# a_3740_7860# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X338 w_390_7590# a_830_7600# a_830_7600# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X339 a_3230_3880# a_2850_3880# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X340 a_670_12430# a_1870_6040# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X341 a_12510_1020# a_11910_970# a_12400_1330# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X342 a_3740_7860# a_3870_7600# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X343 a_3740_7860# a_670_12430# a_4030_8570# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X344 a_3740_7860# a_6460_13890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X345 w_390_7590# a_11910_970# a_11210_990# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X346 a_3740_7860# a_6460_13890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X347 w_1393_10913# a_2020_1290# a_1890_1230# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X348 w_1393_10913# a_3230_10090# a_3230_10090# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X349 w_1393_10913# w_1393_10913# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.625 pd=3.5 as=0 ps=0 w=1.25 l=0.5
X350 w_390_7590# a_6140_1280# a_6800_990# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X351 w_1393_10913# a_7220_1240# a_6800_990# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X352 a_1570_11090# a_670_12430# w_1393_10913# sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X353 a_10530_1430# a_9910_990# a_10230_1150# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X354 w_390_7590# a_6470_3910# a_8430_7380# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X355 w_1393_10913# a_3050_1280# a_2940_1200# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X356 a_3150_3910# a_2250_4530# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X357 w_390_7590# a_6340_3910# a_8580_3960# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X358 a_9230_1430# a_8610_990# a_8930_1150# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X359 a_3740_7860# a_6460_13890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X360 a_670_12430# a_1870_6040# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X361 w_390_7590# a_12480_100# a_13600_130# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X362 w_1393_10913# w_390_7590# a_13000_1330# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X363 a_12510_1020# a_11910_970# a_12400_130# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X364 a_4780_1340# a_4970_990# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X365 a_9910_7150# a_8580_3960# a_8600_8360# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X366 a_3630_5470# w_390_7590# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X367 a_3740_7860# a_3870_7600# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X368 a_2410_1340# a_1760_1030# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X369 a_3630_5470# a_120_12862# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X370 w_1393_10913# a_8500_8330# a_8600_8360# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X371 a_1870_6040# w_390_7590# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X372 a_10230_1150# a_9310_970# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X373 a_2770_3910# a_2250_4530# a_2330_3880# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X374 a_3520_1340# a_3680_910# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X375 a_700_7870# a_1421_8700# a_730_9180# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X376 a_3740_7860# a_6460_13890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X377 a_1421_8700# a_120_12862# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X378 a_8930_1150# a_8010_970# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X379 a_11120_1320# a_11210_990# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X380 a_700_7870# a_120_13680# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X381 a_9910_7150# a_9620_7120# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X382 a_7840_8820# a_7840_8820# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X383 w_1393_10913# a_5440_12430# w_1393_10913# sky130_fd_pr__res_xhigh_po_0p35 l=6
X384 a_6180_2730# a_5790_2730# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X385 w_390_7590# w_390_7590# a_120_12862# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X386 w_390_7590# a_7630_1150# a_7220_1240# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X387 w_1393_10913# w_1393_10913# a_1570_11090# sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X388 w_1393_10913# a_4260_1240# a_3680_910# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X389 a_5400_2730# a_2330_2700# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X390 a_6180_2730# a_5790_2730# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X391 a_4630_3910# a_4190_3910# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X392 w_1393_10913# a_25092_2440# sky130_fd_pr__cap_mim_m3_1 l=60 w=69.8
X393 a_8480_7770# a_8480_7770# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X394 a_1870_6040# w_390_7590# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X395 a_5400_2730# a_2330_2700# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X396 w_390_7590# w_390_7590# a_1421_8700# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X397 a_3870_7600# a_3870_7600# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X398 w_390_7590# a_1870_6040# a_670_12430# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X399 a_2250_2730# a_1760_1030# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X400 w_1393_10913# a_8610_990# a_8520_1320# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X401 a_8580_3960# a_6340_3910# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X402 w_1393_10913# a_2330_3880# a_2250_4530# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X403 a_7840_8820# a_7840_8820# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X404 a_6140_1280# a_8010_970# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X405 a_1870_6040# w_390_7590# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X406 a_2250_3150# a_1760_1030# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X407 a_4030_8570# a_2510_6070# a_3870_7600# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X408 a_700_7870# a_830_7600# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X409 a_3630_5470# a_120_12862# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X410 w_1393_10913# w_1393_10913# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X411 w_1393_10913# a_3630_5470# a_3630_5470# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X412 w_1393_10913# w_1393_10913# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0 ps=0 w=1.25 l=0.5
X413 w_390_7590# a_5670_990# a_3050_1280# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X414 w_1393_10913# w_1393_10913# a_1570_11090# sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X415 a_700_7870# a_120_13680# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X416 a_8250_7150# a_7840_8820# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X417 w_390_7590# a_1870_6040# a_670_12430# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X418 a_3870_7600# a_3870_7600# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X419 a_8480_7770# a_8430_7380# a_8250_7150# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X420 w_390_7590# a_3050_1280# a_3680_910# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X421 a_1421_8700# a_120_12862# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X422 a_700_7870# a_120_13680# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X423 w_1393_10913# w_1393_10913# a_1570_11090# sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X424 w_1393_10913# w_390_7590# a_12400_1330# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X425 w_390_7590# a_6140_1280# a_5670_990# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X426 w_390_7590# a_3870_7600# a_3740_7860# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X427 a_3740_7860# a_6460_13890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X428 a_11120_1320# a_11210_990# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X429 w_390_7590# w_390_7590# a_3630_5470# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X430 a_3740_7860# a_6460_13890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X431 w_390_7590# w_390_7590# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X432 a_11640_8960# a_8770_7150# w_1393_10913# sky130_fd_pr__res_xhigh_po_0p35 l=0.86
X433 a_8600_8360# a_8430_7380# a_9620_7120# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X434 w_390_7590# a_1870_6040# a_1150_10090# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X435 a_4030_8570# a_670_12430# a_3740_7860# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X436 a_5790_3910# a_5400_3910# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X437 a_120_12862# a_700_7870# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X438 a_6360_990# a_6800_990# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X439 w_1393_10913# w_1393_10913# a_1570_11090# sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X440 w_1393_10913# a_8520_1320# a_8010_970# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X441 w_390_7590# w_390_7590# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X442 w_390_7590# a_2330_3880# a_4190_3910# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X443 w_390_7590# a_8610_990# a_8010_970# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X444 w_390_7590# a_2020_1290# a_4970_990# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X445 a_11830_1430# a_11210_990# a_11530_1150# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X446 w_390_7590# w_390_7590# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=1.25 pd=6 as=0 ps=0 w=2.5 l=0.5
X447 a_1870_6040# w_390_7590# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X448 a_6470_3910# a_5790_3910# a_6340_3910# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X449 a_8430_7380# a_6470_3910# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X450 a_3630_5470# a_120_12862# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X451 a_3630_5470# a_3630_5470# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X452 a_3670_3910# a_2850_3880# a_3230_3880# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X453 a_4260_1240# a_3050_1280# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X454 a_1870_6040# w_390_7590# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X455 w_390_7590# a_9620_7120# a_9620_7120# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X456 a_6470_3910# a_6180_3910# sky130_fd_pr__cap_mim_m3_1 l=6.3 w=5.2
X457 a_1870_6040# w_390_7590# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X458 a_120_12862# a_700_7870# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X459 w_390_7590# a_7840_8820# a_8250_7150# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X460 a_4890_1340# a_3050_1280# a_4780_1340# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X461 a_11530_1150# a_10610_970# w_390_7590# w_390_7590# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X462 a_700_7870# a_120_13680# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X463 w_1393_10913# w_1393_10913# w_1393_10913# w_1393_10913# sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
.ends

** .subckt project_magic ua[0] ua[1] VDPWR VGND
Xpll_bgr_magic_flat_0 V_CONT ua[0] VDPWR ua[1] VSUBS pll_bgr_magic_flat
** .ends

