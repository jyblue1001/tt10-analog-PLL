magic
tech sky130A
timestamp 1756893079
<< metal1 >>
rect 13040 9750 13240 9755
rect 13040 9720 13050 9750
rect 13080 9720 13100 9750
rect 13130 9720 13155 9750
rect 13185 9720 13205 9750
rect 13235 9720 13240 9750
rect 13040 4385 13240 9720
rect 13040 4355 13045 4385
rect 13075 4355 13085 4385
rect 13115 4355 13125 4385
rect 13155 4355 13165 4385
rect 13195 4355 13205 4385
rect 13235 4355 13240 4385
rect 13040 4345 13240 4355
rect 13040 4315 13045 4345
rect 13075 4315 13085 4345
rect 13115 4315 13125 4345
rect 13155 4315 13165 4345
rect 13195 4315 13205 4345
rect 13235 4315 13240 4345
rect 13040 4305 13240 4315
rect 13040 4275 13045 4305
rect 13075 4275 13085 4305
rect 13115 4275 13125 4305
rect 13155 4275 13165 4305
rect 13195 4275 13205 4305
rect 13235 4275 13240 4305
rect 9325 3870 9345 3890
rect 13040 3660 13240 4275
rect 13040 3630 13045 3660
rect 13075 3630 13085 3660
rect 13115 3630 13125 3660
rect 13155 3630 13165 3660
rect 13195 3630 13205 3660
rect 13235 3630 13240 3660
rect 5970 3215 6010 3220
rect 5970 3185 5975 3215
rect 6005 3185 6010 3215
rect 5970 665 6010 3185
rect 13040 1215 13240 3630
rect 13000 1175 13240 1215
rect 13040 1140 13240 1175
rect 13040 1110 13045 1140
rect 13075 1110 13085 1140
rect 13115 1110 13125 1140
rect 13155 1110 13165 1140
rect 13195 1110 13205 1140
rect 13235 1110 13240 1140
rect 13040 1105 13240 1110
rect 5970 635 5975 665
rect 6005 635 6010 665
rect 5970 630 6010 635
<< via1 >>
rect 13050 9720 13080 9750
rect 13100 9720 13130 9750
rect 13155 9720 13185 9750
rect 13205 9720 13235 9750
rect 13045 4355 13075 4385
rect 13085 4355 13115 4385
rect 13125 4355 13155 4385
rect 13165 4355 13195 4385
rect 13205 4355 13235 4385
rect 13045 4315 13075 4345
rect 13085 4315 13115 4345
rect 13125 4315 13155 4345
rect 13165 4315 13195 4345
rect 13205 4315 13235 4345
rect 13045 4275 13075 4305
rect 13085 4275 13115 4305
rect 13125 4275 13155 4305
rect 13165 4275 13195 4305
rect 13205 4275 13235 4305
rect 13045 3630 13075 3660
rect 13085 3630 13115 3660
rect 13125 3630 13155 3660
rect 13165 3630 13195 3660
rect 13205 3630 13235 3660
rect 5975 3185 6005 3215
rect 13045 1110 13075 1140
rect 13085 1110 13115 1140
rect 13125 1110 13155 1140
rect 13165 1110 13195 1140
rect 13205 1110 13235 1140
rect 5975 635 6005 665
<< metal2 >>
rect 3730 9940 3860 9945
rect 3730 9910 3735 9940
rect 3765 9910 3780 9940
rect 3810 9910 3825 9940
rect 3855 9910 3860 9940
rect 3730 9895 3860 9910
rect 3730 9865 3735 9895
rect 3765 9865 3780 9895
rect 3810 9865 3825 9895
rect 3855 9865 3860 9895
rect 3730 9850 3860 9865
rect 3730 9820 3735 9850
rect 3765 9820 3780 9850
rect 3810 9820 3825 9850
rect 3855 9820 3860 9850
rect 3730 9815 3860 9820
rect 12995 9750 13240 9755
rect 12995 9720 13050 9750
rect 13080 9720 13100 9750
rect 13130 9720 13155 9750
rect 13185 9720 13205 9750
rect 13235 9720 13240 9750
rect 12995 9715 13240 9720
rect 3730 9525 4225 9545
rect 3730 9495 3735 9525
rect 3765 9495 3780 9525
rect 3810 9495 3825 9525
rect 3855 9495 4225 9525
rect 3730 9475 4225 9495
rect 3730 9445 3735 9475
rect 3765 9445 3780 9475
rect 3810 9445 3825 9475
rect 3855 9445 4225 9475
rect 3730 9425 4225 9445
rect 6635 4845 6655 4865
rect 13040 4385 13240 4390
rect 13040 4355 13045 4385
rect 13075 4355 13085 4385
rect 13115 4355 13125 4385
rect 13155 4355 13165 4385
rect 13195 4355 13205 4385
rect 13235 4355 13240 4385
rect 13040 4345 13240 4355
rect 13040 4315 13045 4345
rect 13075 4315 13085 4345
rect 13115 4315 13125 4345
rect 13155 4315 13165 4345
rect 13195 4315 13205 4345
rect 13235 4315 13240 4345
rect 13040 4305 13240 4315
rect 13040 4275 13045 4305
rect 13075 4275 13085 4305
rect 13115 4275 13125 4305
rect 13155 4275 13165 4305
rect 13195 4275 13205 4305
rect 13235 4275 13240 4305
rect 13040 4270 13240 4275
rect 13040 3660 13240 3665
rect 13040 3630 13045 3660
rect 13075 3630 13085 3660
rect 13115 3630 13125 3660
rect 13155 3630 13165 3660
rect 13195 3630 13205 3660
rect 13235 3630 13240 3660
rect 13040 3625 13240 3630
rect 5970 3215 6010 3220
rect 5970 3185 5975 3215
rect 6005 3185 6010 3215
rect 5970 3180 6010 3185
rect 12705 1700 13335 1710
rect 12705 1660 13275 1700
rect 13315 1660 13335 1700
rect 12705 1640 13335 1660
rect 12705 1600 13275 1640
rect 13315 1600 13335 1640
rect 12705 1590 13335 1600
rect 13040 1110 13045 1140
rect 13075 1110 13085 1140
rect 13115 1110 13125 1140
rect 13155 1110 13165 1140
rect 13195 1110 13205 1140
rect 13235 1110 13240 1140
rect 13040 1105 13240 1110
rect 15185 670 15265 690
rect 5970 665 15205 670
rect 5970 635 5975 665
rect 6005 635 15205 665
rect 5970 630 15205 635
rect 15245 630 15265 670
rect 15185 610 15265 630
<< via2 >>
rect 3735 9910 3765 9940
rect 3780 9910 3810 9940
rect 3825 9910 3855 9940
rect 3735 9865 3765 9895
rect 3780 9865 3810 9895
rect 3825 9865 3855 9895
rect 3735 9820 3765 9850
rect 3780 9820 3810 9850
rect 3825 9820 3855 9850
rect 3735 9495 3765 9525
rect 3780 9495 3810 9525
rect 3825 9495 3855 9525
rect 3735 9445 3765 9475
rect 3780 9445 3810 9475
rect 3825 9445 3855 9475
rect 13275 1660 13315 1700
rect 13275 1600 13315 1640
rect 15205 630 15245 670
<< metal3 >>
rect 400 9940 3860 9945
rect 400 9930 3735 9940
rect 400 9890 405 9930
rect 445 9890 455 9930
rect 495 9890 505 9930
rect 545 9890 555 9930
rect 595 9910 3735 9930
rect 3765 9910 3780 9940
rect 3810 9910 3825 9940
rect 3855 9910 3860 9940
rect 595 9895 3860 9910
rect 595 9890 3735 9895
rect 400 9870 3735 9890
rect 400 9830 405 9870
rect 445 9830 455 9870
rect 495 9830 505 9870
rect 545 9830 555 9870
rect 595 9865 3735 9870
rect 3765 9865 3780 9895
rect 3810 9865 3825 9895
rect 3855 9865 3860 9895
rect 595 9850 3860 9865
rect 595 9830 3735 9850
rect 400 9820 3735 9830
rect 3765 9820 3780 9850
rect 3810 9820 3825 9850
rect 3855 9820 3860 9850
rect 400 9815 3860 9820
rect 400 9530 3860 9545
rect 400 9490 405 9530
rect 445 9490 455 9530
rect 495 9490 505 9530
rect 545 9490 555 9530
rect 595 9525 3860 9530
rect 595 9495 3735 9525
rect 3765 9495 3780 9525
rect 3810 9495 3825 9525
rect 3855 9495 3860 9525
rect 595 9490 3860 9495
rect 400 9480 3860 9490
rect 400 9440 405 9480
rect 445 9440 455 9480
rect 495 9440 505 9480
rect 545 9440 555 9480
rect 595 9475 3860 9480
rect 595 9445 3735 9475
rect 3765 9445 3780 9475
rect 3810 9445 3825 9475
rect 3855 9445 3860 9475
rect 595 9440 3860 9445
rect 400 9425 3860 9440
rect 100 4505 3860 4520
rect 100 4465 105 4505
rect 145 4465 155 4505
rect 195 4465 205 4505
rect 245 4465 255 4505
rect 295 4465 3860 4505
rect 100 4455 3860 4465
rect 100 4415 105 4455
rect 145 4415 155 4455
rect 195 4415 205 4455
rect 245 4415 255 4455
rect 295 4415 3860 4455
rect 100 4400 3860 4415
rect 400 4355 3860 4370
rect 400 4315 405 4355
rect 445 4315 455 4355
rect 495 4315 505 4355
rect 545 4315 555 4355
rect 595 4315 3860 4355
rect 400 4305 3860 4315
rect 400 4265 405 4305
rect 445 4265 455 4305
rect 495 4265 505 4305
rect 545 4265 555 4305
rect 595 4265 3860 4305
rect 400 4250 3860 4265
rect 400 4180 3860 4195
rect 400 4140 405 4180
rect 445 4140 455 4180
rect 495 4140 505 4180
rect 545 4140 555 4180
rect 595 4140 3860 4180
rect 400 4130 3860 4140
rect 400 4090 405 4130
rect 445 4090 455 4130
rect 495 4090 505 4130
rect 545 4090 555 4130
rect 595 4090 3860 4130
rect 400 4075 3860 4090
rect 100 3590 3860 3605
rect 100 3550 105 3590
rect 145 3550 155 3590
rect 195 3550 205 3590
rect 245 3550 255 3590
rect 295 3550 3860 3590
rect 100 3540 3860 3550
rect 100 3500 105 3540
rect 145 3500 155 3540
rect 195 3500 205 3540
rect 245 3500 255 3540
rect 295 3500 3860 3540
rect 100 3485 3860 3500
rect 400 3000 3860 3015
rect 400 2960 405 3000
rect 445 2960 455 3000
rect 495 2960 505 3000
rect 545 2960 555 3000
rect 595 2960 3860 3000
rect 400 2950 3860 2960
rect 400 2910 405 2950
rect 445 2910 455 2950
rect 495 2910 505 2950
rect 545 2910 555 2950
rect 595 2910 3860 2950
rect 400 2895 3860 2910
rect 100 2850 3860 2865
rect 100 2810 105 2850
rect 145 2810 155 2850
rect 195 2810 205 2850
rect 245 2810 255 2850
rect 295 2810 3860 2850
rect 100 2800 3860 2810
rect 100 2760 105 2800
rect 145 2760 155 2800
rect 195 2760 205 2800
rect 245 2760 255 2800
rect 295 2760 3860 2800
rect 100 2745 3860 2760
rect 100 1900 3860 1915
rect 100 1860 105 1900
rect 145 1860 155 1900
rect 195 1860 205 1900
rect 245 1860 255 1900
rect 295 1860 3860 1900
rect 100 1850 3860 1860
rect 100 1810 105 1850
rect 145 1810 155 1850
rect 195 1810 205 1850
rect 245 1810 255 1850
rect 295 1810 3860 1850
rect 100 1795 3860 1810
rect 13255 1700 13335 1710
rect 13255 1660 13275 1700
rect 13315 1660 13335 1700
rect 13255 1640 13335 1660
rect 13255 1600 13275 1640
rect 13315 1600 13335 1640
rect 13255 1590 13335 1600
rect 400 1510 3860 1525
rect 400 1470 405 1510
rect 445 1470 455 1510
rect 495 1470 505 1510
rect 545 1470 555 1510
rect 595 1470 3860 1510
rect 400 1460 3860 1470
rect 400 1420 405 1460
rect 445 1420 455 1460
rect 495 1420 505 1460
rect 545 1420 555 1460
rect 595 1420 3860 1460
rect 400 1405 3860 1420
rect 400 810 3860 825
rect 400 770 405 810
rect 445 770 455 810
rect 495 770 505 810
rect 545 770 555 810
rect 595 770 3860 810
rect 400 760 3860 770
rect 400 720 405 760
rect 445 720 455 760
rect 495 720 505 760
rect 545 720 555 760
rect 595 720 3860 760
rect 400 705 3860 720
rect 15185 670 15265 690
rect 15185 630 15205 670
rect 15245 630 15265 670
rect 15185 610 15265 630
<< via3 >>
rect 405 9890 445 9930
rect 455 9890 495 9930
rect 505 9890 545 9930
rect 555 9890 595 9930
rect 405 9830 445 9870
rect 455 9830 495 9870
rect 505 9830 545 9870
rect 555 9830 595 9870
rect 405 9490 445 9530
rect 455 9490 495 9530
rect 505 9490 545 9530
rect 555 9490 595 9530
rect 405 9440 445 9480
rect 455 9440 495 9480
rect 505 9440 545 9480
rect 555 9440 595 9480
rect 105 4465 145 4505
rect 155 4465 195 4505
rect 205 4465 245 4505
rect 255 4465 295 4505
rect 105 4415 145 4455
rect 155 4415 195 4455
rect 205 4415 245 4455
rect 255 4415 295 4455
rect 405 4315 445 4355
rect 455 4315 495 4355
rect 505 4315 545 4355
rect 555 4315 595 4355
rect 405 4265 445 4305
rect 455 4265 495 4305
rect 505 4265 545 4305
rect 555 4265 595 4305
rect 405 4140 445 4180
rect 455 4140 495 4180
rect 505 4140 545 4180
rect 555 4140 595 4180
rect 405 4090 445 4130
rect 455 4090 495 4130
rect 505 4090 545 4130
rect 555 4090 595 4130
rect 105 3550 145 3590
rect 155 3550 195 3590
rect 205 3550 245 3590
rect 255 3550 295 3590
rect 105 3500 145 3540
rect 155 3500 195 3540
rect 205 3500 245 3540
rect 255 3500 295 3540
rect 405 2960 445 3000
rect 455 2960 495 3000
rect 505 2960 545 3000
rect 555 2960 595 3000
rect 405 2910 445 2950
rect 455 2910 495 2950
rect 505 2910 545 2950
rect 555 2910 595 2950
rect 105 2810 145 2850
rect 155 2810 195 2850
rect 205 2810 245 2850
rect 255 2810 295 2850
rect 105 2760 145 2800
rect 155 2760 195 2800
rect 205 2760 245 2800
rect 255 2760 295 2800
rect 105 1860 145 1900
rect 155 1860 195 1900
rect 205 1860 245 1900
rect 255 1860 295 1900
rect 105 1810 145 1850
rect 155 1810 195 1850
rect 205 1810 245 1850
rect 255 1810 295 1850
rect 13275 1660 13315 1700
rect 13275 1600 13315 1640
rect 405 1470 445 1510
rect 455 1470 495 1510
rect 505 1470 545 1510
rect 555 1470 595 1510
rect 405 1420 445 1460
rect 455 1420 495 1460
rect 505 1420 545 1460
rect 555 1420 595 1460
rect 405 770 445 810
rect 455 770 495 810
rect 505 770 545 810
rect 555 770 595 810
rect 405 720 445 760
rect 455 720 495 760
rect 505 720 545 760
rect 555 720 595 760
rect 15205 630 15245 670
<< metal4 >>
rect 100 4505 300 22076
rect 100 4465 105 4505
rect 145 4465 155 4505
rect 195 4465 205 4505
rect 245 4465 255 4505
rect 295 4465 300 4505
rect 100 4455 300 4465
rect 100 4415 105 4455
rect 145 4415 155 4455
rect 195 4415 205 4455
rect 245 4415 255 4455
rect 295 4415 300 4455
rect 100 3590 300 4415
rect 100 3550 105 3590
rect 145 3550 155 3590
rect 195 3550 205 3590
rect 245 3550 255 3590
rect 295 3550 300 3590
rect 100 3540 300 3550
rect 100 3500 105 3540
rect 145 3500 155 3540
rect 195 3500 205 3540
rect 245 3500 255 3540
rect 295 3500 300 3540
rect 100 2850 300 3500
rect 100 2810 105 2850
rect 145 2810 155 2850
rect 195 2810 205 2850
rect 245 2810 255 2850
rect 295 2810 300 2850
rect 100 2800 300 2810
rect 100 2760 105 2800
rect 145 2760 155 2800
rect 195 2760 205 2800
rect 245 2760 255 2800
rect 295 2760 300 2800
rect 100 1900 300 2760
rect 100 1860 105 1900
rect 145 1860 155 1900
rect 195 1860 205 1900
rect 245 1860 255 1900
rect 295 1860 300 1900
rect 100 1850 300 1860
rect 100 1810 105 1850
rect 145 1810 155 1850
rect 195 1810 205 1850
rect 245 1810 255 1850
rect 295 1810 300 1850
rect 100 500 300 1810
rect 400 9930 600 22076
rect 400 9890 405 9930
rect 445 9890 455 9930
rect 495 9890 505 9930
rect 545 9890 555 9930
rect 595 9890 600 9930
rect 400 9870 600 9890
rect 400 9830 405 9870
rect 445 9830 455 9870
rect 495 9830 505 9870
rect 545 9830 555 9870
rect 595 9830 600 9870
rect 400 9530 600 9830
rect 400 9490 405 9530
rect 445 9490 455 9530
rect 495 9490 505 9530
rect 545 9490 555 9530
rect 595 9490 600 9530
rect 400 9480 600 9490
rect 400 9440 405 9480
rect 445 9440 455 9480
rect 495 9440 505 9480
rect 545 9440 555 9480
rect 595 9440 600 9480
rect 400 4355 600 9440
rect 400 4315 405 4355
rect 445 4315 455 4355
rect 495 4315 505 4355
rect 545 4315 555 4355
rect 595 4315 600 4355
rect 400 4305 600 4315
rect 400 4265 405 4305
rect 445 4265 455 4305
rect 495 4265 505 4305
rect 545 4265 555 4305
rect 595 4265 600 4305
rect 400 4180 600 4265
rect 400 4140 405 4180
rect 445 4140 455 4180
rect 495 4140 505 4180
rect 545 4140 555 4180
rect 595 4140 600 4180
rect 400 4130 600 4140
rect 400 4090 405 4130
rect 445 4090 455 4130
rect 495 4090 505 4130
rect 545 4090 555 4130
rect 595 4090 600 4130
rect 400 3000 600 4090
rect 400 2960 405 3000
rect 445 2960 455 3000
rect 495 2960 505 3000
rect 545 2960 555 3000
rect 595 2960 600 3000
rect 400 2950 600 2960
rect 400 2910 405 2950
rect 445 2910 455 2950
rect 495 2910 505 2950
rect 545 2910 555 2950
rect 595 2910 600 2950
rect 400 1510 600 2910
rect 400 1470 405 1510
rect 445 1470 455 1510
rect 495 1470 505 1510
rect 545 1470 555 1510
rect 595 1470 600 1510
rect 400 1460 600 1470
rect 400 1420 405 1460
rect 445 1420 455 1460
rect 495 1420 505 1460
rect 545 1420 555 1460
rect 595 1420 600 1460
rect 400 810 600 1420
rect 400 770 405 810
rect 445 770 455 810
rect 495 770 505 810
rect 545 770 555 810
rect 595 770 600 810
rect 400 760 600 770
rect 400 720 405 760
rect 445 720 455 760
rect 495 720 505 760
rect 545 720 555 760
rect 595 720 600 760
rect 400 500 600 720
rect 13255 1700 13335 1710
rect 13255 1660 13275 1700
rect 13315 1660 13335 1700
rect 13255 1640 13335 1660
rect 13255 1600 13275 1640
rect 13315 1600 13335 1640
rect 13255 100 13335 1600
rect 15185 670 15265 690
rect 15185 630 15205 670
rect 15245 630 15265 670
rect 15185 100 15265 630
rect 13249 0 13339 100
rect 15181 0 15271 100
use pll_bgr_magic_5_flat  pll_bgr_magic_5_flat_0
timestamp 1756880322
transform 1 0 5995 0 -1 8165
box -2135 -7890 7050 7460
<< labels >>
flabel metal4 s 15181 0 15271 100 0 FreeSans 480 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 13249 0 13339 100 0 FreeSans 480 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 400 500 600 22076 1 FreeSans 200 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 100 500 300 22076 1 FreeSans 200 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal1 13040 1195 13040 1195 3 FreeSans 800 0 400 0 V_CONT
flabel metal1 9325 3880 9325 3880 7 FreeSans 800 0 -400 0 I_IN
flabel metal2 6645 4845 6645 4845 5 FreeSans 800 0 0 -400 PFET_GATE
<< properties >>
string FIXED_BBOX 0 0 16100 22576
<< end >>
