* PEX produced on Sat Aug 30 02:14:21 AM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from project_2.ext - technology: sky130A

.subckt project_2 clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5] ua[6] ua[7] ui_in[0]
+ ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1]
+ uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1]
+ uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1]
+ uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1]
+ uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7] VDPWR VGND
X0 w_23460_23020.t25 w_23460_23020.t22 w_23460_23020.t24 w_23460_23020.t23 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X1 VGND.t209 a_19190_29050.t11 a_14348_27710.t10 VGND.t208 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X2 a_19190_31850.t9 a_19190_31610.t17 VGND.t125 VGND.t124 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X3 VDPWR.t217 a_26300_25010.t3 a_26300_25670.t1 VDPWR.t216 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X4 a_18180_33430.t8 VGND.t334 VDPWR.t210 VDPWR.t209 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X5 a_14348_27710.t14 VGND.t259 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6 a_26640_21760.t1 a_25860_20180.t3 VGND.t120 VGND.t119 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X7 a_23100_30460.t0 a_24280_30060.t2 VGND.t123 VGND.t122 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X8 VDPWR.t235 VDPWR.t288 a_14730_30630.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X9 VDPWR.t299 a_19910_25340.t4 a_19910_25340.t5 VDPWR.t7 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X10 a_20480_25210.t10 a_19910_24200.t6 a_19040_22530.t4 w_20440_23530.t29 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X11 w_20440_23530.t33 a_17884_25798.t9 a_20480_25210.t11 w_20440_23530.t32 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X12 VGND.t193 a_26320_28790.t2 a_26420_30200.t1 VGND.t192 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X13 a_19190_29050.t12 a_13532_27710.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X14 a_19940_23090.t1 a_23100_27770.t2 a_23130_27670.t1 VDPWR.t184 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X15 a_23100_30980.t1 a_23100_30570.t3 a_23550_30490.t1 VGND.t190 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X16 a_19250_24340.t13 a_17884_25190.t9 VDPWR.t157 VDPWR.t1 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X17 VGND.t51 a_19190_29290.t17 a_19190_29050.t3 VGND.t50 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X18 a_17540_31010.t5 a_14348_27710.t15 VGND.t261 VGND.t260 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X19 VGND.t297 VGND.t295 a_14348_27710.t2 VGND.t296 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X20 VGND.t258 a_14348_27710.t16 a_14730_30630.t6 VGND.t257 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X21 a_14348_27710.t7 VGND.t335 VDPWR.t208 VDPWR.t207 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1.01 ps=6.15 w=2.5 l=5
X22 a_14348_27710.t17 VGND.t256 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X23 a_26420_26340.t0 a_26390_26310.t3 a_26420_26230.t0 VDPWR.t317 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X24 a_14730_30630.t5 a_14348_27710.t18 VGND.t255 VGND.t254 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X25 a_19190_29290.t15 a_14730_30630.t8 a_18180_28430.t10 VDPWR.t171 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X26 VGND.t253 a_14348_27710.t19 a_14990_33500.t5 VGND.t252 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X27 VDPWR.t287 VDPWR.t284 VDPWR.t286 VDPWR.t285 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X28 a_26310_26200.t2 a_26390_27520.t2 VDPWR.t149 VDPWR.t148 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X29 a_24310_31390.t0 a_24280_30570.t3 VGND.t302 VGND.t95 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X30 a_14990_33500.t4 a_14348_27710.t20 VGND.t251 VGND.t250 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X31 a_24280_31090.t1 a_23100_30050.t3 VDPWR.t44 VDPWR.t43 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X32 VGND.t191 a_24280_31090.t3 a_24310_31010.t0 VGND.t58 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X33 VDPWR.t48 a_26390_26310.t4 a_26390_28180.t2 VDPWR.t47 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X34 a_25860_21760.t0 a_19910_24460.t8 VDPWR.t121 VDPWR.t36 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X35 a_19940_24490.t1 a_19910_24460.t9 a_19250_24340.t0 VDPWR.t7 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X36 VGND.t25 a_23100_29610.t3 a_23100_29280.t0 VGND.t24 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X37 a_22190_29430.t17 a_14558_34050.t10 VGND.t19 VGND.t18 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X38 VDPWR.t305 a_17884_25190.t10 a_19250_24340.t12 VDPWR.t1 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X39 VGND.t90 a_19190_29290.t18 a_19190_29050.t5 VGND.t89 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X40 VDPWR.t63 a_23100_30570.t4 a_23100_30980.t2 VDPWR.t62 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X41 w_23460_23020.t7 a_23130_27670.t3 a_19910_24460.t6 w_23460_23020.t6 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X42 a_19190_29290.t11 a_19190_29290.t10 VGND.t29 VGND.t28 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X43 VGND.t73 a_19190_31610.t18 a_19190_31850.t8 VGND.t72 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X44 a_14348_27710.t21 VGND.t247 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X45 a_26300_22300.t1 a_26300_23070.t4 VDPWR.t93 VDPWR.t92 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X46 VDPWR.t124 a_26390_27520.t3 a_26420_27440.t0 VDPWR.t123 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X47 VDPWR.t65 a_26310_26200.t3 a_26390_29930.t2 VDPWR.t64 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X48 a_14348_27710.t22 VGND.t246 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X49 a_20480_25210.t8 a_20480_25210.t6 a_20480_25210.t7 w_20440_23530.t27 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X50 VGND.t27 a_14558_34050.t11 a_14140_28370.t12 VGND.t26 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X51 a_26310_26200.t1 a_26390_27520.t4 VGND.t134 VGND.t133 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X52 a_26390_31270.t2 a_26310_26200.t4 VDPWR.t138 VDPWR.t137 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X53 VDPWR.t115 a_19040_22530.t5 a_19940_23090.t9 VDPWR.t114 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X54 VDPWR.t235 VDPWR.t279 a_13370_29270.t8 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X55 a_24280_31990.t1 a_26320_28790.t3 VGND.t305 VGND.t304 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X56 VDPWR.t21 a_23100_29610.t4 a_23100_29280.t1 VDPWR.t20 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X57 VGND.t75 a_19190_31610.t19 a_19190_31850.t7 VGND.t74 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X58 a_26640_21160.t2 VDPWR.t318 VGND.t6 VGND.t5 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X59 a_19910_24200.t1 a_19940_23090.t10 w_23460_23020.t5 w_23460_23020.t4 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X60 a_22190_29430.t4 a_24280_27770.t2 a_24310_27670.t1 VGND.t108 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X61 a_24280_29730.t0 a_23130_29200.t2 VGND.t65 VGND.t64 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X62 a_26300_23600.t1 a_26300_24370.t4 VDPWR.t23 VDPWR.t22 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X63 a_14558_34050.t8 a_19190_31850.t11 VGND.t49 VGND.t48 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X64 VDPWR.t67 a_26390_30500.t2 a_26420_30420.t1 VDPWR.t66 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X65 VDPWR.t206 VGND.t336 a_14558_34050.t2 VDPWR.t205 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X66 a_14348_27710.t23 VGND.t245 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X67 VGND.t294 VGND.t292 a_14348_27710.t4 VGND.t293 sky130_fd_pr__pfet_01v8 ad=0.45 pd=2.9 as=0.2 ps=1.4 w=1 l=0.15
X68 a_25860_21760.t1 ua[1].t2 a_26400_21130.t0 VDPWR.t36 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X69 a_26420_27220.t1 a_26390_27520.t5 VGND.t47 VGND.t46 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X70 w_20440_23530.t9 a_19940_24490.t4 a_19940_24490.t5 w_20440_23530.t8 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X71 a_26390_32300.t3 a_26320_28790.t4 VDPWR.t191 VDPWR.t190 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X72 a_26320_28790.t0 a_26310_26200.t5 VGND.t21 VGND.t20 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X73 VGND.t121 ua[0].t0 a_23550_31910.t0 VGND.t62 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X74 a_14348_27710.t9 a_19190_29050.t13 VGND.t207 VGND.t206 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X75 VGND.t322 a_23100_29280.t2 a_23130_29200.t0 VGND.t321 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X76 a_19190_31850.t2 a_14140_28370.t13 a_18180_33430.t6 VDPWR.t113 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X77 a_17884_25798.t8 a_17884_25190.t8 VDPWR.t303 sky130_fd_pr__res_xhigh_po_5p73 l=1
X78 VGND.t154 a_19190_29290.t8 a_19190_29290.t9 VGND.t153 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X79 a_26300_24900.t1 a_26300_25670.t4 VDPWR.t233 VDPWR.t232 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X80 a_24280_30980.t0 a_24280_30570.t4 a_24310_30490.t0 VGND.t190 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X81 a_26640_20560.t0 a_26400_20530.t2 ua[1].t0 VGND.t16 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X82 a_14348_27710.t24 VGND.t244 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X83 a_22190_29430.t16 a_14558_34050.t12 VGND.t195 VGND.t194 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X84 VDPWR.t283 VDPWR.t280 VDPWR.t282 VDPWR.t281 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X85 a_26740_30530.t0 a_26390_30500.t3 VGND.t67 VGND.t66 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X86 a_17884_25798.t7 a_17884_25798.t6 w_20440_23530.t15 w_20440_23530.t14 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X87 a_23100_30460.t1 a_24280_30060.t3 VDPWR.t111 VDPWR.t110 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X88 a_14140_28370.t2 VGND.t289 VGND.t291 VGND.t290 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X89 VDPWR.t278 VDPWR.t276 VDPWR.t277 VDPWR.t7 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X90 VGND.t307 a_23100_30050.t4 a_23100_29610.t0 VGND.t306 sky130_fd_pr__pfet_01v8 ad=0.805 pd=5 as=0.4 ps=2.4 w=2 l=0.15
X91 VDPWR.t293 ua[0].t1 a_23020_31090.t0 VDPWR.t292 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X92 a_19190_29050.t14 a_13532_27710.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X93 w_23460_23020.t21 w_23460_23020.t18 w_23460_23020.t20 w_23460_23020.t19 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X94 a_19190_31610.t15 a_19190_31610.t14 VGND.t110 VGND.t109 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X95 VDPWR.t79 a_23100_29280.t3 a_23130_29200.t1 VDPWR.t78 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X96 VDPWR.t51 ua[1].t3 a_26300_22410.t2 VDPWR.t50 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X97 VDPWR.t95 a_26390_26310.t5 a_26390_26970.t3 VDPWR.t94 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X98 VGND.t326 a_19190_31850.t12 a_14558_34050.t7 VGND.t325 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X99 a_14348_27710.t25 VGND.t243 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X100 a_19910_24460.t0 a_25350_8708.t0 VDPWR.t9 sky130_fd_pr__res_xhigh_po_0p35 l=7.52
X101 a_19190_29050.t15 a_13532_27710.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X102 VDPWR.t53 a_24280_27770.t3 a_24310_27670.t2 VDPWR.t52 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X103 a_18180_28430.t1 a_14990_33500.t6 a_19190_29050.t1 VDPWR.t16 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X104 w_20440_23530.t61 w_20440_23530.t58 w_20440_23530.t60 w_20440_23530.t59 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0 ps=0 w=2.5 l=0.5
X105 a_23100_30050.t0 a_24280_30570.t5 VDPWR.t88 VDPWR.t87 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X106 VGND.t288 VGND.t286 a_14140_28370.t1 VGND.t287 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X107 a_19190_31850.t13 a_13742_34050.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X108 a_23100_29610.t1 a_23020_29890.t3 VGND.t53 VGND.t52 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X109 VDPWR.t13 a_24280_31090.t4 a_24280_30570.t0 VDPWR.t12 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X110 a_19190_29050.t16 a_13532_27710.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X111 VGND.t205 a_19190_29050.t17 a_14348_27710.t8 VGND.t204 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X112 VDPWR.t225 a_23100_30050.t5 a_23130_29970.t0 VDPWR.t224 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X113 a_18180_33430.t9 a_14140_28370.t14 a_19190_31850.t10 VDPWR.t302 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X114 VDPWR.t6 a_26300_22300.t2 a_26300_23710.t2 VDPWR.t5 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X115 a_19190_29050.t9 a_19190_29290.t19 VGND.t163 VGND.t162 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X116 a_14348_27710.t26 VGND.t242 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X117 VDPWR.t77 a_26390_26310.t6 a_26390_28180.t1 VDPWR.t76 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X118 a_18180_28430.t3 a_14990_33500.t7 a_19190_29050.t8 VDPWR.t142 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X119 a_13532_33810.t0 a_14610_33690.t1 VDPWR.t189 sky130_fd_pr__res_xhigh_po_0p35 l=3.35
X120 a_19190_29050.t18 a_13532_27710.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X121 a_19910_25340.t3 a_19910_25340.t2 VDPWR.t41 VDPWR.t7 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X122 a_19190_31850.t14 a_13742_34050.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X123 a_19040_22530.t3 a_19910_24200.t7 a_20480_25210.t9 w_20440_23530.t28 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X124 a_19910_24460.t5 a_23130_27670.t4 w_23460_23020.t27 w_23460_23020.t26 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X125 a_26300_23070.t2 a_26300_22410.t3 VDPWR.t188 VDPWR.t187 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X126 a_23130_29970.t1 a_23020_29890.t4 a_23100_29610.t2 VDPWR.t70 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X127 a_26640_21760.t2 VDPWR.t319 VGND.t8 VGND.t7 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X128 a_19190_31850.t15 a_13742_34050.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X129 a_17884_25190.t7 a_17884_25190.t6 VDPWR.t97 VDPWR.t1 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X130 VGND.t12 a_19190_31610.t12 a_19190_31610.t13 VGND.t11 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X131 VDPWR.t311 a_26300_23600.t2 a_26300_25010.t2 VDPWR.t310 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X132 a_24280_30060.t1 a_24280_29730.t2 VGND.t329 VGND.t328 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X133 VGND.t63 a_24280_31990.t2 a_24310_31910.t1 VGND.t62 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X134 a_19190_29050.t19 a_13532_27710.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X135 a_19190_31850.t6 a_19190_31610.t20 VGND.t179 VGND.t178 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X136 a_19910_24460.t2 a_24310_27670.t3 VDPWR.t180 VDPWR.t179 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X137 a_22190_29430.t5 a_24310_27960.t3 a_24310_27670.t0 VDPWR.t153 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X138 a_24280_29730.t1 a_23130_29200.t3 VDPWR.t182 VDPWR.t181 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X139 VGND.t94 a_26420_27220.t3 a_26390_28180.t3 VGND.t93 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X140 a_26390_29240.t2 a_26320_28790.t5 VDPWR.t168 VDPWR.t167 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X141 a_19250_24340.t9 a_19910_24200.t8 a_19940_24230.t4 VDPWR.t7 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X142 w_20440_23530.t57 w_20440_23530.t54 w_20440_23530.t56 w_20440_23530.t55 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X143 a_22190_29430.t15 a_14558_34050.t13 VGND.t132 VGND.t131 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X144 a_19190_29050.t20 a_13532_27710.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X145 a_14140_28370.t11 a_14558_34050.t14 VGND.t148 VGND.t147 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X146 a_19190_31850.t16 a_13742_34050.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X147 VDPWR.t275 VDPWR.t272 VDPWR.t274 VDPWR.t273 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0 ps=0 w=1.25 l=0.5
X148 a_23020_29890.t0 a_23020_31090.t3 a_23550_31390.t0 VGND.t2 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X149 a_13370_29270.t0 a_14990_33500.t1 VDPWR.t135 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X150 a_19190_29290.t7 a_19190_29290.t6 VGND.t23 VGND.t22 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X151 a_18180_28430.t0 a_14990_33500.t8 a_19190_29050.t0 VDPWR.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X152 a_19190_31850.t5 a_19190_31610.t21 VGND.t181 VGND.t180 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X153 a_19190_29050.t21 a_13532_27710.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X154 a_26420_27330.t0 a_26390_26310.t7 a_26420_27220.t0 VDPWR.t290 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X155 VGND.t285 VGND.t283 a_14610_33930.t6 VGND.t284 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X156 VDPWR.t295 a_26310_26200.t6 a_26390_29930.t1 VDPWR.t294 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X157 VDPWR.t119 a_22190_29430.t18 a_19910_24200.t2 VDPWR.t118 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X158 a_19190_29290.t16 a_14730_30630.t9 a_18180_28430.t9 VDPWR.t172 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X159 a_13532_33810.t1 a_14610_33930.t0 VDPWR.t192 sky130_fd_pr__res_xhigh_po_0p35 l=3.35
X160 a_14610_33930.t4 a_14348_27710.t27 VGND.t249 VGND.t248 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X161 a_18180_33430.t1 a_14610_33930.t7 a_19190_31610.t1 VDPWR.t71 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X162 a_20480_25210.t1 a_19910_24460.t10 a_19910_25340.t1 w_20440_23530.t5 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X163 VGND.t241 a_14348_27710.t28 a_17540_31010.t4 VGND.t240 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X164 a_26420_29270.t1 a_26390_29240.t3 VDPWR.t59 VDPWR.t58 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X165 VGND.t57 a_14558_34050.t15 a_22190_29430.t14 VGND.t56 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X166 VDPWR.t161 a_24280_30570.t6 a_24280_30980.t1 VDPWR.t160 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X167 VGND.t185 a_14558_34050.t16 a_14140_28370.t10 VGND.t184 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X168 a_14348_27710.t29 VGND.t220 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X169 a_19940_23090.t8 a_19040_22530.t6 VDPWR.t170 VDPWR.t169 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X170 VGND.t189 a_26320_28790.t6 a_26390_29240.t1 VGND.t188 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X171 a_26330_22330.t0 a_26300_22300.t3 VDPWR.t176 VDPWR.t175 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X172 VDPWR.t27 a_23020_31090.t4 a_23020_29890.t1 VDPWR.t26 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X173 w_23460_23020.t9 a_19940_23090.t11 a_19910_24200.t3 w_23460_23020.t8 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X174 a_14558_34050.t6 a_19190_31850.t17 VGND.t161 VGND.t160 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X175 a_19190_29050.t22 a_13532_27710.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X176 a_26390_27410.t1 a_26390_26970.t4 VDPWR.t106 VDPWR.t105 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X177 a_26300_24370.t2 a_26300_23710.t3 VDPWR.t55 VDPWR.t54 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X178 a_18180_33430.t2 a_14140_28370.t15 a_19190_31850.t0 VDPWR.t80 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X179 a_14730_30630.t2 a_17540_31010.t6 a_14348_27710.t6 VGND.t155 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X180 VDPWR.t320 a_25350_8708.t1 sky130_fd_pr__cap_mim_m3_1 l=69.8 w=60
X181 a_26640_21160.t0 a_26400_21130.t2 a_26400_20530.t0 VGND.t5 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X182 a_19250_24340.t7 a_19250_24340.t5 a_19250_24340.t6 VDPWR.t7 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X183 a_19190_31610.t0 a_14610_33930.t8 a_18180_33430.t0 VDPWR.t60 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X184 a_19940_24490.t3 a_19940_24490.t2 w_20440_23530.t31 w_20440_23530.t30 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X185 a_14348_27710.t30 VGND.t219 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X186 VGND.t107 a_26390_29240.t4 a_26420_29380.t1 VGND.t106 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X187 a_19190_31850.t18 a_13742_34050.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X188 w_20440_23530.t35 a_17884_25798.t10 a_20480_25210.t12 w_20440_23530.t34 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X189 a_26330_23630.t1 a_26300_23600.t3 VDPWR.t102 VDPWR.t101 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X190 VDPWR.t235 VDPWR.t242 a_13370_29270.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X191 VGND.t159 a_26300_22300.t4 a_26330_22440.t0 VGND.t158 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X192 a_19190_29290.t13 a_14730_30630.t10 a_18180_28430.t8 VDPWR.t296 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X193 a_26300_25670.t3 a_26300_25010.t4 VDPWR.t215 VDPWR.t214 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X194 VGND.t152 a_19190_31610.t22 a_19190_31850.t4 VGND.t151 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X195 VGND.t81 ua[1].t4 a_26300_22410.t1 VGND.t80 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X196 a_18180_28430.t7 a_14730_30630.t11 a_19190_29290.t14 VDPWR.t297 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X197 VDPWR.t231 a_19040_22530.t7 a_19940_23090.t7 VDPWR.t230 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X198 a_22190_29430.t7 VGND.t280 VGND.t282 VGND.t281 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X199 VDPWR.t156 a_14610_33690.t0 VDPWR.t155 sky130_fd_pr__res_xhigh_po_0p35 l=3.35
X200 w_20440_23530.t21 a_19940_24230.t5 a_19940_23090.t4 w_20440_23530.t20 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X201 VDPWR.t271 VDPWR.t268 VDPWR.t270 VDPWR.t269 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X202 a_17884_25798.t5 a_17884_25798.t4 w_20440_23530.t3 w_20440_23530.t2 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X203 VDPWR.t185 a_17884_25190.t11 a_19250_24340.t11 VDPWR.t1 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X204 VGND.t112 a_23100_27770.t3 a_23130_27960.t0 VGND.t111 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X205 a_26330_24930.t0 a_26300_24900.t2 VDPWR.t38 VDPWR.t37 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X206 VGND.t43 a_26300_23600.t4 a_26330_23740.t1 VGND.t42 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X207 VDPWR.t235 VDPWR.t243 a_13370_29270.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X208 VGND.t177 a_19190_31850.t19 a_14558_34050.t5 VGND.t176 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X209 a_26300_22300.t0 a_26300_22410.t4 VGND.t37 VGND.t36 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X210 a_19190_31610.t16 a_14610_33930.t9 a_18180_33430.t10 VDPWR.t312 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X211 VGND.t98 a_26300_22300.t5 a_26300_23710.t1 VGND.t97 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X212 a_23100_30050.t1 a_24280_31090.t5 a_24310_31390.t1 VGND.t2 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X213 a_24280_30060.t0 a_24280_29730.t3 VDPWR.t100 VDPWR.t99 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X214 VDPWR.t178 a_24280_31990.t3 a_24280_31090.t2 VDPWR.t177 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X215 a_18180_33430.t4 a_14610_33930.t10 a_19190_31610.t3 VDPWR.t90 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X216 a_19940_23090.t12 a_18460_22530.t1 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X217 a_26390_27520.t1 a_26390_28180.t4 VDPWR.t166 VDPWR.t165 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X218 a_19940_23090.t13 a_21386_22530.t1 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X219 VGND.t10 a_14558_34050.t17 a_22190_29430.t13 VGND.t9 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X220 a_17884_25190.t5 a_17884_25190.t4 VDPWR.t139 VDPWR.t1 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X221 VDPWR.t229 a_23100_27770.t4 a_23130_27960.t1 VDPWR.t228 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X222 VGND.t279 VGND.t277 a_14558_34050.t1 VGND.t278 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X223 a_26300_23600.t0 a_26300_23710.t4 VGND.t129 VGND.t128 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X224 a_18180_28430.t6 a_14730_30630.t12 a_19190_29290.t12 VDPWR.t304 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X225 a_19190_31610.t11 a_19190_31610.t10 VGND.t55 VGND.t54 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X226 a_26390_30500.t1 a_26390_29930.t4 VDPWR.t57 VDPWR.t56 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X227 VGND.t31 a_26300_23600.t5 a_26300_25010.t1 VGND.t30 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X228 a_19190_29050.t10 a_14990_33500.t9 a_18180_28430.t4 VDPWR.t152 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X229 a_26420_31640.t1 a_24280_31990.t4 VDPWR.t141 VDPWR.t140 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X230 a_26390_29240.t0 a_26320_28790.t7 VGND.t35 VGND.t34 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X231 a_19190_29050.t23 a_13532_27710.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X232 w_20440_23530.t53 w_20440_23530.t50 w_20440_23530.t52 w_20440_23530.t51 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X233 a_20480_25210.t5 a_20480_25210.t3 a_20480_25210.t4 w_20440_23530.t26 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X234 a_13742_34050.t20 a_14558_34050.t9 VDPWR.t291 sky130_fd_pr__res_high_po_0p35 l=2.05
X235 a_14140_28370.t9 a_14558_34050.t18 VGND.t39 VGND.t38 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X236 VGND.t301 a_26390_27520.t6 a_26310_26200.t0 VGND.t300 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X237 VDPWR.t35 a_26310_26200.t7 a_26390_31270.t1 VDPWR.t34 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X238 a_14348_27710.t31 VGND.t239 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X239 VGND.t84 a_23100_28450.t2 a_23100_27770.t0 VGND.t15 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X240 a_23550_31010.t1 a_23100_30980.t3 a_23100_30570.t1 VGND.t130 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X241 w_23460_23020.t1 a_23130_27670.t5 a_19910_24460.t4 w_23460_23020.t0 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X242 a_19940_24230.t0 a_21386_22530.t0 VDPWR.t30 sky130_fd_pr__res_xhigh_po_0p35 l=1.14
X243 a_24310_27670.t4 a_24310_27960.t0 sky130_fd_pr__cap_mim_m3_1 l=2.7 w=3.8
X244 a_26300_24900.t0 a_26300_25010.t5 VGND.t14 VGND.t13 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X245 VDPWR.t267 VDPWR.t264 VDPWR.t266 VDPWR.t265 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X246 a_26420_30420.t2 a_24280_31990.t5 VDPWR.t309 VDPWR.t308 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X247 a_26640_21760.t0 ua[1].t5 a_26400_21130.t1 VGND.t7 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X248 VDPWR.t263 VDPWR.t260 VDPWR.t262 VDPWR.t261 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X249 a_18180_33430.t3 a_14610_33930.t11 a_19190_31610.t2 VDPWR.t89 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X250 a_19190_29050.t24 a_13532_27710.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X251 VDPWR.t69 a_26300_24900.t3 a_26390_26310.t0 VDPWR.t68 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X252 VGND.t69 a_26300_24900.t4 a_26330_25040.t0 VGND.t68 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X253 a_19190_31850.t1 a_14140_28370.t16 a_18180_33430.t5 VDPWR.t98 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X254 a_19940_24230.t3 a_19910_24200.t9 a_19250_24340.t8 VDPWR.t8 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X255 VGND.t127 a_24280_31990.t6 a_26420_31750.t1 VGND.t126 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X256 VDPWR.t235 VDPWR.t259 a_13370_29270.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X257 a_14348_27710.t32 VGND.t238 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X258 VDPWR.t151 a_26320_28790.t8 a_26390_32300.t2 VDPWR.t150 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X259 VDPWR.t316 a_23100_28450.t3 a_23100_27770.t1 VDPWR.t315 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X260 a_23100_30570.t0 a_23100_30980.t4 VDPWR.t15 VDPWR.t14 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X261 a_19190_31850.t20 a_13742_34050.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X262 a_26300_22410.t0 ua[1].t6 VGND.t167 VGND.t166 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X263 a_14730_30630.t4 a_14348_27710.t33 VGND.t237 VGND.t236 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X264 a_26390_27410.t0 a_26390_26310.t8 VGND.t157 VGND.t156 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X265 a_19190_29050.t2 a_14990_33500.t10 a_18180_28430.t2 VDPWR.t49 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X266 VGND.t316 a_24280_27770.t4 a_24310_27960.t1 VGND.t111 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X267 VGND.t4 a_19190_31610.t8 a_19190_31610.t9 VGND.t3 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X268 a_19190_29050.t25 a_13532_27710.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X269 a_19910_24200.t4 a_22190_29430.t19 VDPWR.t197 VDPWR.t196 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X270 a_19190_31850.t21 a_13742_34050.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X271 a_19910_25340.t0 a_19910_24460.t11 a_20480_25210.t0 w_20440_23530.t4 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X272 VGND.t88 a_26310_26200.t8 a_26420_26340.t1 VGND.t87 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X273 VGND.t197 a_14558_34050.t19 a_22190_29430.t12 VGND.t196 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X274 VDPWR.t235 VDPWR.t258 a_13370_29270.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X275 a_26420_30200.t2 a_24280_31990.t7 a_26740_30530.t1 VGND.t315 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X276 VGND.t333 a_14558_34050.t20 a_14140_28370.t8 VGND.t332 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X277 VGND.t169 a_26300_24900.t5 a_26390_26310.t2 VGND.t168 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X278 VGND.t71 a_23020_29890.t5 a_23100_28450.t0 VGND.t70 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X279 a_19190_31850.t22 a_13742_34050.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X280 a_26300_23710.t0 a_26300_22300.t6 VGND.t310 VGND.t309 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X281 VDPWR.t257 VDPWR.t254 VDPWR.t256 VDPWR.t255 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X282 a_19910_24200.t0 a_19940_23090.t14 w_23460_23020.t3 w_23460_23020.t2 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X283 a_26390_26970.t2 a_26390_26310.t9 VDPWR.t4 VDPWR.t3 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X284 a_19190_29050.t26 a_13532_27710.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X285 a_19190_31850.t23 a_13742_34050.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X286 VDPWR.t11 a_22190_29430.t2 a_22190_29430.t3 VDPWR.t10 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X287 VDPWR.t29 a_14140_28370.t0 VDPWR.t28 sky130_fd_pr__res_xhigh_po_0p35 l=1
X288 a_19190_31850.t3 a_14140_28370.t17 a_18180_33430.t7 VDPWR.t122 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X289 w_20440_23530.t25 a_19940_24490.t6 a_19940_24230.t2 w_20440_23530.t24 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X290 a_22190_29430.t11 a_14558_34050.t21 VGND.t114 VGND.t113 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X291 a_26420_30310.t0 a_26310_26200.t9 a_26420_30200.t0 VDPWR.t183 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X292 VDPWR.t219 a_24280_31090.t6 a_23100_30050.t2 VDPWR.t218 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X293 a_18460_22530.t0 a_19040_22530.t0 VDPWR.t42 sky130_fd_pr__res_xhigh_po_0p35 l=0.86
X294 a_25860_20560.t2 VGND.t337 VDPWR.t204 VDPWR.t107 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X295 VDPWR.t235 VDPWR.t234 a_13370_29270.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X296 a_19190_29050.t27 a_13532_27710.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X297 VDPWR.t147 a_23020_29890.t6 a_23100_28450.t1 VDPWR.t146 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X298 w_20440_23530.t19 a_17884_25798.t2 a_17884_25798.t3 w_20440_23530.t18 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X299 a_26300_25010.t0 a_26300_23600.t6 VGND.t1 VGND.t0 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X300 a_24310_28480.t3 VDPWR.t321 a_24280_27770.t1 VGND.t15 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X301 a_24310_31010.t1 a_24280_30980.t3 a_24280_30570.t2 VGND.t130 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X302 a_19190_29050.t28 a_13532_27710.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X303 a_26390_28180.t0 a_26390_26310.t10 VDPWR.t19 VDPWR.t18 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X304 a_19190_31850.t24 a_13742_34050.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X305 a_14558_34050.t4 a_19190_31850.t25 VGND.t144 VGND.t143 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X306 a_19940_23090.t6 a_19040_22530.t8 VDPWR.t301 VDPWR.t300 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X307 a_19940_23090.t5 a_19940_24230.t6 w_20440_23530.t23 w_20440_23530.t22 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X308 a_19190_29050.t29 a_13532_27710.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X309 a_20480_25210.t13 a_17884_25798.t11 w_20440_23530.t37 w_20440_23530.t36 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X310 a_19190_31850.t26 a_13742_34050.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X311 a_23550_30490.t0 a_23100_30460.t2 VGND.t327 VGND.t145 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X312 VDPWR.t194 a_26300_22410.t5 a_26300_23070.t3 VDPWR.t193 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X313 VDPWR.t91 a_17884_25190.t2 a_17884_25190.t3 VDPWR.t1 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X314 a_14348_27710.t34 VGND.t218 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X315 w_23460_23020.t17 w_23460_23020.t14 w_23460_23020.t16 w_23460_23020.t15 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X316 a_19190_31850.t27 a_13742_34050.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X317 a_26420_26230.t1 a_26310_26200.t10 VDPWR.t221 VDPWR.t220 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X318 a_26640_20560.t1 a_25860_20180.t4 VGND.t312 VGND.t311 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X319 VDPWR.t174 a_26310_26200.t11 a_26390_31270.t0 VDPWR.t173 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X320 w_20440_23530.t49 w_20440_23530.t46 w_20440_23530.t48 w_20440_23530.t47 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X321 a_26390_27520.t0 a_26390_26310.t11 VGND.t175 VGND.t174 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X322 a_24280_31990.t0 a_26390_32300.t4 VDPWR.t25 VDPWR.t24 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X323 VGND.t173 a_14558_34050.t22 a_22190_29430.t10 VGND.t172 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X324 a_19250_24340.t10 a_17884_25190.t12 VDPWR.t186 VDPWR.t1 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X325 VGND.t140 a_14558_34050.t23 a_14140_28370.t7 VGND.t139 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X326 a_14348_27710.t35 VGND.t217 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X327 a_23100_30980.t0 a_23100_30460.t3 VDPWR.t307 VDPWR.t306 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X328 VGND.t303 a_23100_30050.t6 a_24310_28480.t0 VGND.t70 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X329 a_19190_31850.t28 a_13742_34050.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X330 a_26420_27440.t1 a_26390_27410.t2 a_26420_27330.t1 VDPWR.t314 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X331 a_26390_29930.t0 a_26310_26200.t12 VDPWR.t86 VDPWR.t85 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X332 w_20440_23530.t11 a_19940_24230.t7 a_19940_23090.t2 w_20440_23530.t10 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X333 a_26390_26310.t1 a_26300_24900.t6 VGND.t105 VGND.t104 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X334 VDPWR.t227 a_26320_28790.t9 a_26390_32300.t1 VDPWR.t226 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X335 VDPWR.t82 a_24280_27770.t5 a_24310_27960.t2 VDPWR.t81 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X336 a_26420_29380.t0 a_26310_26200.t13 a_26420_29270.t0 VDPWR.t162 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X337 VGND.t331 a_26420_30200.t3 a_26390_31270.t3 VGND.t330 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X338 a_14140_28370.t6 a_14558_34050.t24 VGND.t142 VGND.t141 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X339 a_25860_20560.t1 a_19910_24460.t12 VDPWR.t136 VDPWR.t107 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X340 VDPWR.t128 a_19910_24460.t13 a_25860_20180.t0 VDPWR.t127 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X341 VDPWR.t313 a_19910_25340.t6 a_19040_22530.t2 VDPWR.t7 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X342 a_26330_22440.t1 a_26300_22410.t6 a_26330_22330.t1 VDPWR.t145 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X343 VGND.t203 a_19190_29050.t30 a_14348_27710.t13 VGND.t202 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X344 VDPWR.t33 a_26300_23710.t5 a_26300_24370.t0 VDPWR.t32 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X345 a_14348_27710.t3 a_17540_31010.t7 a_14730_30630.t1 VGND.t101 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X346 VGND.t324 a_26390_27410.t3 a_26420_27220.t2 VGND.t323 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X347 w_20440_23530.t45 w_20440_23530.t42 w_20440_23530.t44 w_20440_23530.t43 sky130_fd_pr__pfet_01v8 ad=1.25 pd=6 as=0 ps=0 w=2.5 l=0.5
X348 a_26390_29930.t3 a_26420_29380.t2 VGND.t116 VGND.t115 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X349 a_14348_27710.t36 VGND.t216 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X350 a_23550_31910.t1 a_23020_29890.t7 a_23020_31090.t2 VGND.t308 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X351 a_26330_23740.t0 a_26300_23710.t6 a_26330_23630.t0 VDPWR.t298 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X352 a_14610_33930.t3 a_14348_27710.t37 VGND.t235 VGND.t234 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X353 a_26300_23070.t0 a_26330_22440.t2 VGND.t83 VGND.t82 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X354 VGND.t233 a_14348_27710.t38 a_14990_33500.t3 VGND.t232 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X355 VDPWR.t213 a_26300_25010.t6 a_26300_25670.t2 VDPWR.t212 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X356 a_24310_30490.t1 a_23100_30460.t4 VGND.t146 VGND.t145 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X357 a_14990_33500.t2 a_14348_27710.t39 VGND.t222 VGND.t221 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X358 VGND.t231 a_14348_27710.t40 a_14730_30630.t3 VGND.t230 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X359 VDPWR.t253 VDPWR.t250 VDPWR.t252 VDPWR.t251 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X360 a_13382_33380.t0 a_14990_33500.t0 VDPWR.t75 sky130_fd_pr__res_xhigh_po_0p35 l=6
X361 a_25860_20560.t0 a_26400_20530.t3 ua[1].t1 VDPWR.t107 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X362 a_24280_30570.t1 a_24280_30980.t4 VDPWR.t40 VDPWR.t39 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X363 a_24310_28480.t2 VGND.t338 a_24280_27770.t0 VDPWR.t203 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X364 VGND.t61 a_14558_34050.t25 a_22190_29430.t9 VGND.t60 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X365 VDPWR.t249 VDPWR.t247 VDPWR.t248 VDPWR.t7 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X366 w_20440_23530.t17 a_17884_25798.t0 a_17884_25798.t1 w_20440_23530.t16 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X367 a_17540_31010.t1 a_17540_31010.t0 a_17540_28930.t0 VDPWR.t96 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X368 a_25860_21160.t2 VGND.t339 VDPWR.t202 VDPWR.t201 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X369 VDPWR.t246 VDPWR.t244 VDPWR.t245 VDPWR.t1 sky130_fd_pr__nfet_01v8 ad=0.625 pd=3.5 as=0 ps=0 w=1.25 l=0.5
X370 a_13532_27710.t0 a_14348_27710.t5 VDPWR.t112 sky130_fd_pr__res_high_po_0p35 l=2.05
X371 a_19190_29290.t5 a_19190_29290.t4 VGND.t320 VGND.t319 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X372 a_23020_31090.t1 a_23020_29890.t8 VDPWR.t84 VDPWR.t83 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X373 a_19190_29050.t6 a_19190_29290.t20 VGND.t92 VGND.t91 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X374 a_14348_27710.t41 VGND.t229 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X375 VDPWR.t144 a_24310_27670.t5 a_19910_24460.t1 VDPWR.t143 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X376 a_13382_28490.t1 a_14990_28610.t0 VDPWR.t74 sky130_fd_pr__res_xhigh_po_0p35 l=6
X377 a_26640_21160.t1 a_25860_20180.t5 VGND.t314 VGND.t313 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X378 a_26300_24370.t1 a_26330_23740.t2 VGND.t45 VGND.t44 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X379 w_20440_23530.t41 w_20440_23530.t38 w_20440_23530.t40 w_20440_23530.t39 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X380 VGND.t228 a_14348_27710.t42 a_14610_33930.t2 VGND.t227 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X381 a_22190_29430.t1 a_22190_29430.t0 VDPWR.t117 VDPWR.t116 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X382 a_19190_31850.t29 a_13742_34050.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X383 a_19940_24230.t1 a_19940_24490.t7 w_20440_23530.t1 w_20440_23530.t0 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X384 a_23130_27670.t6 a_23130_27960.t2 sky130_fd_pr__cap_mim_m3_1 l=5.2 w=6.3
X385 a_14140_28370.t5 a_14558_34050.t26 VGND.t299 VGND.t298 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X386 a_19250_24340.t1 a_19910_24460.t14 a_19940_24490.t0 VDPWR.t7 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X387 VDPWR.t2 a_17884_25190.t0 a_17884_25190.t1 VDPWR.t1 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X388 a_14348_27710.t43 VGND.t215 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X389 a_14558_34050.t0 VGND.t274 VGND.t276 VGND.t275 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X390 VGND.t318 a_25860_20180.t1 a_25860_20180.t2 VGND.t317 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X391 w_23460_23020.t13 w_23460_23020.t10 w_23460_23020.t12 w_23460_23020.t11 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X392 a_26330_25040.t1 a_26300_25010.t7 a_26330_24930.t1 VDPWR.t211 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X393 VDPWR.t223 a_23100_30050.t7 a_24310_28480.t1 VDPWR.t222 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X394 a_26420_31750.t0 a_26320_28790.t10 a_26420_31640.t0 VDPWR.t31 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X395 a_19190_31850.t30 a_13742_34050.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X396 VDPWR.t164 a_14990_33260.t1 VDPWR.t163 sky130_fd_pr__res_xhigh_po_0p35 l=6
X397 a_26320_28790.t1 a_26390_31270.t4 VDPWR.t159 VDPWR.t158 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X398 a_19190_29050.t31 a_13532_27710.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X399 VDPWR.t104 a_26300_22410.t7 a_26300_23070.t1 VDPWR.t103 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X400 VGND.t100 a_19190_29290.t2 a_19190_29290.t3 VGND.t99 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X401 VGND.t138 a_19190_29290.t21 a_19190_29050.t7 VGND.t137 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X402 w_23460_23020.t31 a_19940_23090.t15 a_19910_24200.t5 w_23460_23020.t30 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X403 a_14348_27710.t1 VGND.t271 VGND.t273 VGND.t272 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X404 VDPWR.t132 a_14990_28610.t1 VDPWR.t131 sky130_fd_pr__res_xhigh_po_0p35 l=6
X405 a_24310_31910.t0 a_23100_30050.t8 a_24280_31090.t0 VGND.t308 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X406 a_19190_31850.t31 a_13742_34050.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X407 VDPWR.t241 VDPWR.t238 VDPWR.t240 VDPWR.t239 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X408 a_26300_25670.t0 a_26330_25040.t2 VGND.t103 VGND.t102 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X409 a_26390_32300.t0 a_26420_31750.t2 VGND.t150 VGND.t149 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X410 a_19190_29050.t32 a_13532_27710.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X411 a_26390_30500.t0 a_26310_26200.t14 VGND.t41 VGND.t40 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X412 a_25860_21160.t0 a_19910_24460.t15 VDPWR.t289 VDPWR.t201 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X413 VGND.t183 a_23100_27770.t5 a_23130_27670.t0 VGND.t182 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X414 VGND.t33 a_14558_34050.t27 a_14140_28370.t4 VGND.t32 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X415 a_14348_27710.t44 VGND.t214 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X416 a_19190_31610.t7 a_19190_31610.t6 VGND.t86 VGND.t85 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X417 a_26640_20560.t2 VDPWR.t322 VGND.t17 VGND.t16 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X418 a_23550_31390.t1 a_23100_30570.t5 VGND.t96 VGND.t95 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X419 a_19190_29050.t33 a_13532_27710.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X420 VDPWR.t200 VGND.t340 a_18180_28430.t5 VDPWR.t199 sky130_fd_pr__nfet_01v8 ad=1.01 pd=6.15 as=1 ps=5.8 w=2.5 l=5
X421 a_14348_27710.t12 a_19190_29050.t34 VGND.t201 VGND.t200 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X422 VGND.t79 a_19190_31850.t32 a_14558_34050.t3 VGND.t78 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X423 VGND.t59 a_23020_31090.t5 a_23550_31010.t0 VGND.t58 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X424 VDPWR.t323 a_19910_24460.t7 sky130_fd_pr__cap_mim_m3_1 l=13.8 w=60
X425 a_19190_31850.t33 a_13742_34050.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X426 VDPWR.t235 VDPWR.t236 a_13370_29270.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X427 a_14348_27710.t45 VGND.t213 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X428 a_19940_23090.t0 a_19940_24230.t8 w_20440_23530.t7 w_20440_23530.t6 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X429 a_26390_26970.t0 a_26420_26340.t2 VGND.t136 VGND.t135 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X430 a_22190_29430.t8 a_14558_34050.t28 VGND.t187 VGND.t186 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X431 a_24280_30980.t2 a_23100_30460.t5 VDPWR.t130 VDPWR.t129 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X432 a_13382_33380.t1 a_14990_33260.t0 VDPWR.t154 sky130_fd_pr__res_xhigh_po_0p35 l=6
X433 a_14140_28370.t3 a_14558_34050.t29 VGND.t171 VGND.t170 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X434 a_19190_31850.t34 a_13742_34050.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X435 a_25860_21760.t2 VGND.t341 VDPWR.t198 VDPWR.t36 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X436 a_19040_22530.t1 a_19910_25340.t7 VDPWR.t195 VDPWR.t7 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X437 a_19190_29050.t35 a_13532_27710.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X438 a_19190_29050.t4 a_19190_29290.t22 VGND.t77 VGND.t76 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X439 a_14348_27710.t11 a_19190_29050.t36 VGND.t199 VGND.t198 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X440 a_19910_24460.t3 a_23130_27670.t7 w_23460_23020.t29 w_23460_23020.t28 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X441 VGND.t226 a_14348_27710.t46 a_17540_31010.t3 VGND.t225 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X442 a_23020_29890.t2 a_23100_30570.t6 VDPWR.t126 VDPWR.t125 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X443 a_19190_31850.t35 a_13742_34050.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X444 VDPWR.t46 a_26390_26310.t12 a_26390_26970.t1 VDPWR.t45 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X445 a_17540_31010.t2 a_14348_27710.t47 VGND.t224 VGND.t223 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X446 VDPWR.t109 a_26300_23710.t7 a_26300_24370.t3 VDPWR.t108 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X447 VGND.t212 a_14348_27710.t48 a_14610_33930.t1 VGND.t211 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X448 VGND.t118 a_19190_29290.t0 a_19190_29290.t1 VGND.t117 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X449 VDPWR.t134 a_23020_31090.t6 a_23100_30570.t2 VDPWR.t133 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X450 VDPWR.t235 VDPWR.t237 a_13370_29270.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X451 a_14348_27710.t49 VGND.t210 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X452 a_14610_33930.t5 VGND.t268 VGND.t270 VGND.t269 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X453 a_13382_28490.t0 a_14730_30630.t0 VDPWR.t17 sky130_fd_pr__res_xhigh_po_0p35 l=6
X454 a_14348_27710.t0 VGND.t265 VGND.t267 VGND.t266 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X455 a_17540_28930.t0 a_17540_28930.t1 VDPWR.t73 VDPWR.t72 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X456 VGND.t264 VGND.t262 a_22190_29430.t6 VGND.t263 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X457 a_25860_21160.t1 a_26400_21130.t3 a_26400_20530.t1 VDPWR.t201 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X458 a_19190_31850.t36 a_13742_34050.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X459 a_26420_30420.t0 a_26320_28790.t11 a_26420_30310.t1 VDPWR.t120 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X460 a_19940_23090.t3 a_23130_27960.t3 a_23130_27670.t2 VGND.t108 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X461 a_19250_24340.t4 a_19250_24340.t2 a_19250_24340.t3 VDPWR.t61 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X462 a_20480_25210.t2 a_17884_25798.t12 w_20440_23530.t13 w_20440_23530.t12 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X463 VGND.t165 a_19190_31610.t4 a_19190_31610.t5 VGND.t164 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
R0 w_23460_23020.n46 w_23460_23020.n45 782
R1 w_23460_23020.n72 w_23460_23020.n24 782
R2 w_23460_23020.n47 w_23460_23020.n24 585
R3 w_23460_23020.n49 w_23460_23020.n46 585
R4 w_23460_23020.n48 w_23460_23020.t12 432.038
R5 w_23460_23020.t12 w_23460_23020.n23 432.038
R6 w_23460_23020.t21 w_23460_23020.n57 431.421
R7 w_23460_23020.n58 w_23460_23020.t21 431.421
R8 w_23460_23020.n41 w_23460_23020.t16 431.421
R9 w_23460_23020.t16 w_23460_23020.n40 431.421
R10 w_23460_23020.t30 w_23460_23020.t15 360.346
R11 w_23460_23020.t4 w_23460_23020.t30 360.346
R12 w_23460_23020.t8 w_23460_23020.t4 360.346
R13 w_23460_23020.t2 w_23460_23020.t8 360.346
R14 w_23460_23020.t23 w_23460_23020.t2 360.346
R15 w_23460_23020.t11 w_23460_23020.t6 360.346
R16 w_23460_23020.t6 w_23460_23020.t26 360.346
R17 w_23460_23020.t26 w_23460_23020.t0 360.346
R18 w_23460_23020.t0 w_23460_23020.t28 360.346
R19 w_23460_23020.t28 w_23460_23020.t19 360.346
R20 w_23460_23020.t15 w_23460_23020.n43 343.966
R21 w_23460_23020.n70 w_23460_23020.t23 343.966
R22 w_23460_23020.n70 w_23460_23020.t11 343.966
R23 w_23460_23020.t19 w_23460_23020.n69 343.966
R24 w_23460_23020.n44 w_23460_23020.t22 336.329
R25 w_23460_23020.n44 w_23460_23020.t10 336.329
R26 w_23460_23020.n36 w_23460_23020.t14 320.7
R27 w_23460_23020.n66 w_23460_23020.t18 320.7
R28 w_23460_23020.n57 w_23460_23020.n52 234.355
R29 w_23460_23020.n72 w_23460_23020.n71 230.308
R30 w_23460_23020.n68 w_23460_23020.n67 230.308
R31 w_23460_23020.n51 w_23460_23020.n45 230.308
R32 w_23460_23020.n64 w_23460_23020.n59 196.502
R33 w_23460_23020.n63 w_23460_23020.n60 196.502
R34 w_23460_23020.n62 w_23460_23020.n61 196.502
R35 w_23460_23020.n31 w_23460_23020.n30 196.502
R36 w_23460_23020.n34 w_23460_23020.n33 196.502
R37 w_23460_23020.n75 w_23460_23020.n74 196.502
R38 w_23460_23020.n42 w_23460_23020.n41 189.048
R39 w_23460_23020.n54 w_23460_23020.n53 185
R40 w_23460_23020.n56 w_23460_23020.n55 185
R41 w_23460_23020.n47 w_23460_23020.n25 185
R42 w_23460_23020.n50 w_23460_23020.n49 185
R43 w_23460_23020.n43 w_23460_23020.n42 185
R44 w_23460_23020.n29 w_23460_23020.n28 185
R45 w_23460_23020.n39 w_23460_23020.n38 185
R46 w_23460_23020.n37 w_23460_23020.n27 185
R47 w_23460_23020.n43 w_23460_23020.n27 185
R48 w_23460_23020.n45 w_23460_23020.n44 166.63
R49 w_23460_23020.n50 w_23460_23020.n25 120.001
R50 w_23460_23020.n55 w_23460_23020.n53 120.001
R51 w_23460_23020.n42 w_23460_23020.n28 120.001
R52 w_23460_23020.n38 w_23460_23020.n27 120.001
R53 w_23460_23020.n46 w_23460_23020.t25 98.5005
R54 w_23460_23020.t25 w_23460_23020.n24 98.5005
R55 w_23460_23020.n69 w_23460_23020.n68 69.8479
R56 w_23460_23020.n69 w_23460_23020.n52 69.8479
R57 w_23460_23020.n71 w_23460_23020.n70 69.8479
R58 w_23460_23020.n70 w_23460_23020.n51 69.8479
R59 w_23460_23020.n43 w_23460_23020.n26 69.8479
R60 w_23460_23020.n51 w_23460_23020.n50 45.3071
R61 w_23460_23020.n55 w_23460_23020.n52 45.3071
R62 w_23460_23020.n68 w_23460_23020.n53 45.3071
R63 w_23460_23020.n71 w_23460_23020.n25 45.3071
R64 w_23460_23020.n28 w_23460_23020.n26 45.3071
R65 w_23460_23020.n38 w_23460_23020.n26 45.3071
R66 w_23460_23020.n73 w_23460_23020.n72 32.2291
R67 w_23460_23020.n21 w_23460_23020.n20 43.7643
R68 w_23460_23020.n64 w_23460_23020.n20 21.8824
R69 w_23460_23020.n17 w_23460_23020.n16 43.7643
R70 w_23460_23020.n63 w_23460_23020.n16 9.08242
R71 w_23460_23020.n73 w_23460_23020.n11 21.8824
R72 w_23460_23020.n5 w_23460_23020.n9 41.0489
R73 w_23460_23020.n32 w_23460_23020.n0 37.8824
R74 w_23460_23020.n0 w_23460_23020.n31 34.6824
R75 w_23460_23020.n74 w_23460_23020.n11 34.6824
R76 w_23460_23020.n59 w_23460_23020.t29 24.6255
R77 w_23460_23020.n59 w_23460_23020.t20 24.6255
R78 w_23460_23020.n60 w_23460_23020.t27 24.6255
R79 w_23460_23020.n60 w_23460_23020.t1 24.6255
R80 w_23460_23020.n61 w_23460_23020.t13 24.6255
R81 w_23460_23020.n61 w_23460_23020.t7 24.6255
R82 w_23460_23020.n30 w_23460_23020.t5 24.6255
R83 w_23460_23020.n30 w_23460_23020.t9 24.6255
R84 w_23460_23020.n33 w_23460_23020.t17 24.6255
R85 w_23460_23020.n33 w_23460_23020.t31 24.6255
R86 w_23460_23020.n75 w_23460_23020.t3 24.6255
R87 w_23460_23020.t24 w_23460_23020.n75 24.6255
R88 w_23460_23020.n66 w_23460_23020.n65 24.361
R89 w_23460_23020.n36 w_23460_23020.n35 22.6157
R90 w_23460_23020.n12 w_23460_23020.n14 42.1635
R91 w_23460_23020.n62 w_23460_23020.n14 5.08198
R92 w_23460_23020.n34 w_23460_23020.n32 22.4005
R93 w_23460_23020.n17 w_23460_23020.n62 21.8824
R94 w_23460_23020.n67 w_23460_23020.n66 15.6449
R95 w_23460_23020.n37 w_23460_23020.n36 15.6449
R96 w_23460_23020.n4 w_23460_23020.n5 41.0489
R97 w_23460_23020.n74 w_23460_23020.n9 3.16696
R98 w_23460_23020.n73 w_23460_23020.n12 5.08198
R99 w_23460_23020.n14 w_23460_23020.n13 2.11051
R100 w_23460_23020.n20 w_23460_23020.n19 1.71029
R101 w_23460_23020.n22 w_23460_23020.n21 1.71029
R102 w_23460_23020.n16 w_23460_23020.n15 1.71029
R103 w_23460_23020.n18 w_23460_23020.n17 1.71029
R104 w_23460_23020.n10 w_23460_23020.n12 2.11051
R105 w_23460_23020.n8 w_23460_23020.n11 1.71029
R106 w_23460_23020.n7 w_23460_23020.n5 1.71029
R107 w_23460_23020.n4 w_23460_23020.n1 3.06802
R108 w_23460_23020.n4 w_23460_23020.n31 3.16696
R109 w_23460_23020.n3 w_23460_23020.n0 1.71029
R110 w_23460_23020.n32 w_23460_23020.n2 9.3005
R111 w_23460_23020.n9 w_23460_23020.n6 3.06802
R112 w_23460_23020.n56 w_23460_23020.n54 7.11161
R113 w_23460_23020.n39 w_23460_23020.n29 7.11161
R114 w_23460_23020.n65 w_23460_23020.n64 6.54033
R115 w_23460_23020.n35 w_23460_23020.n34 6.25084
R116 w_23460_23020.n49 w_23460_23020.n47 4.57193
R117 w_23460_23020.n67 w_23460_23020.n58 4.0479
R118 w_23460_23020.n40 w_23460_23020.n37 4.0479
R119 w_23460_23020.n21 w_23460_23020.n63 9.08242
R120 w_23460_23020.n58 w_23460_23020.n54 3.02841
R121 w_23460_23020.n57 w_23460_23020.n56 3.02841
R122 w_23460_23020.n40 w_23460_23020.n39 3.02841
R123 w_23460_23020.n41 w_23460_23020.n29 3.02841
R124 w_23460_23020.n48 w_23460_23020.n45 2.6074
R125 w_23460_23020.n72 w_23460_23020.n23 2.6074
R126 w_23460_23020.n47 w_23460_23020.n23 1.9508
R127 w_23460_23020.n49 w_23460_23020.n48 1.9508
R128 w_23460_23020.n65 w_23460_23020.n19 0.703395
R129 w_23460_23020.n35 w_23460_23020.n2 0.570933
R130 w_23460_23020.n19 w_23460_23020.n22 0.313
R131 w_23460_23020.n22 w_23460_23020.n15 0.313
R132 w_23460_23020.n15 w_23460_23020.n18 0.313
R133 w_23460_23020.n18 w_23460_23020.n13 0.313
R134 w_23460_23020.n13 w_23460_23020.n10 0.313
R135 w_23460_23020.n8 w_23460_23020.n10 0.313
R136 w_23460_23020.n6 w_23460_23020.n8 0.313
R137 w_23460_23020.n7 w_23460_23020.n6 0.313
R138 w_23460_23020.n7 w_23460_23020.n1 0.313
R139 w_23460_23020.n3 w_23460_23020.n1 0.313
R140 w_23460_23020.n3 w_23460_23020.n2 0.313
R141 a_19190_29050.n4 a_19190_29050.t30 363.909
R142 a_19190_29050.n4 a_19190_29050.t36 351.974
R143 a_19190_29050.n12 a_19190_29050.n4 299.252
R144 a_19190_29050.n4 a_19190_29050.n5 299.25
R145 a_19190_29050.n4 a_19190_29050.n7 299.25
R146 a_19190_29050.n3 a_19190_29050.t8 242.968
R147 a_19190_29050.n10 a_19190_29050.n8 200.477
R148 a_19190_29050.n10 a_19190_29050.n9 199.727
R149 a_19190_29050.n6 a_19190_29050.t17 194.809
R150 a_19190_29050.n6 a_19190_29050.t13 194.809
R151 a_19190_29050.n11 a_19190_29050.t11 194.809
R152 a_19190_29050.n11 a_19190_29050.t34 194.809
R153 a_19190_29050.n4 a_19190_29050.n6 163.097
R154 a_19190_29050.n3 a_19190_29050.n11 161.653
R155 a_19190_29050.n8 a_19190_29050.t1 48.0005
R156 a_19190_29050.n8 a_19190_29050.t2 48.0005
R157 a_19190_29050.n9 a_19190_29050.t0 48.0005
R158 a_19190_29050.n9 a_19190_29050.t10 48.0005
R159 a_19190_29050.n5 a_19190_29050.t7 39.4005
R160 a_19190_29050.n5 a_19190_29050.t6 39.4005
R161 a_19190_29050.n7 a_19190_29050.t5 39.4005
R162 a_19190_29050.n7 a_19190_29050.t9 39.4005
R163 a_19190_29050.t3 a_19190_29050.n12 39.4005
R164 a_19190_29050.n12 a_19190_29050.t4 39.4005
R165 a_19190_29050.n3 a_19190_29050.n10 5.2505
R166 a_19190_29050.n0 a_19190_29050.t18 4.8248
R167 a_19190_29050.n1 a_19190_29050.t12 4.5005
R168 a_19190_29050.n1 a_19190_29050.t21 4.5005
R169 a_19190_29050.n0 a_19190_29050.t27 4.5005
R170 a_19190_29050.n0 a_19190_29050.t22 4.5005
R171 a_19190_29050.n0 a_19190_29050.t29 4.5005
R172 a_19190_29050.n0 a_19190_29050.t33 4.5005
R173 a_19190_29050.n0 a_19190_29050.t15 4.5005
R174 a_19190_29050.n0 a_19190_29050.t35 4.5005
R175 a_19190_29050.n1 a_19190_29050.t25 4.5005
R176 a_19190_29050.n1 a_19190_29050.t19 4.5005
R177 a_19190_29050.n1 a_19190_29050.t20 4.5005
R178 a_19190_29050.n1 a_19190_29050.t26 4.5005
R179 a_19190_29050.n1 a_19190_29050.t31 4.5005
R180 a_19190_29050.n2 a_19190_29050.t28 4.5005
R181 a_19190_29050.n2 a_19190_29050.t32 4.5005
R182 a_19190_29050.n2 a_19190_29050.t14 4.5005
R183 a_19190_29050.n2 a_19190_29050.t23 4.5005
R184 a_19190_29050.n2 a_19190_29050.t16 4.5005
R185 a_19190_29050.n2 a_19190_29050.t24 4.5005
R186 a_19190_29050.n4 a_19190_29050.n2 11.6632
R187 a_19190_29050.n2 a_19190_29050.n1 3.5678
R188 a_19190_29050.n4 a_19190_29050.n3 2.7106
R189 a_19190_29050.n1 a_19190_29050.n0 2.3035
R190 a_14348_27710.n2 a_14348_27710.t27 355.784
R191 a_14348_27710.n8 a_14348_27710.t42 355.502
R192 a_14348_27710.n10 a_14348_27710.t48 354.75
R193 a_14348_27710.n0 a_14348_27710.t37 351.002
R194 a_14348_27710.n2 a_14348_27710.t28 310.401
R195 a_14348_27710.n3 a_14348_27710.t15 310.401
R196 a_14348_27710.n4 a_14348_27710.t16 310.401
R197 a_14348_27710.n5 a_14348_27710.t18 310.401
R198 a_14348_27710.n6 a_14348_27710.t19 310.401
R199 a_14348_27710.n7 a_14348_27710.t20 310.401
R200 a_14348_27710.n14 a_14348_27710.t39 310.401
R201 a_14348_27710.n13 a_14348_27710.t40 310.401
R202 a_14348_27710.n12 a_14348_27710.t33 310.401
R203 a_14348_27710.n11 a_14348_27710.t46 310.401
R204 a_14348_27710.n10 a_14348_27710.t47 310.401
R205 a_14348_27710.n27 a_14348_27710.n26 306.808
R206 a_14348_27710.n1 a_14348_27710.t38 305.901
R207 a_14348_27710.n20 a_14348_27710.n19 301.933
R208 a_14348_27710.n22 a_14348_27710.n21 301.933
R209 a_14348_27710.n24 a_14348_27710.n23 301.933
R210 a_14348_27710.n29 a_14348_27710.n28 297.433
R211 a_14348_27710.n27 a_14348_27710.n25 297.433
R212 a_14348_27710.t5 a_14348_27710.n50 149.127
R213 a_14348_27710.n18 a_14348_27710.t7 98.9207
R214 a_14348_27710.n28 a_14348_27710.t13 39.4005
R215 a_14348_27710.n28 a_14348_27710.t1 39.4005
R216 a_14348_27710.n26 a_14348_27710.t4 39.4005
R217 a_14348_27710.n26 a_14348_27710.t3 39.4005
R218 a_14348_27710.n25 a_14348_27710.t6 39.4005
R219 a_14348_27710.n25 a_14348_27710.t0 39.4005
R220 a_14348_27710.n19 a_14348_27710.t2 39.4005
R221 a_14348_27710.n19 a_14348_27710.t11 39.4005
R222 a_14348_27710.n21 a_14348_27710.t8 39.4005
R223 a_14348_27710.n21 a_14348_27710.t9 39.4005
R224 a_14348_27710.n23 a_14348_27710.t10 39.4005
R225 a_14348_27710.n23 a_14348_27710.t12 39.4005
R226 a_14348_27710.n50 a_14348_27710.n30 13.563
R227 a_14348_27710.n50 a_14348_27710.n49 12.3446
R228 a_14348_27710.n20 a_14348_27710.n18 4.90675
R229 a_14348_27710.n31 a_14348_27710.t23 4.8248
R230 a_14348_27710.n38 a_14348_27710.t44 4.5005
R231 a_14348_27710.n37 a_14348_27710.t25 4.5005
R232 a_14348_27710.n36 a_14348_27710.t31 4.5005
R233 a_14348_27710.n35 a_14348_27710.t26 4.5005
R234 a_14348_27710.n34 a_14348_27710.t32 4.5005
R235 a_14348_27710.n33 a_14348_27710.t41 4.5005
R236 a_14348_27710.n32 a_14348_27710.t22 4.5005
R237 a_14348_27710.n31 a_14348_27710.t43 4.5005
R238 a_14348_27710.n40 a_14348_27710.t14 4.5005
R239 a_14348_27710.n39 a_14348_27710.t24 4.5005
R240 a_14348_27710.n41 a_14348_27710.t36 4.5005
R241 a_14348_27710.n42 a_14348_27710.t17 4.5005
R242 a_14348_27710.n43 a_14348_27710.t29 4.5005
R243 a_14348_27710.n44 a_14348_27710.t21 4.5005
R244 a_14348_27710.n45 a_14348_27710.t30 4.5005
R245 a_14348_27710.n46 a_14348_27710.t34 4.5005
R246 a_14348_27710.n47 a_14348_27710.t45 4.5005
R247 a_14348_27710.n48 a_14348_27710.t35 4.5005
R248 a_14348_27710.n49 a_14348_27710.t49 4.5005
R249 a_14348_27710.n15 a_14348_27710.n1 4.5005
R250 a_14348_27710.n9 a_14348_27710.n0 4.5005
R251 a_14348_27710.n17 a_14348_27710.n16 4.5005
R252 a_14348_27710.n30 a_14348_27710.n29 4.5005
R253 a_14348_27710.n29 a_14348_27710.n27 1.59425
R254 a_14348_27710.n18 a_14348_27710.n17 1.28175
R255 a_14348_27710.n22 a_14348_27710.n20 1.1255
R256 a_14348_27710.n24 a_14348_27710.n22 1.1255
R257 a_14348_27710.n30 a_14348_27710.n24 1.1255
R258 a_14348_27710.n32 a_14348_27710.n31 0.3295
R259 a_14348_27710.n33 a_14348_27710.n32 0.3295
R260 a_14348_27710.n34 a_14348_27710.n33 0.3295
R261 a_14348_27710.n35 a_14348_27710.n34 0.3295
R262 a_14348_27710.n36 a_14348_27710.n35 0.3295
R263 a_14348_27710.n37 a_14348_27710.n36 0.3295
R264 a_14348_27710.n38 a_14348_27710.n37 0.3295
R265 a_14348_27710.n40 a_14348_27710.n39 0.3295
R266 a_14348_27710.n48 a_14348_27710.n47 0.3295
R267 a_14348_27710.n47 a_14348_27710.n46 0.3295
R268 a_14348_27710.n46 a_14348_27710.n45 0.3295
R269 a_14348_27710.n45 a_14348_27710.n44 0.3295
R270 a_14348_27710.n44 a_14348_27710.n43 0.3295
R271 a_14348_27710.n43 a_14348_27710.n42 0.3295
R272 a_14348_27710.n42 a_14348_27710.n41 0.3295
R273 a_14348_27710.n49 a_14348_27710.n48 0.3248
R274 a_14348_27710.n39 a_14348_27710.n38 0.306
R275 a_14348_27710.n41 a_14348_27710.n40 0.306
R276 a_14348_27710.n3 a_14348_27710.n2 0.28175
R277 a_14348_27710.n4 a_14348_27710.n3 0.28175
R278 a_14348_27710.n5 a_14348_27710.n4 0.28175
R279 a_14348_27710.n6 a_14348_27710.n5 0.28175
R280 a_14348_27710.n7 a_14348_27710.n6 0.28175
R281 a_14348_27710.n8 a_14348_27710.n7 0.28175
R282 a_14348_27710.n9 a_14348_27710.n8 0.28175
R283 a_14348_27710.n15 a_14348_27710.n14 0.28175
R284 a_14348_27710.n14 a_14348_27710.n13 0.28175
R285 a_14348_27710.n13 a_14348_27710.n12 0.28175
R286 a_14348_27710.n12 a_14348_27710.n11 0.28175
R287 a_14348_27710.n11 a_14348_27710.n10 0.28175
R288 a_14348_27710.n16 a_14348_27710.n9 0.141125
R289 a_14348_27710.n16 a_14348_27710.n15 0.141125
R290 a_14348_27710.n17 a_14348_27710.n0 0.078625
R291 a_14348_27710.n17 a_14348_27710.n1 0.078625
R292 VGND.t40 VGND.t192 2804.76
R293 VGND.t20 VGND.t126 2533.33
R294 VGND.t323 VGND.t156 2307.14
R295 VGND.t13 VGND.t168 2216.67
R296 VGND.t128 VGND.t30 2216.67
R297 VGND.t97 VGND.t36 2216.67
R298 VGND.t133 VGND.t174 2126.19
R299 VGND.t106 VGND.t34 1538.1
R300 VGND.t315 VGND.t330 1492.86
R301 VGND.t93 VGND.t46 1492.86
R302 VGND.t7 VGND.t80 1317.78
R303 VGND.t149 VGND.n22 1289.29
R304 VGND.n252 VGND.t115 1289.29
R305 VGND.t188 VGND.t300 1130.95
R306 VGND.t104 VGND.t87 1130.95
R307 VGND.t0 VGND.t68 1130.95
R308 VGND.t42 VGND.t309 1130.95
R309 VGND.t166 VGND.t158 1130.95
R310 VGND.n251 VGND.t135 927.381
R311 VGND.t102 VGND.n106 927.381
R312 VGND.n206 VGND.t44 927.381
R313 VGND.n205 VGND.t82 927.381
R314 VGND.n749 VGND.n300 831.25
R315 VGND.n339 VGND.n338 831.25
R316 VGND.n326 VGND.n325 831.25
R317 VGND.n332 VGND.n331 831.25
R318 VGND.n148 VGND.n146 831.25
R319 VGND.n154 VGND.n144 831.25
R320 VGND.n62 VGND.t134 733.134
R321 VGND.n56 VGND.t301 733.134
R322 VGND.n575 VGND.t276 708.125
R323 VGND.t276 VGND.n552 708.125
R324 VGND.n572 VGND.t279 708.125
R325 VGND.t279 VGND.n553 708.125
R326 VGND.n601 VGND.t273 708.125
R327 VGND.t273 VGND.n548 708.125
R328 VGND.t297 VGND.n549 708.125
R329 VGND.n598 VGND.t297 708.125
R330 VGND.n677 VGND.t267 708.125
R331 VGND.t267 VGND.n670 708.125
R332 VGND.n705 VGND.t291 708.125
R333 VGND.t291 VGND.n689 708.125
R334 VGND.n723 VGND.t282 708.125
R335 VGND.t282 VGND.n684 708.125
R336 VGND.t294 VGND.n671 694.444
R337 VGND.n674 VGND.t294 694.444
R338 VGND.n253 VGND.t41 663.801
R339 VGND.n21 VGND.t305 663.801
R340 VGND.n250 VGND.t157 663.801
R341 VGND.n105 VGND.t14 663.801
R342 VGND.n207 VGND.t129 663.801
R343 VGND.n204 VGND.t37 663.801
R344 VGND.n574 VGND.t275 657.76
R345 VGND.n600 VGND.t272 657.76
R346 VGND.n243 VGND.n88 654.333
R347 VGND.n237 VGND.n91 654.333
R348 VGND.n97 VGND.n96 654.333
R349 VGND.n100 VGND.n99 654.333
R350 VGND.n117 VGND.n116 654.333
R351 VGND.n125 VGND.n124 654.333
R352 VGND.n197 VGND.n135 654.333
R353 VGND.n191 VGND.n190 654.333
R354 VGND.n77 VGND.n28 654.333
R355 VGND.n70 VGND.n31 654.333
R356 VGND.n54 VGND.n37 654.333
R357 VGND.n47 VGND.n40 654.333
R358 VGND.n7 VGND.n6 654.333
R359 VGND.n11 VGND.n10 654.333
R360 VGND.n265 VGND.n15 653.115
R361 VGND.n676 VGND.t266 640.794
R362 VGND.n704 VGND.t290 640.794
R363 VGND.n722 VGND.t281 640.794
R364 VGND.n22 VGND.t304 610.715
R365 VGND.n252 VGND.t40 610.715
R366 VGND.t156 VGND.n251 610.715
R367 VGND.n106 VGND.t13 610.715
R368 VGND.n206 VGND.t128 610.715
R369 VGND.t36 VGND.n205 610.715
R370 VGND.n653 VGND.n608 587.407
R371 VGND.n654 VGND.n651 587.407
R372 VGND.n641 VGND.n640 587.407
R373 VGND.n642 VGND.n616 587.407
R374 VGND.n338 VGND.n337 585
R375 VGND.n336 VGND.n300 585
R376 VGND.n331 VGND.n330 585
R377 VGND.n329 VGND.n325 585
R378 VGND.n644 VGND.n642 585
R379 VGND.n641 VGND.n618 585
R380 VGND.n655 VGND.n654 585
R381 VGND.n653 VGND.n611 585
R382 VGND.n151 VGND.n144 585
R383 VGND.n150 VGND.n146 585
R384 VGND.t293 VGND.n675 557.783
R385 VGND.t278 VGND.n573 540.818
R386 VGND.t296 VGND.n599 540.818
R387 VGND.n160 VGND.t341 537.492
R388 VGND.n170 VGND.t339 537.491
R389 VGND.n155 VGND.t337 537.491
R390 VGND.t287 VGND.n703 523.855
R391 VGND.t263 VGND.n721 523.855
R392 VGND.t126 VGND.t149 497.62
R393 VGND.t330 VGND.t20 497.62
R394 VGND.t66 VGND.t315 497.62
R395 VGND.t192 VGND.t66 497.62
R396 VGND.t115 VGND.t106 497.62
R397 VGND.t34 VGND.t188 497.62
R398 VGND.t300 VGND.t133 497.62
R399 VGND.t174 VGND.t93 497.62
R400 VGND.t46 VGND.t323 497.62
R401 VGND.t87 VGND.t135 497.62
R402 VGND.t168 VGND.t104 497.62
R403 VGND.t68 VGND.t102 497.62
R404 VGND.t30 VGND.t0 497.62
R405 VGND.t44 VGND.t42 497.62
R406 VGND.t309 VGND.t97 497.62
R407 VGND.t158 VGND.t82 497.62
R408 VGND.t80 VGND.t166 497.62
R409 VGND.t59 VGND.n301 465.079
R410 VGND.n335 VGND.t59 465.079
R411 VGND.n327 VGND.t191 465.079
R412 VGND.t191 VGND.n324 465.079
R413 VGND.n149 VGND.t318 465.079
R414 VGND.t318 VGND.n143 465.079
R415 VGND.n385 VGND.t322 464.281
R416 VGND.t322 VGND.n384 464.281
R417 VGND.n401 VGND.t25 464.281
R418 VGND.t25 VGND.n400 464.281
R419 VGND.t329 VGND.n407 464.281
R420 VGND.n408 VGND.t329 464.281
R421 VGND.t65 VGND.n391 464.281
R422 VGND.n392 VGND.t65 464.281
R423 VGND.t121 VGND.n318 464.281
R424 VGND.n319 VGND.t121 464.281
R425 VGND.t63 VGND.n308 464.281
R426 VGND.n309 VGND.t63 464.281
R427 VGND.n440 VGND.t327 464.281
R428 VGND.t327 VGND.n439 464.281
R429 VGND.t146 VGND.n432 464.281
R430 VGND.n433 VGND.t146 464.281
R431 VGND.n452 VGND.t307 464.281
R432 VGND.t307 VGND.n451 464.281
R433 VGND.t123 VGND.n459 464.281
R434 VGND.n460 VGND.t123 464.281
R435 VGND.n163 VGND.t120 464.281
R436 VGND.n166 VGND.t120 464.281
R437 VGND.t314 VGND.n141 464.281
R438 VGND.n173 VGND.t314 464.281
R439 VGND.t303 VGND.n487 431.421
R440 VGND.n488 VGND.t303 431.421
R441 VGND.n495 VGND.t71 431.421
R442 VGND.t71 VGND.n494 431.421
R443 VGND.n508 VGND.t84 431.421
R444 VGND.t84 VGND.n507 431.421
R445 VGND.t316 VGND.n521 431.421
R446 VGND.n522 VGND.t316 431.421
R447 VGND.n529 VGND.t112 431.421
R448 VGND.t112 VGND.n528 431.421
R449 VGND.t183 VGND.n733 431.421
R450 VGND.n734 VGND.t183 431.421
R451 VGND.n679 VGND.t265 422.384
R452 VGND.n672 VGND.t292 422.384
R453 VGND.n707 VGND.t289 418.368
R454 VGND.n700 VGND.t286 418.368
R455 VGND.n725 VGND.t280 418.368
R456 VGND.n718 VGND.t262 418.368
R457 VGND.n513 VGND.t338 415.336
R458 VGND.t143 VGND.t278 407.144
R459 VGND.t3 VGND.t143 407.144
R460 VGND.t54 VGND.t3 407.144
R461 VGND.t151 VGND.t54 407.144
R462 VGND.t180 VGND.t151 407.144
R463 VGND.t176 VGND.t180 407.144
R464 VGND.t160 VGND.t176 407.144
R465 VGND.t11 VGND.t160 407.144
R466 VGND.t109 VGND.t11 407.144
R467 VGND.t74 VGND.t109 407.144
R468 VGND.t178 VGND.t74 407.144
R469 VGND.t325 VGND.t178 407.144
R470 VGND.t48 VGND.t325 407.144
R471 VGND.t164 VGND.t48 407.144
R472 VGND.t85 VGND.t164 407.144
R473 VGND.t72 VGND.t85 407.144
R474 VGND.t124 VGND.t72 407.144
R475 VGND.t78 VGND.t124 407.144
R476 VGND.t275 VGND.t78 407.144
R477 VGND.t198 VGND.t296 407.144
R478 VGND.t137 VGND.t198 407.144
R479 VGND.t91 VGND.t137 407.144
R480 VGND.t117 VGND.t91 407.144
R481 VGND.t22 VGND.t117 407.144
R482 VGND.t204 VGND.t22 407.144
R483 VGND.t206 VGND.t204 407.144
R484 VGND.t89 VGND.t206 407.144
R485 VGND.t162 VGND.t89 407.144
R486 VGND.t153 VGND.t162 407.144
R487 VGND.t28 VGND.t153 407.144
R488 VGND.t208 VGND.t28 407.144
R489 VGND.t200 VGND.t208 407.144
R490 VGND.t50 VGND.t200 407.144
R491 VGND.t76 VGND.t50 407.144
R492 VGND.t99 VGND.t76 407.144
R493 VGND.t319 VGND.t99 407.144
R494 VGND.t202 VGND.t319 407.144
R495 VGND.t272 VGND.t202 407.144
R496 VGND.n22 VGND.n21 382.8
R497 VGND.n253 VGND.n252 382.8
R498 VGND.n251 VGND.n250 382.8
R499 VGND.n106 VGND.n105 382.8
R500 VGND.n207 VGND.n206 382.8
R501 VGND.n205 VGND.n204 382.8
R502 VGND.t101 VGND.t293 373.214
R503 VGND.t155 VGND.t101 373.214
R504 VGND.t266 VGND.t155 373.214
R505 VGND.t298 VGND.t287 373.214
R506 VGND.t139 VGND.t298 373.214
R507 VGND.t147 VGND.t139 373.214
R508 VGND.t32 VGND.t147 373.214
R509 VGND.t38 VGND.t32 373.214
R510 VGND.t26 VGND.t38 373.214
R511 VGND.t141 VGND.t26 373.214
R512 VGND.t184 VGND.t141 373.214
R513 VGND.t170 VGND.t184 373.214
R514 VGND.t332 VGND.t170 373.214
R515 VGND.t290 VGND.t332 373.214
R516 VGND.t113 VGND.t263 373.214
R517 VGND.t9 VGND.t113 373.214
R518 VGND.t18 VGND.t9 373.214
R519 VGND.t172 VGND.t18 373.214
R520 VGND.t131 VGND.t172 373.214
R521 VGND.t56 VGND.t131 373.214
R522 VGND.t186 VGND.t56 373.214
R523 VGND.t196 VGND.t186 373.214
R524 VGND.t194 VGND.t196 373.214
R525 VGND.t60 VGND.t194 373.214
R526 VGND.t281 VGND.t60 373.214
R527 VGND.n577 VGND.t274 370.168
R528 VGND.n570 VGND.t277 370.168
R529 VGND.n603 VGND.t271 370.168
R530 VGND.n596 VGND.t295 370.168
R531 VGND.n667 VGND.t268 360.868
R532 VGND.n633 VGND.t283 360.868
R533 VGND.n160 VGND.t8 359.752
R534 VGND.n170 VGND.t6 359.752
R535 VGND.n155 VGND.t17 359.752
R536 VGND.n691 VGND.t288 351.793
R537 VGND.n686 VGND.t264 351.793
R538 VGND.n410 VGND.t53 321.649
R539 VGND.t2 VGND.t308 314.113
R540 VGND.t130 VGND.t190 314.113
R541 VGND.n699 VGND.n698 301.933
R542 VGND.n697 VGND.n696 301.933
R543 VGND.n695 VGND.n694 301.933
R544 VGND.n693 VGND.n692 301.933
R545 VGND.n688 VGND.n687 301.933
R546 VGND.n716 VGND.n715 301.933
R547 VGND.n714 VGND.n713 301.933
R548 VGND.n712 VGND.n711 301.933
R549 VGND.n710 VGND.n709 301.933
R550 VGND.n683 VGND.n682 301.933
R551 VGND.n569 VGND.n568 299.231
R552 VGND.n567 VGND.n566 299.231
R553 VGND.n565 VGND.n564 299.231
R554 VGND.n563 VGND.n562 299.231
R555 VGND.n561 VGND.n560 299.231
R556 VGND.n559 VGND.n558 299.231
R557 VGND.n557 VGND.n556 299.231
R558 VGND.n555 VGND.n554 299.231
R559 VGND.n551 VGND.n550 299.231
R560 VGND.n594 VGND.n593 299.231
R561 VGND.n592 VGND.n591 299.231
R562 VGND.n590 VGND.n589 299.231
R563 VGND.n588 VGND.n587 299.231
R564 VGND.n586 VGND.n585 299.231
R565 VGND.n584 VGND.n583 299.231
R566 VGND.n582 VGND.n581 299.231
R567 VGND.n580 VGND.n579 299.231
R568 VGND.n547 VGND.n546 299.231
R569 VGND.t248 VGND.t284 251.471
R570 VGND.t240 VGND.t248 251.471
R571 VGND.t260 VGND.t240 251.471
R572 VGND.t257 VGND.t260 251.471
R573 VGND.t254 VGND.t257 251.471
R574 VGND.t252 VGND.t254 251.471
R575 VGND.t250 VGND.t252 251.471
R576 VGND.t227 VGND.t250 251.471
R577 VGND.t234 VGND.t227 251.471
R578 VGND.t232 VGND.t234 251.471
R579 VGND.t221 VGND.t232 251.471
R580 VGND.t230 VGND.t221 251.471
R581 VGND.t236 VGND.t230 251.471
R582 VGND.t225 VGND.t236 251.471
R583 VGND.t223 VGND.t225 251.471
R584 VGND.t211 VGND.t223 251.471
R585 VGND.t269 VGND.t211 251.471
R586 VGND.n320 VGND.n319 243.698
R587 VGND.n439 VGND.n344 243.698
R588 VGND.n451 VGND.n346 243.698
R589 VGND.n400 VGND.n350 243.698
R590 VGND.n384 VGND.n354 243.698
R591 VGND.n407 VGND.n351 243.698
R592 VGND.n391 VGND.n355 243.698
R593 VGND.n308 VGND.n303 243.698
R594 VGND.n432 VGND.n341 243.698
R595 VGND.n459 VGND.n347 243.698
R596 VGND.n311 VGND.n310 238.367
R597 VGND.n340 VGND.n339 238.367
R598 VGND.n333 VGND.n332 238.367
R599 VGND.n434 VGND.n342 238.367
R600 VGND.n461 VGND.n348 238.367
R601 VGND.n409 VGND.n352 238.367
R602 VGND.n393 VGND.n356 238.367
R603 VGND.n386 VGND.n353 238.367
R604 VGND.n402 VGND.n349 238.367
R605 VGND.n453 VGND.n345 238.367
R606 VGND.n441 VGND.n343 238.367
R607 VGND.n326 VGND.n322 238.367
R608 VGND.n749 VGND.n748 238.367
R609 VGND.n315 VGND.n312 238.367
R610 VGND.n573 VGND.n572 238.367
R611 VGND.n573 VGND.n553 238.367
R612 VGND.n599 VGND.n598 238.367
R613 VGND.n599 VGND.n549 238.367
R614 VGND.n648 VGND.n647 238.367
R615 VGND.n634 VGND.n613 238.367
R616 VGND.n666 VGND.n609 238.367
R617 VGND.n659 VGND.n658 238.367
R618 VGND.n675 VGND.n674 238.367
R619 VGND.n675 VGND.n671 238.367
R620 VGND.n703 VGND.n702 238.367
R621 VGND.n703 VGND.n690 238.367
R622 VGND.n721 VGND.n720 238.367
R623 VGND.n721 VGND.n685 238.367
R624 VGND.n168 VGND.n167 238.367
R625 VGND.n172 VGND.n171 238.367
R626 VGND.n154 VGND.n153 238.367
R627 VGND.n148 VGND.n147 238.367
R628 VGND.n178 VGND.n177 238.367
R629 VGND.n162 VGND.n158 238.367
R630 VGND.t284 VGND.n649 237.5
R631 VGND.n660 VGND.t269 237.5
R632 VGND.n494 VGND.n360 234.355
R633 VGND.n487 VGND.n357 234.355
R634 VGND.n507 VGND.n362 234.355
R635 VGND.n528 VGND.n366 234.355
R636 VGND.n521 VGND.n363 234.355
R637 VGND.n735 VGND.n734 234.355
R638 VGND.n489 VGND.n358 230.308
R639 VGND.n523 VGND.n364 230.308
R640 VGND.n530 VGND.n365 230.308
R641 VGND.n509 VGND.n361 230.308
R642 VGND.n496 VGND.n359 230.308
R643 VGND.n730 VGND.n367 230.308
R644 VGND.t111 VGND.t108 222.178
R645 VGND.n169 VGND.t119 219.232
R646 VGND.t313 VGND.n156 219.232
R647 VGND.t311 VGND.n142 219.232
R648 VGND.n142 VGND.t317 219.232
R649 VGND.n740 VGND.n739 199.195
R650 VGND.n170 VGND.t313 185.002
R651 VGND.t311 VGND.n155 185.002
R652 VGND.n160 VGND.t119 185.002
R653 VGND.n518 VGND.n517 185
R654 VGND.n520 VGND.n519 185
R655 VGND.n527 VGND.n526 185
R656 VGND.n525 VGND.n524 185
R657 VGND.n506 VGND.n505 185
R658 VGND.n504 VGND.n503 185
R659 VGND.n484 VGND.n483 185
R660 VGND.n486 VGND.n485 185
R661 VGND.n493 VGND.n492 185
R662 VGND.n491 VGND.n490 185
R663 VGND.n388 VGND.n387 185
R664 VGND.n390 VGND.n389 185
R665 VGND.n383 VGND.n382 185
R666 VGND.n381 VGND.n380 185
R667 VGND.n404 VGND.n403 185
R668 VGND.n406 VGND.n405 185
R669 VGND.n399 VGND.n398 185
R670 VGND.n397 VGND.n396 185
R671 VGND.n456 VGND.n455 185
R672 VGND.n458 VGND.n457 185
R673 VGND.n450 VGND.n449 185
R674 VGND.n448 VGND.n447 185
R675 VGND.n429 VGND.n428 185
R676 VGND.n431 VGND.n430 185
R677 VGND.n438 VGND.n437 185
R678 VGND.n436 VGND.n435 185
R679 VGND.n330 VGND.n323 185
R680 VGND.n329 VGND.n328 185
R681 VGND.n337 VGND.n334 185
R682 VGND.n336 VGND.n302 185
R683 VGND.n305 VGND.n304 185
R684 VGND.n307 VGND.n306 185
R685 VGND.n314 VGND.n313 185
R686 VGND.n317 VGND.n316 185
R687 VGND.n369 VGND.n368 185
R688 VGND.n732 VGND.n731 185
R689 VGND.n645 VGND.n615 185
R690 VGND.n644 VGND.n643 185
R691 VGND.n637 VGND.n618 185
R692 VGND.n639 VGND.n638 185
R693 VGND.n656 VGND.n650 185
R694 VGND.n655 VGND.n612 185
R695 VGND.n662 VGND.n611 185
R696 VGND.n664 VGND.n663 185
R697 VGND.n152 VGND.n151 185
R698 VGND.n150 VGND.n145 185
R699 VGND.n174 VGND.n157 185
R700 VGND.n176 VGND.n175 185
R701 VGND.n165 VGND.n159 185
R702 VGND.n164 VGND.n161 185
R703 VGND.t70 VGND.n738 172.38
R704 VGND.t15 VGND.n737 172.38
R705 VGND.t108 VGND.n736 172.38
R706 VGND.t5 VGND.n169 158.333
R707 VGND.n156 VGND.t16 158.333
R708 VGND.n316 VGND.n313 150
R709 VGND.n306 VGND.n304 150
R710 VGND.n334 VGND.n302 150
R711 VGND.n328 VGND.n323 150
R712 VGND.n437 VGND.n436 150
R713 VGND.n430 VGND.n429 150
R714 VGND.n449 VGND.n448 150
R715 VGND.n457 VGND.n456 150
R716 VGND.n398 VGND.n397 150
R717 VGND.n405 VGND.n404 150
R718 VGND.n382 VGND.n381 150
R719 VGND.n389 VGND.n388 150
R720 VGND.n638 VGND.n637 150
R721 VGND.n643 VGND.n615 150
R722 VGND.n663 VGND.n662 150
R723 VGND.n650 VGND.n612 150
R724 VGND.n161 VGND.n159 150
R725 VGND.n176 VGND.n157 150
R726 VGND.n152 VGND.n145 150
R727 VGND.n632 VGND.n631 141.709
R728 VGND.n630 VGND.n629 141.709
R729 VGND.n628 VGND.n627 141.709
R730 VGND.n626 VGND.n625 141.709
R731 VGND.n624 VGND.n623 141.709
R732 VGND.n622 VGND.n621 141.709
R733 VGND.n620 VGND.n619 141.709
R734 VGND.n607 VGND.n606 141.709
R735 VGND.n744 VGND.n743 137.904
R736 VGND.n742 VGND.n741 137.904
R737 VGND.n739 VGND.t70 126.412
R738 VGND.n738 VGND.t15 126.412
R739 VGND.n737 VGND.t111 126.412
R740 VGND.n736 VGND.t182 126.412
R741 VGND.t96 VGND.n300 123.126
R742 VGND.n338 VGND.t96 123.126
R743 VGND.n325 VGND.t302 123.126
R744 VGND.n331 VGND.t302 123.126
R745 VGND.t270 VGND.n653 123.126
R746 VGND.n654 VGND.t270 123.126
R747 VGND.t285 VGND.n641 123.126
R748 VGND.n642 VGND.t285 123.126
R749 VGND.n146 VGND.t312 123.126
R750 VGND.t312 VGND.n144 123.126
R751 VGND.n492 VGND.n491 120.001
R752 VGND.n485 VGND.n484 120.001
R753 VGND.n505 VGND.n504 120.001
R754 VGND.n526 VGND.n525 120.001
R755 VGND.n519 VGND.n518 120.001
R756 VGND.n731 VGND.n368 120.001
R757 VGND.t119 VGND.t7 109.615
R758 VGND.t313 VGND.t5 109.615
R759 VGND.t16 VGND.t311 109.615
R760 VGND.n746 VGND.n745 107.258
R761 VGND.t62 VGND.n321 103.427
R762 VGND.n747 VGND.t95 103.427
R763 VGND.n747 VGND.t58 103.427
R764 VGND.t145 VGND.n746 103.427
R765 VGND.n745 VGND.t122 95.7666
R766 VGND.t328 VGND.t24 91.936
R767 VGND.t64 VGND.t321 91.936
R768 VGND.n155 VGND.n154 90.5056
R769 VGND.t308 VGND.t62 84.2747
R770 VGND.t95 VGND.t2 84.2747
R771 VGND.t58 VGND.t130 84.2747
R772 VGND.t190 VGND.t145 84.2747
R773 VGND.t306 VGND.t52 84.2747
R774 VGND.n88 VGND.t136 78.8005
R775 VGND.n88 VGND.t88 78.8005
R776 VGND.n91 VGND.t105 78.8005
R777 VGND.n91 VGND.t169 78.8005
R778 VGND.n96 VGND.t103 78.8005
R779 VGND.n96 VGND.t69 78.8005
R780 VGND.n99 VGND.t1 78.8005
R781 VGND.n99 VGND.t31 78.8005
R782 VGND.n116 VGND.t45 78.8005
R783 VGND.n116 VGND.t43 78.8005
R784 VGND.n124 VGND.t310 78.8005
R785 VGND.n124 VGND.t98 78.8005
R786 VGND.n135 VGND.t83 78.8005
R787 VGND.n135 VGND.t159 78.8005
R788 VGND.n190 VGND.t167 78.8005
R789 VGND.n190 VGND.t81 78.8005
R790 VGND.n28 VGND.t47 78.8005
R791 VGND.n28 VGND.t324 78.8005
R792 VGND.n31 VGND.t175 78.8005
R793 VGND.n31 VGND.t94 78.8005
R794 VGND.n37 VGND.t35 78.8005
R795 VGND.n37 VGND.t189 78.8005
R796 VGND.n40 VGND.t116 78.8005
R797 VGND.n40 VGND.t107 78.8005
R798 VGND.n6 VGND.t150 78.8005
R799 VGND.n6 VGND.t127 78.8005
R800 VGND.n10 VGND.t21 78.8005
R801 VGND.n10 VGND.t331 78.8005
R802 VGND.n15 VGND.t67 78.8005
R803 VGND.n15 VGND.t193 78.8005
R804 VGND.n172 VGND.n170 74.7688
R805 VGND.n167 VGND.n160 74.7688
R806 VGND.n737 VGND.n364 69.8479
R807 VGND.n737 VGND.n363 69.8479
R808 VGND.n737 VGND.n366 69.8479
R809 VGND.n737 VGND.n365 69.8479
R810 VGND.n738 VGND.n362 69.8479
R811 VGND.n738 VGND.n361 69.8479
R812 VGND.n739 VGND.n358 69.8479
R813 VGND.n739 VGND.n357 69.8479
R814 VGND.n739 VGND.n360 69.8479
R815 VGND.n739 VGND.n359 69.8479
R816 VGND.n736 VGND.n735 69.8479
R817 VGND.n736 VGND.n367 69.8479
R818 VGND.n740 VGND.n356 65.8183
R819 VGND.n740 VGND.n355 65.8183
R820 VGND.n741 VGND.n354 65.8183
R821 VGND.n741 VGND.n353 65.8183
R822 VGND.n742 VGND.n352 65.8183
R823 VGND.n742 VGND.n351 65.8183
R824 VGND.n743 VGND.n350 65.8183
R825 VGND.n743 VGND.n349 65.8183
R826 VGND.n744 VGND.n348 65.8183
R827 VGND.n744 VGND.n347 65.8183
R828 VGND.n745 VGND.n346 65.8183
R829 VGND.n745 VGND.n345 65.8183
R830 VGND.n746 VGND.n342 65.8183
R831 VGND.n746 VGND.n341 65.8183
R832 VGND.n746 VGND.n344 65.8183
R833 VGND.n746 VGND.n343 65.8183
R834 VGND.n747 VGND.n333 65.8183
R835 VGND.n747 VGND.n322 65.8183
R836 VGND.n747 VGND.n340 65.8183
R837 VGND.n748 VGND.n747 65.8183
R838 VGND.n321 VGND.n311 65.8183
R839 VGND.n321 VGND.n303 65.8183
R840 VGND.n321 VGND.n320 65.8183
R841 VGND.n321 VGND.n312 65.8183
R842 VGND.n649 VGND.n648 65.8183
R843 VGND.n649 VGND.n614 65.8183
R844 VGND.n649 VGND.n613 65.8183
R845 VGND.n660 VGND.n659 65.8183
R846 VGND.n661 VGND.n660 65.8183
R847 VGND.n660 VGND.n609 65.8183
R848 VGND.n153 VGND.n142 65.8183
R849 VGND.n147 VGND.n142 65.8183
R850 VGND.n171 VGND.n156 65.8183
R851 VGND.n177 VGND.n156 65.8183
R852 VGND.n169 VGND.n168 65.8183
R853 VGND.n169 VGND.n158 65.8183
R854 VGND.n315 VGND.n292 64.4576
R855 VGND.n310 VGND.n292 64.4576
R856 VGND.n442 VGND.n441 64.4576
R857 VGND.n442 VGND.n434 64.4576
R858 VGND.n454 VGND.n453 64.4576
R859 VGND.n462 VGND.n461 64.4576
R860 VGND.n497 VGND.n496 63.6449
R861 VGND.n497 VGND.n489 63.6449
R862 VGND.n510 VGND.n509 63.6449
R863 VGND.n531 VGND.n530 63.6449
R864 VGND.n531 VGND.n523 63.6449
R865 VGND.n730 VGND.n729 63.6449
R866 VGND.n751 VGND.n298 60.8005
R867 VGND.n751 VGND.n750 60.8005
R868 VGND.n299 VGND.n298 60.8005
R869 VGND.n750 VGND.n299 60.8005
R870 VGND.n21 VGND.n2 60.8005
R871 VGND.n254 VGND.n253 60.8005
R872 VGND.n250 VGND.n249 60.8005
R873 VGND.n105 VGND.n94 60.8005
R874 VGND.n208 VGND.n207 60.8005
R875 VGND.n204 VGND.n203 60.8005
R876 VGND.n542 VGND.t335 58.8
R877 VGND.n541 VGND.t336 58.8
R878 VGND.n476 VGND.n386 58.0576
R879 VGND.n469 VGND.n402 58.0576
R880 VGND.n468 VGND.n409 58.0576
R881 VGND.n475 VGND.n393 58.0576
R882 VGND.n316 VGND.n312 53.3664
R883 VGND.n306 VGND.n303 53.3664
R884 VGND.n748 VGND.n302 53.3664
R885 VGND.n328 VGND.n322 53.3664
R886 VGND.n436 VGND.n343 53.3664
R887 VGND.n430 VGND.n341 53.3664
R888 VGND.n448 VGND.n345 53.3664
R889 VGND.n457 VGND.n347 53.3664
R890 VGND.n397 VGND.n349 53.3664
R891 VGND.n405 VGND.n351 53.3664
R892 VGND.n381 VGND.n353 53.3664
R893 VGND.n389 VGND.n355 53.3664
R894 VGND.n388 VGND.n356 53.3664
R895 VGND.n382 VGND.n354 53.3664
R896 VGND.n404 VGND.n352 53.3664
R897 VGND.n398 VGND.n350 53.3664
R898 VGND.n456 VGND.n348 53.3664
R899 VGND.n449 VGND.n346 53.3664
R900 VGND.n429 VGND.n342 53.3664
R901 VGND.n437 VGND.n344 53.3664
R902 VGND.n333 VGND.n323 53.3664
R903 VGND.n340 VGND.n334 53.3664
R904 VGND.n311 VGND.n304 53.3664
R905 VGND.n320 VGND.n313 53.3664
R906 VGND.n638 VGND.n613 53.3664
R907 VGND.n643 VGND.n614 53.3664
R908 VGND.n648 VGND.n615 53.3664
R909 VGND.n637 VGND.n614 53.3664
R910 VGND.n662 VGND.n661 53.3664
R911 VGND.n659 VGND.n650 53.3664
R912 VGND.n661 VGND.n612 53.3664
R913 VGND.n663 VGND.n609 53.3664
R914 VGND.n161 VGND.n158 53.3664
R915 VGND.n177 VGND.n176 53.3664
R916 VGND.n147 VGND.n145 53.3664
R917 VGND.n153 VGND.n152 53.3664
R918 VGND.n171 VGND.n157 53.3664
R919 VGND.n168 VGND.n159 53.3664
R920 VGND.n541 VGND.t334 49.164
R921 VGND.n543 VGND.t340 48.5159
R922 VGND.n491 VGND.n359 45.3071
R923 VGND.n485 VGND.n357 45.3071
R924 VGND.n504 VGND.n361 45.3071
R925 VGND.n525 VGND.n365 45.3071
R926 VGND.n519 VGND.n363 45.3071
R927 VGND.n518 VGND.n364 45.3071
R928 VGND.n526 VGND.n366 45.3071
R929 VGND.n505 VGND.n362 45.3071
R930 VGND.n484 VGND.n358 45.3071
R931 VGND.n492 VGND.n360 45.3071
R932 VGND.n735 VGND.n368 45.3071
R933 VGND.n731 VGND.n367 45.3071
R934 VGND.n568 VGND.t144 39.4005
R935 VGND.n568 VGND.t4 39.4005
R936 VGND.n566 VGND.t55 39.4005
R937 VGND.n566 VGND.t152 39.4005
R938 VGND.n564 VGND.t181 39.4005
R939 VGND.n564 VGND.t177 39.4005
R940 VGND.n562 VGND.t161 39.4005
R941 VGND.n562 VGND.t12 39.4005
R942 VGND.n560 VGND.t110 39.4005
R943 VGND.n560 VGND.t75 39.4005
R944 VGND.n558 VGND.t179 39.4005
R945 VGND.n558 VGND.t326 39.4005
R946 VGND.n556 VGND.t49 39.4005
R947 VGND.n556 VGND.t165 39.4005
R948 VGND.n554 VGND.t86 39.4005
R949 VGND.n554 VGND.t73 39.4005
R950 VGND.n550 VGND.t125 39.4005
R951 VGND.n550 VGND.t79 39.4005
R952 VGND.n593 VGND.t199 39.4005
R953 VGND.n593 VGND.t138 39.4005
R954 VGND.n591 VGND.t92 39.4005
R955 VGND.n591 VGND.t118 39.4005
R956 VGND.n589 VGND.t23 39.4005
R957 VGND.n589 VGND.t205 39.4005
R958 VGND.n587 VGND.t207 39.4005
R959 VGND.n587 VGND.t90 39.4005
R960 VGND.n585 VGND.t163 39.4005
R961 VGND.n585 VGND.t154 39.4005
R962 VGND.n583 VGND.t29 39.4005
R963 VGND.n583 VGND.t209 39.4005
R964 VGND.n581 VGND.t201 39.4005
R965 VGND.n581 VGND.t51 39.4005
R966 VGND.n579 VGND.t77 39.4005
R967 VGND.n579 VGND.t100 39.4005
R968 VGND.n546 VGND.t320 39.4005
R969 VGND.n546 VGND.t203 39.4005
R970 VGND.n698 VGND.t299 39.4005
R971 VGND.n698 VGND.t140 39.4005
R972 VGND.n696 VGND.t148 39.4005
R973 VGND.n696 VGND.t33 39.4005
R974 VGND.n694 VGND.t39 39.4005
R975 VGND.n694 VGND.t27 39.4005
R976 VGND.n692 VGND.t142 39.4005
R977 VGND.n692 VGND.t185 39.4005
R978 VGND.n687 VGND.t171 39.4005
R979 VGND.n687 VGND.t333 39.4005
R980 VGND.n715 VGND.t114 39.4005
R981 VGND.n715 VGND.t10 39.4005
R982 VGND.n713 VGND.t19 39.4005
R983 VGND.n713 VGND.t173 39.4005
R984 VGND.n711 VGND.t132 39.4005
R985 VGND.n711 VGND.t57 39.4005
R986 VGND.n709 VGND.t187 39.4005
R987 VGND.n709 VGND.t197 39.4005
R988 VGND.n682 VGND.t195 39.4005
R989 VGND.n682 VGND.t61 39.4005
R990 VGND.n511 VGND.n374 32.0005
R991 VGND.n516 VGND.n374 32.0005
R992 VGND.n532 VGND.n372 32.0005
R993 VGND.n536 VGND.n372 32.0005
R994 VGND.n537 VGND.n536 32.0005
R995 VGND.n538 VGND.n537 32.0005
R996 VGND.n538 VGND.n370 32.0005
R997 VGND.n759 VGND.n292 32.0005
R998 VGND.n759 VGND.n758 32.0005
R999 VGND.n758 VGND.n757 32.0005
R1000 VGND.n757 VGND.n294 32.0005
R1001 VGND.n753 VGND.n294 32.0005
R1002 VGND.n753 VGND.n752 32.0005
R1003 VGND.n752 VGND.n751 32.0005
R1004 VGND.n416 VGND.n299 32.0005
R1005 VGND.n421 VGND.n416 32.0005
R1006 VGND.n422 VGND.n421 32.0005
R1007 VGND.n423 VGND.n422 32.0005
R1008 VGND.n423 VGND.n414 32.0005
R1009 VGND.n427 VGND.n414 32.0005
R1010 VGND.n442 VGND.n427 32.0005
R1011 VGND.n443 VGND.n412 32.0005
R1012 VGND.n462 VGND.n454 32.0005
R1013 VGND.n467 VGND.n466 32.0005
R1014 VGND.n470 VGND.n394 32.0005
R1015 VGND.n474 VGND.n394 32.0005
R1016 VGND.n478 VGND.n477 32.0005
R1017 VGND.n478 VGND.n378 32.0005
R1018 VGND.n482 VGND.n378 32.0005
R1019 VGND.n497 VGND.n482 32.0005
R1020 VGND.n498 VGND.n376 32.0005
R1021 VGND.n502 VGND.n376 32.0005
R1022 VGND.n245 VGND.n23 32.0005
R1023 VGND.n245 VGND.n244 32.0005
R1024 VGND.n242 VGND.n89 32.0005
R1025 VGND.n238 VGND.n89 32.0005
R1026 VGND.n236 VGND.n92 32.0005
R1027 VGND.n232 VGND.n92 32.0005
R1028 VGND.n232 VGND.n231 32.0005
R1029 VGND.n231 VGND.n230 32.0005
R1030 VGND.n226 VGND.n225 32.0005
R1031 VGND.n225 VGND.n224 32.0005
R1032 VGND.n221 VGND.n220 32.0005
R1033 VGND.n220 VGND.n219 32.0005
R1034 VGND.n215 VGND.n214 32.0005
R1035 VGND.n214 VGND.n213 32.0005
R1036 VGND.n213 VGND.n102 32.0005
R1037 VGND.n209 VGND.n102 32.0005
R1038 VGND.n115 VGND.n104 32.0005
R1039 VGND.n118 VGND.n115 32.0005
R1040 VGND.n122 VGND.n112 32.0005
R1041 VGND.n123 VGND.n122 32.0005
R1042 VGND.n129 VGND.n110 32.0005
R1043 VGND.n130 VGND.n129 32.0005
R1044 VGND.n131 VGND.n130 32.0005
R1045 VGND.n131 VGND.n107 32.0005
R1046 VGND.n199 VGND.n108 32.0005
R1047 VGND.n199 VGND.n198 32.0005
R1048 VGND.n196 VGND.n136 32.0005
R1049 VGND.n192 VGND.n136 32.0005
R1050 VGND.n186 VGND.n185 32.0005
R1051 VGND.n185 VGND.n184 32.0005
R1052 VGND.n184 VGND.n139 32.0005
R1053 VGND.n180 VGND.n139 32.0005
R1054 VGND.n78 VGND.n26 32.0005
R1055 VGND.n82 VGND.n26 32.0005
R1056 VGND.n83 VGND.n82 32.0005
R1057 VGND.n84 VGND.n83 32.0005
R1058 VGND.n84 VGND.n24 32.0005
R1059 VGND.n71 VGND.n29 32.0005
R1060 VGND.n75 VGND.n29 32.0005
R1061 VGND.n76 VGND.n75 32.0005
R1062 VGND.n64 VGND.n63 32.0005
R1063 VGND.n64 VGND.n32 32.0005
R1064 VGND.n68 VGND.n32 32.0005
R1065 VGND.n69 VGND.n68 32.0005
R1066 VGND.n61 VGND.n34 32.0005
R1067 VGND.n57 VGND.n55 32.0005
R1068 VGND.n49 VGND.n48 32.0005
R1069 VGND.n49 VGND.n38 32.0005
R1070 VGND.n53 VGND.n38 32.0005
R1071 VGND.n289 VGND.n288 32.0005
R1072 VGND.n288 VGND.n287 32.0005
R1073 VGND.n287 VGND.n4 32.0005
R1074 VGND.n283 VGND.n282 32.0005
R1075 VGND.n282 VGND.n281 32.0005
R1076 VGND.n281 VGND.n8 32.0005
R1077 VGND.n277 VGND.n8 32.0005
R1078 VGND.n277 VGND.n276 32.0005
R1079 VGND.n276 VGND.n275 32.0005
R1080 VGND.n272 VGND.n271 32.0005
R1081 VGND.n271 VGND.n270 32.0005
R1082 VGND.n270 VGND.n13 32.0005
R1083 VGND.n266 VGND.n13 32.0005
R1084 VGND.n264 VGND.n16 32.0005
R1085 VGND.n260 VGND.n16 32.0005
R1086 VGND.n260 VGND.n259 32.0005
R1087 VGND.n259 VGND.n258 32.0005
R1088 VGND.n258 VGND.n18 32.0005
R1089 VGND.n254 VGND.n18 32.0005
R1090 VGND.n42 VGND.n20 32.0005
R1091 VGND.n42 VGND.n41 32.0005
R1092 VGND.n46 VGND.n41 32.0005
R1093 VGND.n148 VGND.n140 30.2632
R1094 VGND.n510 VGND.n502 28.8005
R1095 VGND.n249 VGND.n23 28.8005
R1096 VGND.n237 VGND.n236 28.8005
R1097 VGND.n226 VGND.n94 28.8005
R1098 VGND.n215 VGND.n100 28.8005
R1099 VGND.n208 VGND.n104 28.8005
R1100 VGND.n125 VGND.n110 28.8005
R1101 VGND.n203 VGND.n108 28.8005
R1102 VGND.n55 VGND.n54 28.8005
R1103 VGND.n266 VGND.n265 28.8005
R1104 VGND.n531 VGND.n516 25.6005
R1105 VGND.n532 VGND.n531 25.6005
R1106 VGND.n475 VGND.n474 25.6005
R1107 VGND.n179 VGND.n178 24.991
R1108 VGND.n162 VGND.n137 24.991
R1109 VGND.n189 VGND.n188 24.1894
R1110 VGND.n634 VGND.n633 22.8576
R1111 VGND.n667 VGND.n666 22.8576
R1112 VGND.n511 VGND.n510 22.4005
R1113 VGND.n238 VGND.n237 22.4005
R1114 VGND.n230 VGND.n94 22.4005
R1115 VGND.n219 VGND.n100 22.4005
R1116 VGND.n209 VGND.n208 22.4005
R1117 VGND.n125 VGND.n123 22.4005
R1118 VGND.n203 VGND.n107 22.4005
R1119 VGND.n192 VGND.n191 22.4005
R1120 VGND.n186 VGND.n137 22.4005
R1121 VGND.n180 VGND.n179 22.4005
R1122 VGND.n249 VGND.n24 22.4005
R1123 VGND.n54 VGND.n53 22.4005
R1124 VGND.n265 VGND.n264 22.4005
R1125 VGND.n729 VGND.n370 19.2005
R1126 VGND.n751 VGND.n297 19.2005
R1127 VGND.n299 VGND.n297 19.2005
R1128 VGND.n443 VGND.n442 19.2005
R1129 VGND.n454 VGND.n412 19.2005
R1130 VGND.n463 VGND.n462 19.2005
R1131 VGND.n498 VGND.n497 19.2005
R1132 VGND.n254 VGND.n20 19.2005
R1133 VGND.n291 VGND.n2 17.0989
R1134 VGND.n545 VGND.t245 17.0848
R1135 VGND.n468 VGND.n467 16.0005
R1136 VGND.n243 VGND.n242 16.0005
R1137 VGND.n221 VGND.n97 16.0005
R1138 VGND.n117 VGND.n112 16.0005
R1139 VGND.n197 VGND.n196 16.0005
R1140 VGND.n71 VGND.n70 16.0005
R1141 VGND.n77 VGND.n76 16.0005
R1142 VGND.n7 VGND.n4 16.0005
R1143 VGND.n762 VGND.n291 13.3726
R1144 VGND.n631 VGND.t249 13.1338
R1145 VGND.n631 VGND.t241 13.1338
R1146 VGND.n629 VGND.t261 13.1338
R1147 VGND.n629 VGND.t258 13.1338
R1148 VGND.n627 VGND.t255 13.1338
R1149 VGND.n627 VGND.t253 13.1338
R1150 VGND.n625 VGND.t251 13.1338
R1151 VGND.n625 VGND.t228 13.1338
R1152 VGND.n623 VGND.t235 13.1338
R1153 VGND.n623 VGND.t233 13.1338
R1154 VGND.n621 VGND.t222 13.1338
R1155 VGND.n621 VGND.t231 13.1338
R1156 VGND.n619 VGND.t237 13.1338
R1157 VGND.n619 VGND.t226 13.1338
R1158 VGND.n606 VGND.t224 13.1338
R1159 VGND.n606 VGND.t212 13.1338
R1160 VGND.n466 VGND.n410 12.8005
R1161 VGND.n470 VGND.n469 12.8005
R1162 VGND.n56 VGND.n34 12.8005
R1163 VGND.n62 VGND.n61 12.8005
R1164 VGND.n272 VGND.n11 12.8005
R1165 VGND.n762 VGND.n761 11.8717
R1166 VGND.t52 VGND.n744 11.4924
R1167 VGND.n743 VGND.t328 11.4924
R1168 VGND.t24 VGND.n742 11.4924
R1169 VGND.n741 VGND.t64 11.4924
R1170 VGND.t321 VGND.n740 11.4924
R1171 VGND.n633 VGND.n632 11.0565
R1172 VGND.n668 VGND.n667 10.8682
R1173 VGND.n48 VGND.n47 9.6005
R1174 VGND.n289 VGND.n2 9.6005
R1175 VGND.n47 VGND.n46 9.6005
R1176 VGND.n576 VGND.n552 9.50883
R1177 VGND.n602 VGND.n548 9.50883
R1178 VGND.n666 VGND.n665 9.50883
R1179 VGND.n658 VGND.n657 9.50883
R1180 VGND.n636 VGND.n634 9.50883
R1181 VGND.n647 VGND.n646 9.50883
R1182 VGND.n678 VGND.n670 9.50883
R1183 VGND.n728 VGND.n727 9.34188
R1184 VGND.n576 VGND.n575 9.3005
R1185 VGND.n602 VGND.n601 9.3005
R1186 VGND.n639 VGND.n636 9.3005
R1187 VGND.n635 VGND.n618 9.3005
R1188 VGND.n644 VGND.n617 9.3005
R1189 VGND.n646 VGND.n645 9.3005
R1190 VGND.n665 VGND.n664 9.3005
R1191 VGND.n611 VGND.n610 9.3005
R1192 VGND.n655 VGND.n652 9.3005
R1193 VGND.n657 VGND.n656 9.3005
R1194 VGND.n678 VGND.n677 9.3005
R1195 VGND.n417 VGND.n297 9.3005
R1196 VGND.n540 VGND.n370 9.3005
R1197 VGND.n539 VGND.n538 9.3005
R1198 VGND.n537 VGND.n371 9.3005
R1199 VGND.n536 VGND.n535 9.3005
R1200 VGND.n534 VGND.n372 9.3005
R1201 VGND.n533 VGND.n532 9.3005
R1202 VGND.n531 VGND.n373 9.3005
R1203 VGND.n516 VGND.n515 9.3005
R1204 VGND.n514 VGND.n374 9.3005
R1205 VGND.n512 VGND.n511 9.3005
R1206 VGND.n510 VGND.n375 9.3005
R1207 VGND.n502 VGND.n501 9.3005
R1208 VGND.n500 VGND.n376 9.3005
R1209 VGND.n499 VGND.n498 9.3005
R1210 VGND.n497 VGND.n377 9.3005
R1211 VGND.n482 VGND.n481 9.3005
R1212 VGND.n480 VGND.n378 9.3005
R1213 VGND.n479 VGND.n478 9.3005
R1214 VGND.n477 VGND.n379 9.3005
R1215 VGND.n474 VGND.n473 9.3005
R1216 VGND.n472 VGND.n394 9.3005
R1217 VGND.n471 VGND.n470 9.3005
R1218 VGND.n467 VGND.n395 9.3005
R1219 VGND.n466 VGND.n465 9.3005
R1220 VGND.n464 VGND.n463 9.3005
R1221 VGND.n462 VGND.n411 9.3005
R1222 VGND.n454 VGND.n446 9.3005
R1223 VGND.n445 VGND.n412 9.3005
R1224 VGND.n444 VGND.n443 9.3005
R1225 VGND.n442 VGND.n413 9.3005
R1226 VGND.n427 VGND.n426 9.3005
R1227 VGND.n425 VGND.n414 9.3005
R1228 VGND.n424 VGND.n423 9.3005
R1229 VGND.n422 VGND.n415 9.3005
R1230 VGND.n421 VGND.n420 9.3005
R1231 VGND.n419 VGND.n416 9.3005
R1232 VGND.n418 VGND.n299 9.3005
R1233 VGND.n751 VGND.n296 9.3005
R1234 VGND.n752 VGND.n295 9.3005
R1235 VGND.n754 VGND.n753 9.3005
R1236 VGND.n755 VGND.n294 9.3005
R1237 VGND.n757 VGND.n756 9.3005
R1238 VGND.n758 VGND.n293 9.3005
R1239 VGND.n760 VGND.n759 9.3005
R1240 VGND.n181 VGND.n180 9.3005
R1241 VGND.n182 VGND.n139 9.3005
R1242 VGND.n184 VGND.n183 9.3005
R1243 VGND.n185 VGND.n138 9.3005
R1244 VGND.n187 VGND.n186 9.3005
R1245 VGND.n193 VGND.n192 9.3005
R1246 VGND.n194 VGND.n136 9.3005
R1247 VGND.n196 VGND.n195 9.3005
R1248 VGND.n198 VGND.n134 9.3005
R1249 VGND.n200 VGND.n199 9.3005
R1250 VGND.n201 VGND.n108 9.3005
R1251 VGND.n203 VGND.n202 9.3005
R1252 VGND.n133 VGND.n107 9.3005
R1253 VGND.n132 VGND.n131 9.3005
R1254 VGND.n130 VGND.n109 9.3005
R1255 VGND.n129 VGND.n128 9.3005
R1256 VGND.n127 VGND.n110 9.3005
R1257 VGND.n126 VGND.n125 9.3005
R1258 VGND.n123 VGND.n111 9.3005
R1259 VGND.n122 VGND.n121 9.3005
R1260 VGND.n120 VGND.n112 9.3005
R1261 VGND.n119 VGND.n118 9.3005
R1262 VGND.n115 VGND.n114 9.3005
R1263 VGND.n113 VGND.n104 9.3005
R1264 VGND.n208 VGND.n103 9.3005
R1265 VGND.n210 VGND.n209 9.3005
R1266 VGND.n211 VGND.n102 9.3005
R1267 VGND.n213 VGND.n212 9.3005
R1268 VGND.n214 VGND.n101 9.3005
R1269 VGND.n216 VGND.n215 9.3005
R1270 VGND.n217 VGND.n100 9.3005
R1271 VGND.n219 VGND.n218 9.3005
R1272 VGND.n220 VGND.n98 9.3005
R1273 VGND.n222 VGND.n221 9.3005
R1274 VGND.n224 VGND.n223 9.3005
R1275 VGND.n225 VGND.n95 9.3005
R1276 VGND.n227 VGND.n226 9.3005
R1277 VGND.n228 VGND.n94 9.3005
R1278 VGND.n230 VGND.n229 9.3005
R1279 VGND.n231 VGND.n93 9.3005
R1280 VGND.n233 VGND.n232 9.3005
R1281 VGND.n234 VGND.n92 9.3005
R1282 VGND.n236 VGND.n235 9.3005
R1283 VGND.n237 VGND.n90 9.3005
R1284 VGND.n239 VGND.n238 9.3005
R1285 VGND.n240 VGND.n89 9.3005
R1286 VGND.n242 VGND.n241 9.3005
R1287 VGND.n244 VGND.n87 9.3005
R1288 VGND.n246 VGND.n245 9.3005
R1289 VGND.n247 VGND.n23 9.3005
R1290 VGND.n249 VGND.n248 9.3005
R1291 VGND.n86 VGND.n24 9.3005
R1292 VGND.n85 VGND.n84 9.3005
R1293 VGND.n83 VGND.n25 9.3005
R1294 VGND.n82 VGND.n81 9.3005
R1295 VGND.n80 VGND.n26 9.3005
R1296 VGND.n79 VGND.n78 9.3005
R1297 VGND.n76 VGND.n27 9.3005
R1298 VGND.n75 VGND.n74 9.3005
R1299 VGND.n73 VGND.n29 9.3005
R1300 VGND.n72 VGND.n71 9.3005
R1301 VGND.n69 VGND.n30 9.3005
R1302 VGND.n68 VGND.n67 9.3005
R1303 VGND.n66 VGND.n32 9.3005
R1304 VGND.n65 VGND.n64 9.3005
R1305 VGND.n63 VGND.n33 9.3005
R1306 VGND.n61 VGND.n60 9.3005
R1307 VGND.n59 VGND.n34 9.3005
R1308 VGND.n58 VGND.n57 9.3005
R1309 VGND.n55 VGND.n35 9.3005
R1310 VGND.n54 VGND.n36 9.3005
R1311 VGND.n53 VGND.n52 9.3005
R1312 VGND.n51 VGND.n38 9.3005
R1313 VGND.n50 VGND.n49 9.3005
R1314 VGND.n48 VGND.n39 9.3005
R1315 VGND.n46 VGND.n45 9.3005
R1316 VGND.n44 VGND.n41 9.3005
R1317 VGND.n43 VGND.n42 9.3005
R1318 VGND.n20 VGND.n19 9.3005
R1319 VGND.n255 VGND.n254 9.3005
R1320 VGND.n256 VGND.n18 9.3005
R1321 VGND.n258 VGND.n257 9.3005
R1322 VGND.n259 VGND.n17 9.3005
R1323 VGND.n261 VGND.n260 9.3005
R1324 VGND.n262 VGND.n16 9.3005
R1325 VGND.n264 VGND.n263 9.3005
R1326 VGND.n265 VGND.n14 9.3005
R1327 VGND.n267 VGND.n266 9.3005
R1328 VGND.n268 VGND.n13 9.3005
R1329 VGND.n270 VGND.n269 9.3005
R1330 VGND.n271 VGND.n12 9.3005
R1331 VGND.n273 VGND.n272 9.3005
R1332 VGND.n275 VGND.n274 9.3005
R1333 VGND.n276 VGND.n9 9.3005
R1334 VGND.n278 VGND.n277 9.3005
R1335 VGND.n279 VGND.n8 9.3005
R1336 VGND.n281 VGND.n280 9.3005
R1337 VGND.n282 VGND.n5 9.3005
R1338 VGND.n284 VGND.n283 9.3005
R1339 VGND.n285 VGND.n4 9.3005
R1340 VGND.n287 VGND.n286 9.3005
R1341 VGND.n288 VGND.n3 9.3005
R1342 VGND.n290 VGND.n289 9.3005
R1343 VGND.n383 VGND.n380 9.14336
R1344 VGND.n399 VGND.n396 9.14336
R1345 VGND.n406 VGND.n403 9.14336
R1346 VGND.n390 VGND.n387 9.14336
R1347 VGND.n317 VGND.n314 9.14336
R1348 VGND.n307 VGND.n305 9.14336
R1349 VGND.n438 VGND.n435 9.14336
R1350 VGND.n431 VGND.n428 9.14336
R1351 VGND.n450 VGND.n447 9.14336
R1352 VGND.n458 VGND.n455 9.14336
R1353 VGND.n639 VGND.n618 9.14336
R1354 VGND.n644 VGND.n618 9.14336
R1355 VGND.n645 VGND.n644 9.14336
R1356 VGND.n664 VGND.n611 9.14336
R1357 VGND.n655 VGND.n611 9.14336
R1358 VGND.n656 VGND.n655 9.14336
R1359 VGND.n175 VGND.n174 9.14336
R1360 VGND.n165 VGND.n164 9.14336
R1361 VGND.t122 VGND.t306 7.66179
R1362 VGND.n729 VGND.n728 7.49891
R1363 VGND.n191 VGND.n189 7.37605
R1364 VGND.n493 VGND.n490 7.11161
R1365 VGND.n486 VGND.n483 7.11161
R1366 VGND.n506 VGND.n503 7.11161
R1367 VGND.n527 VGND.n524 7.11161
R1368 VGND.n520 VGND.n517 7.11161
R1369 VGND.n732 VGND.n369 7.11161
R1370 VGND.n727 VGND.n726 7.098
R1371 VGND.n188 VGND.n137 7.05969
R1372 VGND.n179 VGND.n140 7.05957
R1373 VGND.n761 VGND.n292 6.87881
R1374 VGND.n463 VGND.n410 6.4005
R1375 VGND.n63 VGND.n62 6.4005
R1376 VGND.n57 VGND.n56 6.4005
R1377 VGND.n275 VGND.n11 6.4005
R1378 VGND.n337 VGND.n336 5.81868
R1379 VGND.n330 VGND.n329 5.81868
R1380 VGND.n151 VGND.n150 5.81868
R1381 VGND.n386 VGND.n385 5.33286
R1382 VGND.n402 VGND.n401 5.33286
R1383 VGND.n409 VGND.n408 5.33286
R1384 VGND.n393 VGND.n392 5.33286
R1385 VGND.n318 VGND.n315 5.33286
R1386 VGND.n310 VGND.n309 5.33286
R1387 VGND.n441 VGND.n440 5.33286
R1388 VGND.n434 VGND.n433 5.33286
R1389 VGND.n453 VGND.n452 5.33286
R1390 VGND.n461 VGND.n460 5.33286
R1391 VGND.n640 VGND.n634 5.33286
R1392 VGND.n647 VGND.n616 5.33286
R1393 VGND.n666 VGND.n608 5.33286
R1394 VGND.n658 VGND.n651 5.33286
R1395 VGND.n167 VGND.n166 5.33286
R1396 VGND.n178 VGND.n141 5.33286
R1397 VGND.n173 VGND.n172 5.33286
R1398 VGND.n163 VGND.n162 5.33286
R1399 VGND.n700 VGND.n699 4.84425
R1400 VGND.n702 VGND.n701 4.73979
R1401 VGND.n706 VGND.n689 4.73979
R1402 VGND.n720 VGND.n719 4.73979
R1403 VGND.n724 VGND.n684 4.73979
R1404 VGND.n771 VGND.n762 4.73554
R1405 VGND.n701 VGND.n690 4.6505
R1406 VGND.n706 VGND.n705 4.6505
R1407 VGND.n719 VGND.n685 4.6505
R1408 VGND.n724 VGND.n723 4.6505
R1409 VGND.n702 VGND.n691 4.54311
R1410 VGND.n691 VGND.n690 4.54311
R1411 VGND.n720 VGND.n686 4.54311
R1412 VGND.n686 VGND.n685 4.54311
R1413 VGND.n726 VGND.n725 4.5005
R1414 VGND.n718 VGND.n717 4.5005
R1415 VGND.n708 VGND.n707 4.5005
R1416 VGND.n575 VGND.n574 4.48641
R1417 VGND.n574 VGND.n552 4.48641
R1418 VGND.n601 VGND.n600 4.48641
R1419 VGND.n600 VGND.n548 4.48641
R1420 VGND.n677 VGND.n676 4.48641
R1421 VGND.n676 VGND.n670 4.48641
R1422 VGND.n705 VGND.n704 4.48641
R1423 VGND.n704 VGND.n689 4.48641
R1424 VGND.n723 VGND.n722 4.48641
R1425 VGND.n722 VGND.n684 4.48641
R1426 VGND.n496 VGND.n495 4.0479
R1427 VGND.n489 VGND.n488 4.0479
R1428 VGND.n509 VGND.n508 4.0479
R1429 VGND.n530 VGND.n529 4.0479
R1430 VGND.n523 VGND.n522 4.0479
R1431 VGND.n733 VGND.n730 4.0479
R1432 VGND VGND.n772 4.02487
R1433 VGND.n384 VGND.n383 3.75335
R1434 VGND.n385 VGND.n380 3.75335
R1435 VGND.n400 VGND.n399 3.75335
R1436 VGND.n401 VGND.n396 3.75335
R1437 VGND.n408 VGND.n403 3.75335
R1438 VGND.n407 VGND.n406 3.75335
R1439 VGND.n392 VGND.n387 3.75335
R1440 VGND.n391 VGND.n390 3.75335
R1441 VGND.n319 VGND.n314 3.75335
R1442 VGND.n318 VGND.n317 3.75335
R1443 VGND.n309 VGND.n305 3.75335
R1444 VGND.n308 VGND.n307 3.75335
R1445 VGND.n439 VGND.n438 3.75335
R1446 VGND.n440 VGND.n435 3.75335
R1447 VGND.n433 VGND.n428 3.75335
R1448 VGND.n432 VGND.n431 3.75335
R1449 VGND.n451 VGND.n450 3.75335
R1450 VGND.n452 VGND.n447 3.75335
R1451 VGND.n460 VGND.n455 3.75335
R1452 VGND.n459 VGND.n458 3.75335
R1453 VGND.n645 VGND.n616 3.75335
R1454 VGND.n640 VGND.n639 3.75335
R1455 VGND.n656 VGND.n651 3.75335
R1456 VGND.n664 VGND.n608 3.75335
R1457 VGND.n174 VGND.n173 3.75335
R1458 VGND.n175 VGND.n141 3.75335
R1459 VGND.n166 VGND.n165 3.75335
R1460 VGND.n164 VGND.n163 3.75335
R1461 VGND.n673 VGND.n672 3.46433
R1462 VGND.n571 VGND.n570 3.41464
R1463 VGND.n597 VGND.n596 3.41464
R1464 VGND.n767 VGND.n764 3.4105
R1465 VGND.n769 VGND.n764 3.4105
R1466 VGND.n771 VGND.n764 3.4105
R1467 VGND.n770 VGND.n769 3.4105
R1468 VGND.n771 VGND.n770 3.4105
R1469 VGND.n769 VGND.n763 3.4105
R1470 VGND.n771 VGND.n763 3.4105
R1471 VGND.n772 VGND.n771 3.4105
R1472 VGND.n749 VGND.n301 3.40194
R1473 VGND.n339 VGND.n335 3.40194
R1474 VGND.n327 VGND.n326 3.40194
R1475 VGND.n332 VGND.n324 3.40194
R1476 VGND.n149 VGND.n148 3.40194
R1477 VGND.n154 VGND.n143 3.40194
R1478 VGND.n469 VGND.n468 3.2005
R1479 VGND.n476 VGND.n475 3.2005
R1480 VGND.n477 VGND.n476 3.2005
R1481 VGND.n244 VGND.n243 3.2005
R1482 VGND.n224 VGND.n97 3.2005
R1483 VGND.n118 VGND.n117 3.2005
R1484 VGND.n198 VGND.n197 3.2005
R1485 VGND.n78 VGND.n77 3.2005
R1486 VGND.n70 VGND.n69 3.2005
R1487 VGND.n283 VGND.n7 3.2005
R1488 VGND.n571 VGND.n553 3.11118
R1489 VGND.n598 VGND.n597 3.11118
R1490 VGND.n572 VGND.n571 3.04304
R1491 VGND.n597 VGND.n549 3.04304
R1492 VGND.n494 VGND.n493 3.02841
R1493 VGND.n495 VGND.n490 3.02841
R1494 VGND.n488 VGND.n483 3.02841
R1495 VGND.n487 VGND.n486 3.02841
R1496 VGND.n507 VGND.n506 3.02841
R1497 VGND.n508 VGND.n503 3.02841
R1498 VGND.n528 VGND.n527 3.02841
R1499 VGND.n529 VGND.n524 3.02841
R1500 VGND.n522 VGND.n517 3.02841
R1501 VGND.n521 VGND.n520 3.02841
R1502 VGND.n734 VGND.n369 3.02841
R1503 VGND.n733 VGND.n732 3.02841
R1504 VGND.n674 VGND.n673 2.96855
R1505 VGND.n673 VGND.n671 2.90353
R1506 VGND.n605 VGND.n545 2.47421
R1507 VGND.n337 VGND.n335 2.39444
R1508 VGND.n336 VGND.n301 2.39444
R1509 VGND.n330 VGND.n324 2.39444
R1510 VGND.n329 VGND.n327 2.39444
R1511 VGND.n151 VGND.n143 2.39444
R1512 VGND.n150 VGND.n149 2.39444
R1513 VGND.n681 VGND.n680 2.36621
R1514 VGND.n605 VGND.n604 2.35058
R1515 VGND.n750 VGND.n749 2.32777
R1516 VGND.n332 VGND.n298 2.32777
R1517 VGND.n680 VGND.n679 2.00667
R1518 VGND.n672 VGND.n669 1.94319
R1519 VGND.n570 VGND.n569 1.90331
R1520 VGND.n604 VGND.n603 1.82095
R1521 VGND.n578 VGND.n577 1.77831
R1522 VGND.n596 VGND.n595 1.77831
R1523 VGND.n766 VGND.n765 1.70307
R1524 VGND.n768 VGND.n767 1.70307
R1525 VGND.n772 VGND.n1 1.70307
R1526 VGND.n765 VGND.n0 1.70307
R1527 VGND.n545 VGND.n543 1.05389
R1528 VGND.n717 VGND.n708 0.90675
R1529 VGND.n542 VGND.n541 0.75233
R1530 VGND.n681 VGND.n605 0.682678
R1531 VGND.n543 VGND.n542 0.648391
R1532 VGND.n699 VGND.n697 0.34425
R1533 VGND.n697 VGND.n695 0.34425
R1534 VGND.n695 VGND.n693 0.34425
R1535 VGND.n693 VGND.n688 0.34425
R1536 VGND.n708 VGND.n688 0.34425
R1537 VGND.n717 VGND.n716 0.34425
R1538 VGND.n716 VGND.n714 0.34425
R1539 VGND.n714 VGND.n712 0.34425
R1540 VGND.n712 VGND.n710 0.34425
R1541 VGND.n710 VGND.n683 0.34425
R1542 VGND.n726 VGND.n683 0.34425
R1543 VGND.n595 VGND.n578 0.333833
R1544 VGND.n669 VGND.n668 0.328625
R1545 VGND.n577 VGND.n576 0.2505
R1546 VGND.n603 VGND.n602 0.2505
R1547 VGND.n679 VGND.n678 0.2505
R1548 VGND.n727 VGND.n681 0.245239
R1549 VGND.n680 VGND.n669 0.229667
R1550 VGND.n665 VGND.n610 0.208833
R1551 VGND.n652 VGND.n610 0.208833
R1552 VGND.n657 VGND.n652 0.208833
R1553 VGND.n636 VGND.n635 0.208833
R1554 VGND.n635 VGND.n617 0.208833
R1555 VGND.n646 VGND.n617 0.208833
R1556 VGND.n761 VGND.n760 0.206321
R1557 VGND.n181 VGND.n140 0.203053
R1558 VGND.n188 VGND.n187 0.202927
R1559 VGND.n193 VGND.n189 0.196005
R1560 VGND.n728 VGND.n540 0.193961
R1561 VGND.n291 VGND.n290 0.193958
R1562 VGND.n632 VGND.n630 0.188
R1563 VGND.n630 VGND.n628 0.188
R1564 VGND.n628 VGND.n626 0.188
R1565 VGND.n626 VGND.n624 0.188
R1566 VGND.n624 VGND.n622 0.188
R1567 VGND.n622 VGND.n620 0.188
R1568 VGND.n620 VGND.n607 0.188
R1569 VGND.n668 VGND.n607 0.188
R1570 VGND.n707 VGND.n706 0.182048
R1571 VGND.n725 VGND.n724 0.182048
R1572 VGND.n701 VGND.n700 0.182048
R1573 VGND.n719 VGND.n718 0.182048
R1574 VGND.t217 VGND.t210 0.1603
R1575 VGND.t213 VGND.t217 0.1603
R1576 VGND.t218 VGND.t213 0.1603
R1577 VGND.t219 VGND.t218 0.1603
R1578 VGND.t247 VGND.t219 0.1603
R1579 VGND.t220 VGND.t247 0.1603
R1580 VGND.t256 VGND.t220 0.1603
R1581 VGND.t216 VGND.t256 0.1603
R1582 VGND.t243 VGND.t214 0.1603
R1583 VGND.t239 VGND.t243 0.1603
R1584 VGND.t242 VGND.t239 0.1603
R1585 VGND.t238 VGND.t242 0.1603
R1586 VGND.t229 VGND.t238 0.1603
R1587 VGND.t246 VGND.t229 0.1603
R1588 VGND.t215 VGND.t246 0.1603
R1589 VGND.t245 VGND.t215 0.1603
R1590 VGND.t244 VGND.n544 0.159278
R1591 VGND.n760 VGND.n293 0.15675
R1592 VGND.n756 VGND.n293 0.15675
R1593 VGND.n756 VGND.n755 0.15675
R1594 VGND.n755 VGND.n754 0.15675
R1595 VGND.n754 VGND.n295 0.15675
R1596 VGND.n296 VGND.n295 0.15675
R1597 VGND.n417 VGND.n296 0.15675
R1598 VGND.n418 VGND.n417 0.15675
R1599 VGND.n419 VGND.n418 0.15675
R1600 VGND.n420 VGND.n419 0.15675
R1601 VGND.n420 VGND.n415 0.15675
R1602 VGND.n424 VGND.n415 0.15675
R1603 VGND.n425 VGND.n424 0.15675
R1604 VGND.n426 VGND.n425 0.15675
R1605 VGND.n426 VGND.n413 0.15675
R1606 VGND.n444 VGND.n413 0.15675
R1607 VGND.n445 VGND.n444 0.15675
R1608 VGND.n446 VGND.n445 0.15675
R1609 VGND.n446 VGND.n411 0.15675
R1610 VGND.n464 VGND.n411 0.15675
R1611 VGND.n465 VGND.n464 0.15675
R1612 VGND.n465 VGND.n395 0.15675
R1613 VGND.n471 VGND.n395 0.15675
R1614 VGND.n472 VGND.n471 0.15675
R1615 VGND.n473 VGND.n472 0.15675
R1616 VGND.n473 VGND.n379 0.15675
R1617 VGND.n479 VGND.n379 0.15675
R1618 VGND.n480 VGND.n479 0.15675
R1619 VGND.n481 VGND.n480 0.15675
R1620 VGND.n481 VGND.n377 0.15675
R1621 VGND.n499 VGND.n377 0.15675
R1622 VGND.n500 VGND.n499 0.15675
R1623 VGND.n501 VGND.n500 0.15675
R1624 VGND.n501 VGND.n375 0.15675
R1625 VGND.n512 VGND.n375 0.15675
R1626 VGND.n515 VGND.n514 0.15675
R1627 VGND.n515 VGND.n373 0.15675
R1628 VGND.n533 VGND.n373 0.15675
R1629 VGND.n534 VGND.n533 0.15675
R1630 VGND.n535 VGND.n534 0.15675
R1631 VGND.n535 VGND.n371 0.15675
R1632 VGND.n539 VGND.n371 0.15675
R1633 VGND.n540 VGND.n539 0.15675
R1634 VGND.n187 VGND.n138 0.15675
R1635 VGND.n183 VGND.n138 0.15675
R1636 VGND.n183 VGND.n182 0.15675
R1637 VGND.n182 VGND.n181 0.15675
R1638 VGND.n290 VGND.n3 0.15675
R1639 VGND.n286 VGND.n3 0.15675
R1640 VGND.n286 VGND.n285 0.15675
R1641 VGND.n285 VGND.n284 0.15675
R1642 VGND.n284 VGND.n5 0.15675
R1643 VGND.n280 VGND.n5 0.15675
R1644 VGND.n280 VGND.n279 0.15675
R1645 VGND.n279 VGND.n278 0.15675
R1646 VGND.n278 VGND.n9 0.15675
R1647 VGND.n274 VGND.n9 0.15675
R1648 VGND.n274 VGND.n273 0.15675
R1649 VGND.n273 VGND.n12 0.15675
R1650 VGND.n269 VGND.n12 0.15675
R1651 VGND.n269 VGND.n268 0.15675
R1652 VGND.n268 VGND.n267 0.15675
R1653 VGND.n267 VGND.n14 0.15675
R1654 VGND.n263 VGND.n14 0.15675
R1655 VGND.n263 VGND.n262 0.15675
R1656 VGND.n262 VGND.n261 0.15675
R1657 VGND.n261 VGND.n17 0.15675
R1658 VGND.n257 VGND.n17 0.15675
R1659 VGND.n257 VGND.n256 0.15675
R1660 VGND.n256 VGND.n255 0.15675
R1661 VGND.n255 VGND.n19 0.15675
R1662 VGND.n43 VGND.n19 0.15675
R1663 VGND.n44 VGND.n43 0.15675
R1664 VGND.n45 VGND.n44 0.15675
R1665 VGND.n45 VGND.n39 0.15675
R1666 VGND.n50 VGND.n39 0.15675
R1667 VGND.n51 VGND.n50 0.15675
R1668 VGND.n52 VGND.n51 0.15675
R1669 VGND.n52 VGND.n36 0.15675
R1670 VGND.n36 VGND.n35 0.15675
R1671 VGND.n58 VGND.n35 0.15675
R1672 VGND.n59 VGND.n58 0.15675
R1673 VGND.n60 VGND.n59 0.15675
R1674 VGND.n60 VGND.n33 0.15675
R1675 VGND.n65 VGND.n33 0.15675
R1676 VGND.n66 VGND.n65 0.15675
R1677 VGND.n67 VGND.n66 0.15675
R1678 VGND.n67 VGND.n30 0.15675
R1679 VGND.n72 VGND.n30 0.15675
R1680 VGND.n73 VGND.n72 0.15675
R1681 VGND.n74 VGND.n73 0.15675
R1682 VGND.n74 VGND.n27 0.15675
R1683 VGND.n79 VGND.n27 0.15675
R1684 VGND.n80 VGND.n79 0.15675
R1685 VGND.n81 VGND.n80 0.15675
R1686 VGND.n81 VGND.n25 0.15675
R1687 VGND.n85 VGND.n25 0.15675
R1688 VGND.n86 VGND.n85 0.15675
R1689 VGND.n248 VGND.n86 0.15675
R1690 VGND.n248 VGND.n247 0.15675
R1691 VGND.n247 VGND.n246 0.15675
R1692 VGND.n246 VGND.n87 0.15675
R1693 VGND.n241 VGND.n87 0.15675
R1694 VGND.n241 VGND.n240 0.15675
R1695 VGND.n240 VGND.n239 0.15675
R1696 VGND.n239 VGND.n90 0.15675
R1697 VGND.n235 VGND.n90 0.15675
R1698 VGND.n235 VGND.n234 0.15675
R1699 VGND.n234 VGND.n233 0.15675
R1700 VGND.n233 VGND.n93 0.15675
R1701 VGND.n229 VGND.n93 0.15675
R1702 VGND.n229 VGND.n228 0.15675
R1703 VGND.n228 VGND.n227 0.15675
R1704 VGND.n227 VGND.n95 0.15675
R1705 VGND.n223 VGND.n95 0.15675
R1706 VGND.n223 VGND.n222 0.15675
R1707 VGND.n222 VGND.n98 0.15675
R1708 VGND.n218 VGND.n98 0.15675
R1709 VGND.n218 VGND.n217 0.15675
R1710 VGND.n217 VGND.n216 0.15675
R1711 VGND.n216 VGND.n101 0.15675
R1712 VGND.n212 VGND.n101 0.15675
R1713 VGND.n212 VGND.n211 0.15675
R1714 VGND.n211 VGND.n210 0.15675
R1715 VGND.n210 VGND.n103 0.15675
R1716 VGND.n113 VGND.n103 0.15675
R1717 VGND.n114 VGND.n113 0.15675
R1718 VGND.n119 VGND.n114 0.15675
R1719 VGND.n120 VGND.n119 0.15675
R1720 VGND.n121 VGND.n120 0.15675
R1721 VGND.n121 VGND.n111 0.15675
R1722 VGND.n126 VGND.n111 0.15675
R1723 VGND.n127 VGND.n126 0.15675
R1724 VGND.n128 VGND.n127 0.15675
R1725 VGND.n128 VGND.n109 0.15675
R1726 VGND.n132 VGND.n109 0.15675
R1727 VGND.n133 VGND.n132 0.15675
R1728 VGND.n202 VGND.n133 0.15675
R1729 VGND.n202 VGND.n201 0.15675
R1730 VGND.n201 VGND.n200 0.15675
R1731 VGND.n200 VGND.n134 0.15675
R1732 VGND.n195 VGND.n134 0.15675
R1733 VGND.n195 VGND.n194 0.15675
R1734 VGND.n194 VGND.n193 0.15675
R1735 VGND.t214 VGND.t244 0.137822
R1736 VGND.n544 VGND.t216 0.1368
R1737 VGND.n569 VGND.n567 0.1255
R1738 VGND.n567 VGND.n565 0.1255
R1739 VGND.n565 VGND.n563 0.1255
R1740 VGND.n563 VGND.n561 0.1255
R1741 VGND.n561 VGND.n559 0.1255
R1742 VGND.n559 VGND.n557 0.1255
R1743 VGND.n557 VGND.n555 0.1255
R1744 VGND.n555 VGND.n551 0.1255
R1745 VGND.n578 VGND.n551 0.1255
R1746 VGND.n595 VGND.n594 0.1255
R1747 VGND.n594 VGND.n592 0.1255
R1748 VGND.n592 VGND.n590 0.1255
R1749 VGND.n590 VGND.n588 0.1255
R1750 VGND.n588 VGND.n586 0.1255
R1751 VGND.n586 VGND.n584 0.1255
R1752 VGND.n584 VGND.n582 0.1255
R1753 VGND.n582 VGND.n580 0.1255
R1754 VGND.n580 VGND.n547 0.1255
R1755 VGND.n604 VGND.n547 0.1255
R1756 VGND.n513 VGND.n512 0.078625
R1757 VGND.n514 VGND.n513 0.078625
R1758 VGND.n771 VGND.n765 0.01225
R1759 VGND.n769 VGND.n765 0.01225
R1760 VGND.n767 VGND.n1 0.0068649
R1761 VGND.n770 VGND.n766 0.0068649
R1762 VGND.n768 VGND.n763 0.0068649
R1763 VGND.n772 VGND.n0 0.0068649
R1764 VGND.n766 VGND.n764 0.0068649
R1765 VGND.n770 VGND.n768 0.0068649
R1766 VGND.n763 VGND.n0 0.0068649
R1767 VGND.n769 VGND.n1 0.0068649
R1768 VGND.n544 VGND.t259 0.00152174
R1769 a_19190_31610.n15 a_19190_31610.t20 310.488
R1770 a_19190_31610.n1 a_19190_31610.t21 310.488
R1771 a_19190_31610.n6 a_19190_31610.t17 310.488
R1772 a_19190_31610.n4 a_19190_31610.n0 297.433
R1773 a_19190_31610.n9 a_19190_31610.n5 297.433
R1774 a_19190_31610.n19 a_19190_31610.n18 297.433
R1775 a_19190_31610.n13 a_19190_31610.t1 248.133
R1776 a_19190_31610.n13 a_19190_31610.n12 199.383
R1777 a_19190_31610.n14 a_19190_31610.n11 194.883
R1778 a_19190_31610.n17 a_19190_31610.t12 184.097
R1779 a_19190_31610.n3 a_19190_31610.t8 184.097
R1780 a_19190_31610.n8 a_19190_31610.t4 184.097
R1781 a_19190_31610.n16 a_19190_31610.n15 167.094
R1782 a_19190_31610.n2 a_19190_31610.n1 167.094
R1783 a_19190_31610.n7 a_19190_31610.n6 167.094
R1784 a_19190_31610.n18 a_19190_31610.n17 161.3
R1785 a_19190_31610.n4 a_19190_31610.n3 161.3
R1786 a_19190_31610.n9 a_19190_31610.n8 161.3
R1787 a_19190_31610.n16 a_19190_31610.t14 120.501
R1788 a_19190_31610.n15 a_19190_31610.t19 120.501
R1789 a_19190_31610.n2 a_19190_31610.t10 120.501
R1790 a_19190_31610.n1 a_19190_31610.t22 120.501
R1791 a_19190_31610.n7 a_19190_31610.t6 120.501
R1792 a_19190_31610.n6 a_19190_31610.t18 120.501
R1793 a_19190_31610.n12 a_19190_31610.t3 48.0005
R1794 a_19190_31610.n12 a_19190_31610.t0 48.0005
R1795 a_19190_31610.n11 a_19190_31610.t2 48.0005
R1796 a_19190_31610.n11 a_19190_31610.t16 48.0005
R1797 a_19190_31610.n17 a_19190_31610.n16 40.7027
R1798 a_19190_31610.n3 a_19190_31610.n2 40.7027
R1799 a_19190_31610.n8 a_19190_31610.n7 40.7027
R1800 a_19190_31610.n0 a_19190_31610.t9 39.4005
R1801 a_19190_31610.n0 a_19190_31610.t11 39.4005
R1802 a_19190_31610.n5 a_19190_31610.t5 39.4005
R1803 a_19190_31610.n5 a_19190_31610.t7 39.4005
R1804 a_19190_31610.n19 a_19190_31610.t13 39.4005
R1805 a_19190_31610.t15 a_19190_31610.n19 39.4005
R1806 a_19190_31610.n10 a_19190_31610.n4 6.6255
R1807 a_19190_31610.n10 a_19190_31610.n9 6.6255
R1808 a_19190_31610.n14 a_19190_31610.n13 5.2505
R1809 a_19190_31610.n18 a_19190_31610.n10 4.5005
R1810 a_19190_31610.n18 a_19190_31610.n14 0.78175
R1811 a_19190_31850.n9 a_19190_31850.t25 362.342
R1812 a_19190_31850.n23 a_19190_31850.t32 355.094
R1813 a_19190_31850.n11 a_19190_31850.n10 302.183
R1814 a_19190_31850.n20 a_19190_31850.n19 302.183
R1815 a_19190_31850.n24 a_19190_31850.n23 302.183
R1816 a_19190_31850.n16 a_19190_31850.t3 242.968
R1817 a_19190_31850.n15 a_19190_31850.n13 200.477
R1818 a_19190_31850.n15 a_19190_31850.n14 199.727
R1819 a_19190_31850.n12 a_19190_31850.t19 194.809
R1820 a_19190_31850.n12 a_19190_31850.t17 194.809
R1821 a_19190_31850.n21 a_19190_31850.t12 194.809
R1822 a_19190_31850.n21 a_19190_31850.t11 194.809
R1823 a_19190_31850.n22 a_19190_31850.n21 166.03
R1824 a_19190_31850.n17 a_19190_31850.n12 161.53
R1825 a_19190_31850.n14 a_19190_31850.t0 48.0005
R1826 a_19190_31850.n14 a_19190_31850.t1 48.0005
R1827 a_19190_31850.n13 a_19190_31850.t10 48.0005
R1828 a_19190_31850.n13 a_19190_31850.t2 48.0005
R1829 a_19190_31850.n9 a_19190_31850.n8 40.0791
R1830 a_19190_31850.n10 a_19190_31850.t4 39.4005
R1831 a_19190_31850.n10 a_19190_31850.t5 39.4005
R1832 a_19190_31850.n19 a_19190_31850.t7 39.4005
R1833 a_19190_31850.n19 a_19190_31850.t6 39.4005
R1834 a_19190_31850.n24 a_19190_31850.t8 39.4005
R1835 a_19190_31850.t9 a_19190_31850.n24 39.4005
R1836 a_19190_31850.n16 a_19190_31850.n15 5.2505
R1837 a_19190_31850.n0 a_19190_31850.t23 4.8248
R1838 a_19190_31850.n3 a_19190_31850.t18 4.5005
R1839 a_19190_31850.n3 a_19190_31850.t27 4.5005
R1840 a_19190_31850.n2 a_19190_31850.t34 4.5005
R1841 a_19190_31850.n2 a_19190_31850.t28 4.5005
R1842 a_19190_31850.n1 a_19190_31850.t36 4.5005
R1843 a_19190_31850.n1 a_19190_31850.t15 4.5005
R1844 a_19190_31850.n0 a_19190_31850.t21 4.5005
R1845 a_19190_31850.n0 a_19190_31850.t16 4.5005
R1846 a_19190_31850.n7 a_19190_31850.t31 4.5005
R1847 a_19190_31850.n3 a_19190_31850.t24 4.5005
R1848 a_19190_31850.n7 a_19190_31850.t26 4.5005
R1849 a_19190_31850.n6 a_19190_31850.t33 4.5005
R1850 a_19190_31850.n6 a_19190_31850.t13 4.5005
R1851 a_19190_31850.n4 a_19190_31850.t35 4.5005
R1852 a_19190_31850.n4 a_19190_31850.t14 4.5005
R1853 a_19190_31850.n5 a_19190_31850.t20 4.5005
R1854 a_19190_31850.n5 a_19190_31850.t29 4.5005
R1855 a_19190_31850.n8 a_19190_31850.t22 4.5005
R1856 a_19190_31850.n8 a_19190_31850.t30 4.5005
R1857 a_19190_31850.n18 a_19190_31850.n17 4.5005
R1858 a_19190_31850.n11 a_19190_31850.n9 2.93757
R1859 a_19190_31850.n1 a_19190_31850.n0 0.9875
R1860 a_19190_31850.n8 a_19190_31850.n5 0.9828
R1861 a_19190_31850.n20 a_19190_31850.n18 0.7505
R1862 a_19190_31850.n23 a_19190_31850.n22 0.7505
R1863 a_19190_31850.n4 a_19190_31850.n6 0.6585
R1864 a_19190_31850.n5 a_19190_31850.n4 0.6585
R1865 a_19190_31850.n3 a_19190_31850.n2 0.6585
R1866 a_19190_31850.n2 a_19190_31850.n1 0.6585
R1867 a_19190_31850.n6 a_19190_31850.n7 0.635
R1868 a_19190_31850.n7 a_19190_31850.n3 0.635
R1869 a_19190_31850.n17 a_19190_31850.n16 0.422375
R1870 a_19190_31850.n18 a_19190_31850.n11 0.3755
R1871 a_19190_31850.n22 a_19190_31850.n20 0.3755
R1872 a_26300_25010.n5 a_26300_25010.t1 758.734
R1873 a_26300_25010.n4 a_26300_25010.t0 758.734
R1874 a_26300_25010.n0 a_26300_25010.t5 538.234
R1875 a_26300_25010.n3 a_26300_25010.n2 342.757
R1876 a_26300_25010.t2 a_26300_25010.n5 260.733
R1877 a_26300_25010.n3 a_26300_25010.t7 190.123
R1878 a_26300_25010.n4 a_26300_25010.n3 180.8
R1879 a_26300_25010.n0 a_26300_25010.t6 136.567
R1880 a_26300_25010.n1 a_26300_25010.t4 136.567
R1881 a_26300_25010.n2 a_26300_25010.t3 136.567
R1882 a_26300_25010.n1 a_26300_25010.n0 128.534
R1883 a_26300_25010.n2 a_26300_25010.n1 128.534
R1884 a_26300_25010.n5 a_26300_25010.n4 57.6005
R1885 a_26300_25670.n2 a_26300_25670.t0 755.889
R1886 a_26300_25670.n1 a_26300_25670.t4 343.034
R1887 a_26300_25670.t1 a_26300_25670.n2 270.334
R1888 a_26300_25670.n1 a_26300_25670.n0 212.733
R1889 a_26300_25670.n0 a_26300_25670.t2 48.0005
R1890 a_26300_25670.n0 a_26300_25670.t3 48.0005
R1891 a_26300_25670.n2 a_26300_25670.n1 35.2005
R1892 VDPWR.n448 VDPWR.n447 1.97032e+06
R1893 VDPWR.n451 VDPWR.n450 589600
R1894 VDPWR.n449 VDPWR.n448 533500
R1895 VDPWR.n450 VDPWR.n449 478500
R1896 VDPWR.n46 VDPWR.n7 312538
R1897 VDPWR.n449 VDPWR.n369 286825
R1898 VDPWR.n2739 VDPWR.n9 263120
R1899 VDPWR.n2739 VDPWR.n8 132880
R1900 VDPWR.n291 VDPWR.n9 88572
R1901 VDPWR.n49 VDPWR.n48 65639.8
R1902 VDPWR.n48 VDPWR.n33 53957.9
R1903 VDPWR.n447 VDPWR.n369 40085.8
R1904 VDPWR.n369 VDPWR.t9 27530.6
R1905 VDPWR.n2734 VDPWR.n7 24406.2
R1906 VDPWR.n2727 VDPWR.n2726 19915.8
R1907 VDPWR.n46 VDPWR.n33 11350.7
R1908 VDPWR.n33 VDPWR.n15 9588.98
R1909 VDPWR.n47 VDPWR.n5 7758.04
R1910 VDPWR.n2728 VDPWR.n2727 6037.79
R1911 VDPWR.n471 VDPWR.n19 5433.26
R1912 VDPWR.n2727 VDPWR.n18 5222.9
R1913 VDPWR.n2740 VDPWR.n7 4738.46
R1914 VDPWR.n2732 VDPWR.n2731 4533.62
R1915 VDPWR.n2733 VDPWR.n15 4447.11
R1916 VDPWR.t235 VDPWR.n33 4106.67
R1917 VDPWR.n2731 VDPWR.n15 3693.93
R1918 VDPWR.n471 VDPWR.t127 3396.4
R1919 VDPWR.n2733 VDPWR.n2732 3257.69
R1920 VDPWR.t235 VDPWR.t291 3181.05
R1921 VDPWR.n2668 VDPWR.t112 2808.61
R1922 VDPWR.n2730 VDPWR.n2729 2551.48
R1923 VDPWR.n2729 VDPWR.n9 1998.47
R1924 VDPWR.n2726 VDPWR.n2725 1910.53
R1925 VDPWR.t303 VDPWR.n2669 1895.12
R1926 VDPWR.t83 VDPWR.t26 1751.46
R1927 VDPWR.n2742 VDPWR.n5 1452.43
R1928 VDPWR.t9 VDPWR.n19 1444.58
R1929 VDPWR.n2734 VDPWR.n2733 1337.98
R1930 VDPWR.n1800 VDPWR.n880 1214.72
R1931 VDPWR.n1807 VDPWR.n880 1214.72
R1932 VDPWR.n1807 VDPWR.n865 1214.72
R1933 VDPWR.n1820 VDPWR.n865 1214.72
R1934 VDPWR.n1820 VDPWR.n20 1214.72
R1935 VDPWR.n1827 VDPWR.n21 1214.72
R1936 VDPWR.n1827 VDPWR.n851 1214.72
R1937 VDPWR.n2449 VDPWR.n851 1214.72
R1938 VDPWR.n2449 VDPWR.n2448 1214.72
R1939 VDPWR.n2448 VDPWR.n22 1214.72
R1940 VDPWR.n1600 VDPWR.n1599 1214.72
R1941 VDPWR.n1599 VDPWR.n1598 1214.72
R1942 VDPWR.n1598 VDPWR.n1462 1214.72
R1943 VDPWR.n1592 VDPWR.n1462 1214.72
R1944 VDPWR.n1592 VDPWR.n23 1214.72
R1945 VDPWR.n1500 VDPWR.n24 1214.72
R1946 VDPWR.n1515 VDPWR.n1500 1214.72
R1947 VDPWR.n1515 VDPWR.n1494 1214.72
R1948 VDPWR.n1521 VDPWR.n1494 1214.72
R1949 VDPWR.n1521 VDPWR.n25 1214.72
R1950 VDPWR.n2260 VDPWR.n2123 1214.72
R1951 VDPWR.n2267 VDPWR.n2123 1214.72
R1952 VDPWR.n2267 VDPWR.n2044 1214.72
R1953 VDPWR.n2280 VDPWR.n2044 1214.72
R1954 VDPWR.n2280 VDPWR.n26 1214.72
R1955 VDPWR.n2039 VDPWR.n27 1214.72
R1956 VDPWR.n2289 VDPWR.n2039 1214.72
R1957 VDPWR.n2289 VDPWR.n2028 1214.72
R1958 VDPWR.n2325 VDPWR.n2028 1214.72
R1959 VDPWR.n2325 VDPWR.n28 1214.72
R1960 VDPWR.n2257 VDPWR.n2126 1214.72
R1961 VDPWR.n2130 VDPWR.n2126 1214.72
R1962 VDPWR.n2250 VDPWR.n2130 1214.72
R1963 VDPWR.n2250 VDPWR.n2249 1214.72
R1964 VDPWR.n2249 VDPWR.n29 1214.72
R1965 VDPWR.n2163 VDPWR.n30 1214.72
R1966 VDPWR.n2173 VDPWR.n2163 1214.72
R1967 VDPWR.n2173 VDPWR.n2020 1214.72
R1968 VDPWR.n2356 VDPWR.n2020 1214.72
R1969 VDPWR.n2356 VDPWR.n31 1214.72
R1970 VDPWR.n292 VDPWR.n213 1210.53
R1971 VDPWR.n368 VDPWR.n225 1210.53
R1972 VDPWR.n366 VDPWR.n237 1210.53
R1973 VDPWR.t7 VDPWR.n2658 1186
R1974 VDPWR.t7 VDPWR.n2667 1186
R1975 VDPWR.n2716 VDPWR.n2715 1186
R1976 VDPWR.n2723 VDPWR.n2722 1186
R1977 VDPWR.n170 VDPWR.n92 1182.8
R1978 VDPWR.n582 VDPWR.n581 1182.8
R1979 VDPWR.n463 VDPWR.n462 1173.78
R1980 VDPWR.n470 VDPWR.n469 1173.78
R1981 VDPWR.n457 VDPWR.n456 1173.78
R1982 VDPWR.n472 VDPWR.n471 1170
R1983 VDPWR.t112 VDPWR.t235 1115.59
R1984 VDPWR.n2740 VDPWR.n2739 1110.68
R1985 VDPWR.n2670 VDPWR.t303 979.318
R1986 VDPWR.t228 VDPWR.t184 974.047
R1987 VDPWR.t70 VDPWR.n2736 833.01
R1988 VDPWR.t20 VDPWR.n2735 833.01
R1989 VDPWR.t167 VDPWR.t203 808.649
R1990 VDPWR.n49 VDPWR.n5 806.668
R1991 VDPWR.n690 VDPWR.t315 789.313
R1992 VDPWR.t173 VDPWR.t308 784.865
R1993 VDPWR.n47 VDPWR.n46 755.076
R1994 VDPWR.n446 VDPWR.n8 745.129
R1995 VDPWR.n462 VDPWR.t318 728.524
R1996 VDPWR.n469 VDPWR.t322 728.524
R1997 VDPWR.n456 VDPWR.t319 728.524
R1998 VDPWR.n2724 VDPWR.t235 704.505
R1999 VDPWR.n2579 VDPWR.n2578 686.717
R2000 VDPWR.n2587 VDPWR.n2586 686.717
R2001 VDPWR.n2600 VDPWR.n2599 686.717
R2002 VDPWR.n2609 VDPWR.n2608 686.717
R2003 VDPWR.n2614 VDPWR.n2612 686.717
R2004 VDPWR.n452 VDPWR.n247 686.717
R2005 VDPWR.n458 VDPWR.n251 686.717
R2006 VDPWR.n465 VDPWR.n464 686.717
R2007 VDPWR.n467 VDPWR.n464 686.717
R2008 VDPWR.n460 VDPWR.n458 686.717
R2009 VDPWR.n454 VDPWR.n452 686.717
R2010 VDPWR.n2615 VDPWR.n2614 686.717
R2011 VDPWR.n296 VDPWR.n295 673.669
R2012 VDPWR.n364 VDPWR.n363 673.669
R2013 VDPWR.n2732 VDPWR.t146 671.756
R2014 VDPWR.n2560 VDPWR.n2559 669.307
R2015 VDPWR.n2538 VDPWR.n2535 669.307
R2016 VDPWR.n278 VDPWR.n277 669.307
R2017 VDPWR.n334 VDPWR.n257 669.307
R2018 VDPWR.n359 VDPWR.n258 669.307
R2019 VDPWR.n341 VDPWR.n256 669.307
R2020 VDPWR.n284 VDPWR.n283 669.307
R2021 VDPWR.n301 VDPWR.n300 669.307
R2022 VDPWR.n2623 VDPWR.n2622 654.962
R2023 VDPWR.t235 VDPWR.n21 634.356
R2024 VDPWR.t235 VDPWR.n24 634.356
R2025 VDPWR.t235 VDPWR.n27 634.356
R2026 VDPWR.t235 VDPWR.n30 634.356
R2027 VDPWR.n2671 VDPWR.t7 629.396
R2028 VDPWR.n2734 VDPWR.n14 621.375
R2029 VDPWR.t105 VDPWR.t290 616.66
R2030 VDPWR.n2738 VDPWR.n2737 598.058
R2031 VDPWR.n2657 VDPWR.n2656 589.889
R2032 VDPWR.n2741 VDPWR.n6 585.003
R2033 VDPWR.n444 VDPWR.n371 585.003
R2034 VDPWR.n94 VDPWR.n93 585.001
R2035 VDPWR.n583 VDPWR.n86 585.001
R2036 VDPWR.n585 VDPWR.n584 585.001
R2037 VDPWR.n423 VDPWR.n422 585.001
R2038 VDPWR.n421 VDPWR.n418 585.001
R2039 VDPWR.n442 VDPWR.n441 585.001
R2040 VDPWR.n443 VDPWR.n372 585.001
R2041 VDPWR.n445 VDPWR.n370 585.001
R2042 VDPWR.n691 VDPWR.n690 585.001
R2043 VDPWR.n683 VDPWR.n16 585.001
R2044 VDPWR.n676 VDPWR.n14 585.001
R2045 VDPWR.n2735 VDPWR.n13 585.001
R2046 VDPWR.n2736 VDPWR.n12 585.001
R2047 VDPWR.n2737 VDPWR.n11 585.001
R2048 VDPWR.n2738 VDPWR.n10 585.001
R2049 VDPWR.n2743 VDPWR.n2742 585.001
R2050 VDPWR.n2714 VDPWR.n2713 585.001
R2051 VDPWR.n1578 VDPWR.n1223 585
R2052 VDPWR.n1600 VDPWR.n1223 585
R2053 VDPWR.n1580 VDPWR.n1460 585
R2054 VDPWR.n1599 VDPWR.n1460 585
R2055 VDPWR.n1581 VDPWR.n1461 585
R2056 VDPWR.n1598 VDPWR.n1461 585
R2057 VDPWR.n1471 VDPWR.n1466 585
R2058 VDPWR.n1466 VDPWR.n1462 585
R2059 VDPWR.n1591 VDPWR.n1590 585
R2060 VDPWR.n1592 VDPWR.n1591 585
R2061 VDPWR.n1469 VDPWR.n1467 585
R2062 VDPWR.n1467 VDPWR.n23 585
R2063 VDPWR.n1505 VDPWR.n1504 585
R2064 VDPWR.n1504 VDPWR.n24 585
R2065 VDPWR.n1502 VDPWR.n1501 585
R2066 VDPWR.n1501 VDPWR.n1500 585
R2067 VDPWR.n1514 VDPWR.n1513 585
R2068 VDPWR.n1515 VDPWR.n1514 585
R2069 VDPWR.n1493 VDPWR.n1490 585
R2070 VDPWR.n1494 VDPWR.n1493 585
R2071 VDPWR.n1523 VDPWR.n1522 585
R2072 VDPWR.n1522 VDPWR.n1521 585
R2073 VDPWR.n1491 VDPWR.n819 585
R2074 VDPWR.n819 VDPWR.n25 585
R2075 VDPWR.n815 VDPWR.n811 585
R2076 VDPWR.n811 VDPWR.n25 585
R2077 VDPWR.n1520 VDPWR.n1519 585
R2078 VDPWR.n1521 VDPWR.n1520 585
R2079 VDPWR.n1518 VDPWR.n1495 585
R2080 VDPWR.n1495 VDPWR.n1494 585
R2081 VDPWR.n1517 VDPWR.n1516 585
R2082 VDPWR.n1516 VDPWR.n1515 585
R2083 VDPWR.n1499 VDPWR.n1496 585
R2084 VDPWR.n1500 VDPWR.n1499 585
R2085 VDPWR.n1498 VDPWR.n1497 585
R2086 VDPWR.n1498 VDPWR.n24 585
R2087 VDPWR.n1465 VDPWR.n1464 585
R2088 VDPWR.n1465 VDPWR.n23 585
R2089 VDPWR.n1594 VDPWR.n1593 585
R2090 VDPWR.n1593 VDPWR.n1592 585
R2091 VDPWR.n1595 VDPWR.n1463 585
R2092 VDPWR.n1463 VDPWR.n1462 585
R2093 VDPWR.n1597 VDPWR.n1596 585
R2094 VDPWR.n1598 VDPWR.n1597 585
R2095 VDPWR.n1459 VDPWR.n1226 585
R2096 VDPWR.n1599 VDPWR.n1459 585
R2097 VDPWR.n1602 VDPWR.n1601 585
R2098 VDPWR.n1601 VDPWR.n1600 585
R2099 VDPWR.n2328 VDPWR.n2327 585
R2100 VDPWR.n2327 VDPWR.n28 585
R2101 VDPWR.n2326 VDPWR.n2026 585
R2102 VDPWR.n2326 VDPWR.n2325 585
R2103 VDPWR.n2286 VDPWR.n2027 585
R2104 VDPWR.n2028 VDPWR.n2027 585
R2105 VDPWR.n2288 VDPWR.n2287 585
R2106 VDPWR.n2289 VDPWR.n2288 585
R2107 VDPWR.n2285 VDPWR.n2040 585
R2108 VDPWR.n2040 VDPWR.n2039 585
R2109 VDPWR.n2284 VDPWR.n2283 585
R2110 VDPWR.n2283 VDPWR.n27 585
R2111 VDPWR.n2282 VDPWR.n2041 585
R2112 VDPWR.n2282 VDPWR.n26 585
R2113 VDPWR.n2281 VDPWR.n2043 585
R2114 VDPWR.n2281 VDPWR.n2280 585
R2115 VDPWR.n2264 VDPWR.n2042 585
R2116 VDPWR.n2044 VDPWR.n2042 585
R2117 VDPWR.n2266 VDPWR.n2265 585
R2118 VDPWR.n2267 VDPWR.n2266 585
R2119 VDPWR.n2263 VDPWR.n2124 585
R2120 VDPWR.n2124 VDPWR.n2123 585
R2121 VDPWR.n2262 VDPWR.n2261 585
R2122 VDPWR.n2261 VDPWR.n2260 585
R2123 VDPWR.n2358 VDPWR.n2017 585
R2124 VDPWR.n2358 VDPWR.n31 585
R2125 VDPWR.n2357 VDPWR.n2019 585
R2126 VDPWR.n2357 VDPWR.n2356 585
R2127 VDPWR.n2170 VDPWR.n2018 585
R2128 VDPWR.n2020 VDPWR.n2018 585
R2129 VDPWR.n2172 VDPWR.n2171 585
R2130 VDPWR.n2173 VDPWR.n2172 585
R2131 VDPWR.n2169 VDPWR.n2164 585
R2132 VDPWR.n2164 VDPWR.n2163 585
R2133 VDPWR.n2168 VDPWR.n2167 585
R2134 VDPWR.n2167 VDPWR.n30 585
R2135 VDPWR.n2166 VDPWR.n2165 585
R2136 VDPWR.n2166 VDPWR.n29 585
R2137 VDPWR.n2129 VDPWR.n2128 585
R2138 VDPWR.n2249 VDPWR.n2129 585
R2139 VDPWR.n2252 VDPWR.n2251 585
R2140 VDPWR.n2251 VDPWR.n2250 585
R2141 VDPWR.n2253 VDPWR.n2127 585
R2142 VDPWR.n2130 VDPWR.n2127 585
R2143 VDPWR.n2255 VDPWR.n2254 585
R2144 VDPWR.n2255 VDPWR.n2126 585
R2145 VDPWR.n2256 VDPWR.n816 585
R2146 VDPWR.n2257 VDPWR.n2256 585
R2147 VDPWR.n2233 VDPWR.n2125 585
R2148 VDPWR.n2257 VDPWR.n2125 585
R2149 VDPWR.n2236 VDPWR.n2235 585
R2150 VDPWR.n2236 VDPWR.n2126 585
R2151 VDPWR.n2238 VDPWR.n2237 585
R2152 VDPWR.n2237 VDPWR.n2130 585
R2153 VDPWR.n2136 VDPWR.n2131 585
R2154 VDPWR.n2250 VDPWR.n2131 585
R2155 VDPWR.n2248 VDPWR.n2247 585
R2156 VDPWR.n2249 VDPWR.n2248 585
R2157 VDPWR.n2134 VDPWR.n2132 585
R2158 VDPWR.n2132 VDPWR.n29 585
R2159 VDPWR.n2161 VDPWR.n2160 585
R2160 VDPWR.n2161 VDPWR.n30 585
R2161 VDPWR.n2162 VDPWR.n2157 585
R2162 VDPWR.n2163 VDPWR.n2162 585
R2163 VDPWR.n2175 VDPWR.n2174 585
R2164 VDPWR.n2174 VDPWR.n2173 585
R2165 VDPWR.n2153 VDPWR.n2021 585
R2166 VDPWR.n2021 VDPWR.n2020 585
R2167 VDPWR.n2355 VDPWR.n2354 585
R2168 VDPWR.n2356 VDPWR.n2355 585
R2169 VDPWR.n2352 VDPWR.n2022 585
R2170 VDPWR.n2022 VDPWR.n31 585
R2171 VDPWR.n2479 VDPWR.n814 585
R2172 VDPWR.n812 VDPWR.n809 585
R2173 VDPWR.n2484 VDPWR.n808 585
R2174 VDPWR.n2485 VDPWR.n806 585
R2175 VDPWR.n2486 VDPWR.n805 585
R2176 VDPWR.n803 VDPWR.n800 585
R2177 VDPWR.n2491 VDPWR.n799 585
R2178 VDPWR.n2492 VDPWR.n797 585
R2179 VDPWR.n2493 VDPWR.n796 585
R2180 VDPWR.n794 VDPWR.n790 585
R2181 VDPWR.n793 VDPWR.n789 585
R2182 VDPWR.n2500 VDPWR.n788 585
R2183 VDPWR.n2456 VDPWR.n845 585
R2184 VDPWR.n2457 VDPWR.n843 585
R2185 VDPWR.n2458 VDPWR.n842 585
R2186 VDPWR.n840 VDPWR.n837 585
R2187 VDPWR.n2463 VDPWR.n836 585
R2188 VDPWR.n2464 VDPWR.n834 585
R2189 VDPWR.n2465 VDPWR.n833 585
R2190 VDPWR.n831 VDPWR.n828 585
R2191 VDPWR.n2470 VDPWR.n827 585
R2192 VDPWR.n2471 VDPWR.n825 585
R2193 VDPWR.n2472 VDPWR.n824 585
R2194 VDPWR.n822 VDPWR.n820 585
R2195 VDPWR.n2477 VDPWR.n817 585
R2196 VDPWR.n817 VDPWR.n36 585
R2197 VDPWR.n2480 VDPWR.n2479 585
R2198 VDPWR.n2482 VDPWR.n809 585
R2199 VDPWR.n2484 VDPWR.n2483 585
R2200 VDPWR.n2485 VDPWR.n802 585
R2201 VDPWR.n2487 VDPWR.n2486 585
R2202 VDPWR.n2489 VDPWR.n800 585
R2203 VDPWR.n2491 VDPWR.n2490 585
R2204 VDPWR.n2492 VDPWR.n791 585
R2205 VDPWR.n2494 VDPWR.n2493 585
R2206 VDPWR.n2496 VDPWR.n790 585
R2207 VDPWR.n2497 VDPWR.n789 585
R2208 VDPWR.n2500 VDPWR.n2499 585
R2209 VDPWR.n2456 VDPWR.n2455 585
R2210 VDPWR.n2457 VDPWR.n839 585
R2211 VDPWR.n2459 VDPWR.n2458 585
R2212 VDPWR.n2461 VDPWR.n837 585
R2213 VDPWR.n2463 VDPWR.n2462 585
R2214 VDPWR.n2464 VDPWR.n830 585
R2215 VDPWR.n2466 VDPWR.n2465 585
R2216 VDPWR.n2468 VDPWR.n828 585
R2217 VDPWR.n2470 VDPWR.n2469 585
R2218 VDPWR.n2471 VDPWR.n821 585
R2219 VDPWR.n2473 VDPWR.n2472 585
R2220 VDPWR.n2475 VDPWR.n820 585
R2221 VDPWR.n2477 VDPWR.n2476 585
R2222 VDPWR.n2476 VDPWR.n34 585
R2223 VDPWR.n1458 VDPWR.n1225 585
R2224 VDPWR.n1456 VDPWR.n1455 585
R2225 VDPWR.n1228 VDPWR.n1227 585
R2226 VDPWR.n1368 VDPWR.n1367 585
R2227 VDPWR.n1369 VDPWR.n1365 585
R2228 VDPWR.n1363 VDPWR.n1359 585
R2229 VDPWR.n1374 VDPWR.n1358 585
R2230 VDPWR.n1375 VDPWR.n1356 585
R2231 VDPWR.n1376 VDPWR.n1355 585
R2232 VDPWR.n1353 VDPWR.n1350 585
R2233 VDPWR.n1381 VDPWR.n1349 585
R2234 VDPWR.n1382 VDPWR.n1347 585
R2235 VDPWR.n1452 VDPWR.n1225 585
R2236 VDPWR.n1455 VDPWR.n1454 585
R2237 VDPWR.n1229 VDPWR.n1228 585
R2238 VDPWR.n1368 VDPWR.n1362 585
R2239 VDPWR.n1370 VDPWR.n1369 585
R2240 VDPWR.n1372 VDPWR.n1359 585
R2241 VDPWR.n1374 VDPWR.n1373 585
R2242 VDPWR.n1375 VDPWR.n1352 585
R2243 VDPWR.n1377 VDPWR.n1376 585
R2244 VDPWR.n1379 VDPWR.n1350 585
R2245 VDPWR.n1381 VDPWR.n1380 585
R2246 VDPWR.n1382 VDPWR.n1343 585
R2247 VDPWR.n2388 VDPWR.n2387 585
R2248 VDPWR.n2390 VDPWR.n2389 585
R2249 VDPWR.n2392 VDPWR.n2391 585
R2250 VDPWR.n2394 VDPWR.n2393 585
R2251 VDPWR.n2396 VDPWR.n2395 585
R2252 VDPWR.n2398 VDPWR.n2397 585
R2253 VDPWR.n2400 VDPWR.n2399 585
R2254 VDPWR.n2402 VDPWR.n2401 585
R2255 VDPWR.n2404 VDPWR.n2403 585
R2256 VDPWR.n2406 VDPWR.n2405 585
R2257 VDPWR.n2408 VDPWR.n2407 585
R2258 VDPWR.n2410 VDPWR.n2409 585
R2259 VDPWR.n1711 VDPWR.n1710 585
R2260 VDPWR.n1709 VDPWR.n1708 585
R2261 VDPWR.n1707 VDPWR.n1706 585
R2262 VDPWR.n1705 VDPWR.n1704 585
R2263 VDPWR.n1703 VDPWR.n1702 585
R2264 VDPWR.n1701 VDPWR.n1700 585
R2265 VDPWR.n1699 VDPWR.n1698 585
R2266 VDPWR.n1697 VDPWR.n1696 585
R2267 VDPWR.n1695 VDPWR.n1694 585
R2268 VDPWR.n1693 VDPWR.n1692 585
R2269 VDPWR.n1691 VDPWR.n1690 585
R2270 VDPWR.n1689 VDPWR.n1688 585
R2271 VDPWR.n260 VDPWR.n259 585
R2272 VDPWR.n361 VDPWR.n360 585
R2273 VDPWR.n338 VDPWR.n337 585
R2274 VDPWR.n336 VDPWR.n332 585
R2275 VDPWR.n280 VDPWR.n274 585
R2276 VDPWR.n282 VDPWR.n281 585
R2277 VDPWR.n297 VDPWR.n294 585
R2278 VDPWR.n299 VDPWR.n298 585
R2279 VDPWR.n2670 VDPWR.n2657 585
R2280 VDPWR.n2673 VDPWR.n2672 585
R2281 VDPWR.n2672 VDPWR.n2671 585
R2282 VDPWR.n2360 VDPWR.n2359 585
R2283 VDPWR.n2362 VDPWR.n2361 585
R2284 VDPWR.n2364 VDPWR.n2363 585
R2285 VDPWR.n2366 VDPWR.n2365 585
R2286 VDPWR.n2368 VDPWR.n2367 585
R2287 VDPWR.n2370 VDPWR.n2369 585
R2288 VDPWR.n2372 VDPWR.n2371 585
R2289 VDPWR.n2374 VDPWR.n2373 585
R2290 VDPWR.n2376 VDPWR.n2375 585
R2291 VDPWR.n2378 VDPWR.n2377 585
R2292 VDPWR.n2380 VDPWR.n2379 585
R2293 VDPWR.n2384 VDPWR.n2383 585
R2294 VDPWR.n2329 VDPWR.n1877 585
R2295 VDPWR.n2384 VDPWR.n1877 585
R2296 VDPWR.n2331 VDPWR.n2330 585
R2297 VDPWR.n2333 VDPWR.n2332 585
R2298 VDPWR.n2335 VDPWR.n2334 585
R2299 VDPWR.n2337 VDPWR.n2336 585
R2300 VDPWR.n2339 VDPWR.n2338 585
R2301 VDPWR.n2341 VDPWR.n2340 585
R2302 VDPWR.n2343 VDPWR.n2342 585
R2303 VDPWR.n2345 VDPWR.n2344 585
R2304 VDPWR.n2347 VDPWR.n2346 585
R2305 VDPWR.n2349 VDPWR.n2348 585
R2306 VDPWR.n2351 VDPWR.n2025 585
R2307 VDPWR.n2351 VDPWR.n2350 585
R2308 VDPWR.n2386 VDPWR.n1869 585
R2309 VDPWR.n2301 VDPWR.n1870 585
R2310 VDPWR.n2303 VDPWR.n2302 585
R2311 VDPWR.n2305 VDPWR.n2304 585
R2312 VDPWR.n2307 VDPWR.n2306 585
R2313 VDPWR.n2309 VDPWR.n2308 585
R2314 VDPWR.n2311 VDPWR.n2310 585
R2315 VDPWR.n2313 VDPWR.n2312 585
R2316 VDPWR.n2315 VDPWR.n2314 585
R2317 VDPWR.n2317 VDPWR.n2316 585
R2318 VDPWR.n2319 VDPWR.n2318 585
R2319 VDPWR.n2607 VDPWR.n2594 585
R2320 VDPWR.n2606 VDPWR.n2605 585
R2321 VDPWR.n2606 VDPWR.t0 585
R2322 VDPWR.n2601 VDPWR.n2596 585
R2323 VDPWR.n2541 VDPWR.n2536 585
R2324 VDPWR.n2543 VDPWR.n2542 585
R2325 VDPWR.n2544 VDPWR.n2543 585
R2326 VDPWR.n1978 VDPWR.n787 585
R2327 VDPWR.n1979 VDPWR.n1978 585
R2328 VDPWR.n1977 VDPWR.n786 585
R2329 VDPWR.n1980 VDPWR.n1977 585
R2330 VDPWR.n1983 VDPWR.n1982 585
R2331 VDPWR.n1982 VDPWR.n1981 585
R2332 VDPWR.n1984 VDPWR.n1905 585
R2333 VDPWR.n1905 VDPWR.n1904 585
R2334 VDPWR.n1993 VDPWR.n1992 585
R2335 VDPWR.n1994 VDPWR.n1993 585
R2336 VDPWR.n1908 VDPWR.n1903 585
R2337 VDPWR.n1995 VDPWR.n1903 585
R2338 VDPWR.n1997 VDPWR.n1902 585
R2339 VDPWR.n1997 VDPWR.n1996 585
R2340 VDPWR.n1999 VDPWR.n1998 585
R2341 VDPWR.n1998 VDPWR.n53 585
R2342 VDPWR.n1899 VDPWR.n1895 585
R2343 VDPWR.n1895 VDPWR.n1894 585
R2344 VDPWR.n2009 VDPWR.n2008 585
R2345 VDPWR.n2010 VDPWR.n2009 585
R2346 VDPWR.n1897 VDPWR.n1893 585
R2347 VDPWR.n2011 VDPWR.n1893 585
R2348 VDPWR.n2014 VDPWR.n2013 585
R2349 VDPWR.n2013 VDPWR.n2012 585
R2350 VDPWR.n2016 VDPWR.n1890 585
R2351 VDPWR.n1890 VDPWR.n52 585
R2352 VDPWR.n2561 VDPWR.n703 585
R2353 VDPWR.n2557 VDPWR.n702 585
R2354 VDPWR.n2558 VDPWR.n2557 585
R2355 VDPWR.n2585 VDPWR.n2584 585
R2356 VDPWR.n2582 VDPWR.n2574 585
R2357 VDPWR.n2574 VDPWR.t98 585
R2358 VDPWR.n2577 VDPWR.n2575 585
R2359 VDPWR.n1384 VDPWR.n1344 585
R2360 VDPWR.n1344 VDPWR.n44 585
R2361 VDPWR.n1346 VDPWR.n706 585
R2362 VDPWR.n706 VDPWR.n704 585
R2363 VDPWR.n2555 VDPWR.n2554 585
R2364 VDPWR.n2556 VDPWR.n2555 585
R2365 VDPWR.n709 VDPWR.n707 585
R2366 VDPWR.n707 VDPWR.n705 585
R2367 VDPWR.n2513 VDPWR.n2512 585
R2368 VDPWR.n2512 VDPWR.n2511 585
R2369 VDPWR.n2516 VDPWR.n2508 585
R2370 VDPWR.n2510 VDPWR.n2508 585
R2371 VDPWR.n2521 VDPWR.n2520 585
R2372 VDPWR.n2521 VDPWR.n32 585
R2373 VDPWR.n2524 VDPWR.n2523 585
R2374 VDPWR.n2523 VDPWR.n2522 585
R2375 VDPWR.n2506 VDPWR.n2505 585
R2376 VDPWR.n2505 VDPWR.n2504 585
R2377 VDPWR.n2531 VDPWR.n2530 585
R2378 VDPWR.n2532 VDPWR.n2531 585
R2379 VDPWR.n784 VDPWR.n730 585
R2380 VDPWR.n2533 VDPWR.n784 585
R2381 VDPWR.n2547 VDPWR.n2546 585
R2382 VDPWR.n2546 VDPWR.n2545 585
R2383 VDPWR.n2503 VDPWR.n2502 585
R2384 VDPWR.n2534 VDPWR.n2503 585
R2385 VDPWR.n787 VDPWR.n785 585
R2386 VDPWR.n785 VDPWR.n35 585
R2387 VDPWR.n1404 VDPWR.n1403 585
R2388 VDPWR.n1403 VDPWR.n38 585
R2389 VDPWR.n1402 VDPWR.n1238 585
R2390 VDPWR.n1402 VDPWR.n1401 585
R2391 VDPWR.n1264 VDPWR.n1237 585
R2392 VDPWR.n1400 VDPWR.n1237 585
R2393 VDPWR.n1398 VDPWR.n1397 585
R2394 VDPWR.n1399 VDPWR.n1398 585
R2395 VDPWR.n1242 VDPWR.n1240 585
R2396 VDPWR.n1240 VDPWR.n1239 585
R2397 VDPWR.n1326 VDPWR.n1325 585
R2398 VDPWR.n1325 VDPWR.n40 585
R2399 VDPWR.n1329 VDPWR.n1323 585
R2400 VDPWR.n1323 VDPWR.n1322 585
R2401 VDPWR.n1337 VDPWR.n1336 585
R2402 VDPWR.n1338 VDPWR.n1337 585
R2403 VDPWR.n1332 VDPWR.n1321 585
R2404 VDPWR.n1339 VDPWR.n1321 585
R2405 VDPWR.n1341 VDPWR.n1263 585
R2406 VDPWR.n1341 VDPWR.n1340 585
R2407 VDPWR.n1390 VDPWR.n1389 585
R2408 VDPWR.n1389 VDPWR.n1388 585
R2409 VDPWR.n1345 VDPWR.n1342 585
R2410 VDPWR.n1387 VDPWR.n1342 585
R2411 VDPWR.n1385 VDPWR.n1384 585
R2412 VDPWR.n1386 VDPWR.n1385 585
R2413 VDPWR.n1451 VDPWR.n1224 585
R2414 VDPWR.n1449 VDPWR.n1448 585
R2415 VDPWR.n1447 VDPWR.n1230 585
R2416 VDPWR.n1446 VDPWR.n1445 585
R2417 VDPWR.n1443 VDPWR.n1231 585
R2418 VDPWR.n1441 VDPWR.n1440 585
R2419 VDPWR.n1439 VDPWR.n1232 585
R2420 VDPWR.n1438 VDPWR.n1437 585
R2421 VDPWR.n1435 VDPWR.n1233 585
R2422 VDPWR.n1433 VDPWR.n1432 585
R2423 VDPWR.n1431 VDPWR.n1234 585
R2424 VDPWR.n1430 VDPWR.n1429 585
R2425 VDPWR.n1054 VDPWR.n934 585
R2426 VDPWR.n1052 VDPWR.n1051 585
R2427 VDPWR.n1049 VDPWR.n1048 585
R2428 VDPWR.n966 VDPWR.n938 585
R2429 VDPWR.n970 VDPWR.n969 585
R2430 VDPWR.n972 VDPWR.n965 585
R2431 VDPWR.n975 VDPWR.n974 585
R2432 VDPWR.n961 VDPWR.n957 585
R2433 VDPWR.n985 VDPWR.n984 585
R2434 VDPWR.n987 VDPWR.n956 585
R2435 VDPWR.n991 VDPWR.n990 585
R2436 VDPWR.n988 VDPWR.n885 585
R2437 VDPWR.n1427 VDPWR.n1426 585
R2438 VDPWR.n1425 VDPWR.n1424 585
R2439 VDPWR.n1423 VDPWR.n1422 585
R2440 VDPWR.n1421 VDPWR.n1420 585
R2441 VDPWR.n1419 VDPWR.n1418 585
R2442 VDPWR.n1417 VDPWR.n1416 585
R2443 VDPWR.n1415 VDPWR.n1414 585
R2444 VDPWR.n1413 VDPWR.n1412 585
R2445 VDPWR.n1411 VDPWR.n1410 585
R2446 VDPWR.n1409 VDPWR.n1408 585
R2447 VDPWR.n1407 VDPWR.n1406 585
R2448 VDPWR.n1685 VDPWR.n915 585
R2449 VDPWR.n1687 VDPWR.n913 585
R2450 VDPWR.n1055 VDPWR.n914 585
R2451 VDPWR.n1057 VDPWR.n1056 585
R2452 VDPWR.n1059 VDPWR.n1058 585
R2453 VDPWR.n1061 VDPWR.n1060 585
R2454 VDPWR.n1063 VDPWR.n1062 585
R2455 VDPWR.n1065 VDPWR.n1064 585
R2456 VDPWR.n1067 VDPWR.n1066 585
R2457 VDPWR.n1069 VDPWR.n1068 585
R2458 VDPWR.n1071 VDPWR.n1070 585
R2459 VDPWR.n1073 VDPWR.n1072 585
R2460 VDPWR.n1685 VDPWR.n1076 585
R2461 VDPWR.n1685 VDPWR.n1684 585
R2462 VDPWR.n1685 VDPWR.n922 585
R2463 VDPWR.n1132 VDPWR.n1131 585
R2464 VDPWR.n1129 VDPWR.n1128 585
R2465 VDPWR.n1193 VDPWR.n1192 585
R2466 VDPWR.n1195 VDPWR.n1127 585
R2467 VDPWR.n1198 VDPWR.n1197 585
R2468 VDPWR.n1125 VDPWR.n1124 585
R2469 VDPWR.n1205 VDPWR.n1204 585
R2470 VDPWR.n1207 VDPWR.n1122 585
R2471 VDPWR.n1210 VDPWR.n1209 585
R2472 VDPWR.n1102 VDPWR.n1101 585
R2473 VDPWR.n1218 VDPWR.n1217 585
R2474 VDPWR.n1221 VDPWR.n1220 585
R2475 VDPWR.n1663 VDPWR.n928 585
R2476 VDPWR.n1685 VDPWR.n928 585
R2477 VDPWR.n1665 VDPWR.n1664 585
R2478 VDPWR.n1667 VDPWR.n1666 585
R2479 VDPWR.n1669 VDPWR.n1668 585
R2480 VDPWR.n1671 VDPWR.n1670 585
R2481 VDPWR.n1673 VDPWR.n1672 585
R2482 VDPWR.n1675 VDPWR.n1674 585
R2483 VDPWR.n1677 VDPWR.n1676 585
R2484 VDPWR.n1679 VDPWR.n1678 585
R2485 VDPWR.n1681 VDPWR.n1680 585
R2486 VDPWR.n1683 VDPWR.n1682 585
R2487 VDPWR.n1642 VDPWR.n1641 585
R2488 VDPWR.n1644 VDPWR.n1085 585
R2489 VDPWR.n1646 VDPWR.n1645 585
R2490 VDPWR.n1647 VDPWR.n1084 585
R2491 VDPWR.n1649 VDPWR.n1648 585
R2492 VDPWR.n1651 VDPWR.n1082 585
R2493 VDPWR.n1653 VDPWR.n1652 585
R2494 VDPWR.n1654 VDPWR.n1081 585
R2495 VDPWR.n1656 VDPWR.n1655 585
R2496 VDPWR.n1658 VDPWR.n1080 585
R2497 VDPWR.n1659 VDPWR.n1079 585
R2498 VDPWR.n1662 VDPWR.n1661 585
R2499 VDPWR.n2454 VDPWR.n2453 585
R2500 VDPWR.n2454 VDPWR.n22 585
R2501 VDPWR.n2452 VDPWR.n848 585
R2502 VDPWR.n2448 VDPWR.n848 585
R2503 VDPWR.n2451 VDPWR.n2450 585
R2504 VDPWR.n2450 VDPWR.n2449 585
R2505 VDPWR.n850 VDPWR.n849 585
R2506 VDPWR.n851 VDPWR.n850 585
R2507 VDPWR.n1826 VDPWR.n1825 585
R2508 VDPWR.n1827 VDPWR.n1826 585
R2509 VDPWR.n1824 VDPWR.n862 585
R2510 VDPWR.n862 VDPWR.n21 585
R2511 VDPWR.n1823 VDPWR.n1822 585
R2512 VDPWR.n1822 VDPWR.n20 585
R2513 VDPWR.n1821 VDPWR.n863 585
R2514 VDPWR.n1821 VDPWR.n1820 585
R2515 VDPWR.n1804 VDPWR.n864 585
R2516 VDPWR.n865 VDPWR.n864 585
R2517 VDPWR.n1806 VDPWR.n1805 585
R2518 VDPWR.n1807 VDPWR.n1806 585
R2519 VDPWR.n1803 VDPWR.n881 585
R2520 VDPWR.n881 VDPWR.n880 585
R2521 VDPWR.n1802 VDPWR.n1801 585
R2522 VDPWR.n1801 VDPWR.n1800 585
R2523 VDPWR.n1639 VDPWR.n883 585
R2524 VDPWR.n1638 VDPWR.n1090 585
R2525 VDPWR.n1630 VDPWR.n1088 585
R2526 VDPWR.n1633 VDPWR.n1632 585
R2527 VDPWR.n1629 VDPWR.n1092 585
R2528 VDPWR.n1627 VDPWR.n1626 585
R2529 VDPWR.n1094 VDPWR.n1093 585
R2530 VDPWR.n1620 VDPWR.n1619 585
R2531 VDPWR.n1617 VDPWR.n1096 585
R2532 VDPWR.n1615 VDPWR.n1614 585
R2533 VDPWR.n1098 VDPWR.n1097 585
R2534 VDPWR.n1608 VDPWR.n1607 585
R2535 VDPWR.n1605 VDPWR.n1604 585
R2536 VDPWR.n1605 VDPWR.n45 585
R2537 VDPWR.n1640 VDPWR.n1639 585
R2538 VDPWR.n1638 VDPWR.n1637 585
R2539 VDPWR.n1636 VDPWR.n1088 585
R2540 VDPWR.n1634 VDPWR.n1633 585
R2541 VDPWR.n1092 VDPWR.n1091 585
R2542 VDPWR.n1626 VDPWR.n1625 585
R2543 VDPWR.n1623 VDPWR.n1094 585
R2544 VDPWR.n1621 VDPWR.n1620 585
R2545 VDPWR.n1096 VDPWR.n1095 585
R2546 VDPWR.n1614 VDPWR.n1613 585
R2547 VDPWR.n1611 VDPWR.n1098 585
R2548 VDPWR.n1609 VDPWR.n1608 585
R2549 VDPWR.n1604 VDPWR.n1099 585
R2550 VDPWR.n1099 VDPWR.n43 585
R2551 VDPWR.n1712 VDPWR.n73 585
R2552 VDPWR.n911 VDPWR.n910 585
R2553 VDPWR.n1717 VDPWR.n908 585
R2554 VDPWR.n1718 VDPWR.n906 585
R2555 VDPWR.n1719 VDPWR.n905 585
R2556 VDPWR.n903 VDPWR.n900 585
R2557 VDPWR.n1724 VDPWR.n899 585
R2558 VDPWR.n1725 VDPWR.n897 585
R2559 VDPWR.n1726 VDPWR.n896 585
R2560 VDPWR.n894 VDPWR.n890 585
R2561 VDPWR.n893 VDPWR.n888 585
R2562 VDPWR.n1733 VDPWR.n887 585
R2563 VDPWR.n886 VDPWR.n884 585
R2564 VDPWR.n884 VDPWR.n45 585
R2565 VDPWR.n1713 VDPWR.n1712 585
R2566 VDPWR.n1715 VDPWR.n911 585
R2567 VDPWR.n1717 VDPWR.n1716 585
R2568 VDPWR.n1718 VDPWR.n902 585
R2569 VDPWR.n1720 VDPWR.n1719 585
R2570 VDPWR.n1722 VDPWR.n900 585
R2571 VDPWR.n1724 VDPWR.n1723 585
R2572 VDPWR.n1725 VDPWR.n891 585
R2573 VDPWR.n1727 VDPWR.n1726 585
R2574 VDPWR.n1729 VDPWR.n890 585
R2575 VDPWR.n1730 VDPWR.n888 585
R2576 VDPWR.n1733 VDPWR.n1732 585
R2577 VDPWR.n889 VDPWR.n886 585
R2578 VDPWR.n889 VDPWR.n43 585
R2579 VDPWR.n1799 VDPWR.n1798 585
R2580 VDPWR.n1800 VDPWR.n1799 585
R2581 VDPWR.n879 VDPWR.n878 585
R2582 VDPWR.n880 VDPWR.n879 585
R2583 VDPWR.n1809 VDPWR.n1808 585
R2584 VDPWR.n1808 VDPWR.n1807 585
R2585 VDPWR.n875 VDPWR.n866 585
R2586 VDPWR.n866 VDPWR.n865 585
R2587 VDPWR.n1819 VDPWR.n1818 585
R2588 VDPWR.n1820 VDPWR.n1819 585
R2589 VDPWR.n869 VDPWR.n867 585
R2590 VDPWR.n867 VDPWR.n20 585
R2591 VDPWR.n872 VDPWR.n861 585
R2592 VDPWR.n861 VDPWR.n21 585
R2593 VDPWR.n1828 VDPWR.n860 585
R2594 VDPWR.n1828 VDPWR.n1827 585
R2595 VDPWR.n1830 VDPWR.n1829 585
R2596 VDPWR.n1829 VDPWR.n851 585
R2597 VDPWR.n857 VDPWR.n852 585
R2598 VDPWR.n2449 VDPWR.n852 585
R2599 VDPWR.n2447 VDPWR.n2446 585
R2600 VDPWR.n2448 VDPWR.n2447 585
R2601 VDPWR.n2444 VDPWR.n853 585
R2602 VDPWR.n853 VDPWR.n22 585
R2603 VDPWR.n2259 VDPWR.n1839 585
R2604 VDPWR.n2260 VDPWR.n2259 585
R2605 VDPWR.n2122 VDPWR.n2121 585
R2606 VDPWR.n2123 VDPWR.n2122 585
R2607 VDPWR.n2269 VDPWR.n2268 585
R2608 VDPWR.n2268 VDPWR.n2267 585
R2609 VDPWR.n2055 VDPWR.n2045 585
R2610 VDPWR.n2045 VDPWR.n2044 585
R2611 VDPWR.n2279 VDPWR.n2278 585
R2612 VDPWR.n2280 VDPWR.n2279 585
R2613 VDPWR.n2048 VDPWR.n2046 585
R2614 VDPWR.n2046 VDPWR.n26 585
R2615 VDPWR.n2052 VDPWR.n2051 585
R2616 VDPWR.n2051 VDPWR.n27 585
R2617 VDPWR.n2038 VDPWR.n2037 585
R2618 VDPWR.n2039 VDPWR.n2038 585
R2619 VDPWR.n2291 VDPWR.n2290 585
R2620 VDPWR.n2290 VDPWR.n2289 585
R2621 VDPWR.n2034 VDPWR.n2029 585
R2622 VDPWR.n2029 VDPWR.n2028 585
R2623 VDPWR.n2324 VDPWR.n2323 585
R2624 VDPWR.n2325 VDPWR.n2324 585
R2625 VDPWR.n2321 VDPWR.n2030 585
R2626 VDPWR.n2030 VDPWR.n28 585
R2627 VDPWR.n2384 VDPWR.n1883 585
R2628 VDPWR.n2421 VDPWR.n1868 585
R2629 VDPWR.n1866 VDPWR.n1863 585
R2630 VDPWR.n2426 VDPWR.n1862 585
R2631 VDPWR.n2427 VDPWR.n1860 585
R2632 VDPWR.n2428 VDPWR.n1859 585
R2633 VDPWR.n1857 VDPWR.n1854 585
R2634 VDPWR.n2433 VDPWR.n1853 585
R2635 VDPWR.n2434 VDPWR.n1851 585
R2636 VDPWR.n2435 VDPWR.n1850 585
R2637 VDPWR.n1848 VDPWR.n1844 585
R2638 VDPWR.n1847 VDPWR.n1842 585
R2639 VDPWR.n2442 VDPWR.n1841 585
R2640 VDPWR.n2258 VDPWR.n1840 585
R2641 VDPWR.n2258 VDPWR.n36 585
R2642 VDPWR.n2422 VDPWR.n2421 585
R2643 VDPWR.n2424 VDPWR.n1863 585
R2644 VDPWR.n2426 VDPWR.n2425 585
R2645 VDPWR.n2427 VDPWR.n1856 585
R2646 VDPWR.n2429 VDPWR.n2428 585
R2647 VDPWR.n2431 VDPWR.n1854 585
R2648 VDPWR.n2433 VDPWR.n2432 585
R2649 VDPWR.n2434 VDPWR.n1845 585
R2650 VDPWR.n2436 VDPWR.n2435 585
R2651 VDPWR.n2438 VDPWR.n1844 585
R2652 VDPWR.n2439 VDPWR.n1842 585
R2653 VDPWR.n2442 VDPWR.n2441 585
R2654 VDPWR.n1843 VDPWR.n1840 585
R2655 VDPWR.n1843 VDPWR.n34 585
R2656 VDPWR.n2419 VDPWR.n1865 585
R2657 VDPWR.n2418 VDPWR.n2417 585
R2658 VDPWR.n2416 VDPWR.n64 585
R2659 VDPWR.n2640 VDPWR.n64 585
R2660 VDPWR.n2415 VDPWR.n2414 585
R2661 VDPWR.n2413 VDPWR.n2412 585
R2662 VDPWR.n2411 VDPWR.n76 585
R2663 VDPWR.n2630 VDPWR.n2629 585
R2664 VDPWR.n2632 VDPWR.n2631 585
R2665 VDPWR.n2634 VDPWR.n2633 585
R2666 VDPWR.n2636 VDPWR.n2635 585
R2667 VDPWR.n2637 VDPWR.n74 585
R2668 VDPWR.n2639 VDPWR.n2638 585
R2669 VDPWR.n2640 VDPWR.n2639 585
R2670 VDPWR.n2621 VDPWR.n78 585
R2671 VDPWR.n2627 VDPWR.n77 585
R2672 VDPWR.n77 VDPWR.n72 585
R2673 VDPWR.t235 VDPWR.n20 580.369
R2674 VDPWR.t235 VDPWR.n23 580.369
R2675 VDPWR.t235 VDPWR.n26 580.369
R2676 VDPWR.t235 VDPWR.n29 580.369
R2677 VDPWR.n2742 VDPWR.t292 576.699
R2678 VDPWR.t125 VDPWR.n2741 576.699
R2679 VDPWR.n2741 VDPWR.t133 576.699
R2680 VDPWR.t306 VDPWR.n2738 576.699
R2681 VDPWR.n2737 VDPWR.t224 576.699
R2682 VDPWR.n2736 VDPWR.t20 576.699
R2683 VDPWR.n2735 VDPWR.t78 576.699
R2684 VDPWR.n591 VDPWR.t321 566.966
R2685 VDPWR.t235 VDPWR.t72 541.827
R2686 VDPWR.t235 VDPWR.t96 541.827
R2687 VDPWR.n2739 VDPWR.t62 533.981
R2688 VDPWR.n293 VDPWR.t94 524.22
R2689 VDPWR.t183 VDPWR.t110 523.244
R2690 VDPWR.t146 VDPWR.n14 520.611
R2691 VDPWR.t315 VDPWR.n16 520.611
R2692 VDPWR.n690 VDPWR.t228 520.611
R2693 VDPWR.t148 VDPWR.n583 487.568
R2694 VDPWR.t292 VDPWR.t83 469.904
R2695 VDPWR.t26 VDPWR.t125 469.904
R2696 VDPWR.t133 VDPWR.t14 469.904
R2697 VDPWR.t62 VDPWR.t306 469.904
R2698 VDPWR.t224 VDPWR.t70 469.904
R2699 VDPWR.t181 VDPWR.n421 463.784
R2700 VDPWR.t201 VDPWR.n457 459.776
R2701 VDPWR.t107 VDPWR.n463 459.776
R2702 VDPWR.t36 VDPWR.t50 454.832
R2703 VDPWR.t30 VDPWR.t42 449.502
R2704 VDPWR.t7 VDPWR.n17 433.072
R2705 VDPWR.t78 VDPWR.n2734 422.62
R2706 VDPWR.t42 VDPWR.n2724 415.76
R2707 VDPWR.n584 VDPWR.t222 392.433
R2708 VDPWR.t43 VDPWR.t31 380.541
R2709 VDPWR.t255 VDPWR.t143 378.125
R2710 VDPWR.n2730 VDPWR.n17 347.368
R2711 VDPWR.n276 VDPWR.t284 336.329
R2712 VDPWR.n276 VDPWR.t238 336.329
R2713 VDPWR.n333 VDPWR.t250 336.329
R2714 VDPWR.n333 VDPWR.t254 336.329
R2715 VDPWR.t140 VDPWR.t218 332.974
R2716 VDPWR.t235 VDPWR.n49 324.967
R2717 VDPWR.n1800 VDPWR.t235 323.926
R2718 VDPWR.n1600 VDPWR.t235 323.926
R2719 VDPWR.n2260 VDPWR.t235 323.926
R2720 VDPWR.t235 VDPWR.n2257 323.926
R2721 VDPWR.t58 VDPWR.n92 321.082
R2722 VDPWR.n358 VDPWR.t260 320.7
R2723 VDPWR.n302 VDPWR.t268 320.7
R2724 VDPWR.t68 VDPWR.t10 317.969
R2725 VDPWR.t310 VDPWR.t196 317.969
R2726 VDPWR.t5 VDPWR.t261 317.969
R2727 VDPWR.n292 VDPWR.t116 309.375
R2728 VDPWR.n368 VDPWR.t251 309.375
R2729 VDPWR.t110 VDPWR.t56 309.19
R2730 VDPWR.n284 VDPWR.n272 305
R2731 VDPWR.n278 VDPWR.n275 305
R2732 VDPWR.n341 VDPWR.n331 305
R2733 VDPWR.n335 VDPWR.n334 305
R2734 VDPWR.n2721 VDPWR.t264 304.634
R2735 VDPWR.n2660 VDPWR.t276 304.634
R2736 VDPWR.n2666 VDPWR.t247 304.634
R2737 VDPWR.n2717 VDPWR.t280 304.634
R2738 VDPWR.n133 VDPWR.t141 302.334
R2739 VDPWR.n102 VDPWR.t168 302.334
R2740 VDPWR.n100 VDPWR.t149 302.334
R2741 VDPWR.n451 VDPWR.t103 301.574
R2742 VDPWR.n2712 VDPWR.t272 292.584
R2743 VDPWR.n2674 VDPWR.t244 292.584
R2744 VDPWR.n366 VDPWR.n365 292.188
R2745 VDPWR.n2672 VDPWR.n2657 275.8
R2746 VDPWR.t153 VDPWR.n582 273.514
R2747 VDPWR.t24 VDPWR.n446 270.493
R2748 VDPWR.t235 VDPWR.n22 269.94
R2749 VDPWR.t235 VDPWR.n25 269.94
R2750 VDPWR.t235 VDPWR.n28 269.94
R2751 VDPWR.t235 VDPWR.n31 269.94
R2752 VDPWR.n2622 VDPWR.n72 267.485
R2753 VDPWR.t31 VDPWR.t140 261.623
R2754 VDPWR.t218 VDPWR.t87 261.623
R2755 VDPWR.t294 VDPWR.t85 261.623
R2756 VDPWR.t165 VDPWR.t47 261.623
R2757 VDPWR.t18 VDPWR.t76 261.623
R2758 VDPWR.n582 VDPWR.n94 261.623
R2759 VDPWR.t314 VDPWR.t123 261.623
R2760 VDPWR.n124 VDPWR.n123 260.199
R2761 VDPWR.n2615 VDPWR.t73 260
R2762 VDPWR.t73 VDPWR.n2612 260
R2763 VDPWR.n467 VDPWR.t136 260
R2764 VDPWR.n465 VDPWR.t136 260
R2765 VDPWR.n2669 VDPWR.n2668 259.844
R2766 VDPWR.n2639 VDPWR.n73 259.416
R2767 VDPWR.n1429 VDPWR.n1427 259.416
R2768 VDPWR.n2256 VDPWR.n814 259.416
R2769 VDPWR.n2261 VDPWR.n845 259.416
R2770 VDPWR.n1801 VDPWR.n883 259.416
R2771 VDPWR.n1601 VDPWR.n1458 259.416
R2772 VDPWR.n1688 VDPWR.n1687 259.416
R2773 VDPWR.n2409 VDPWR.n1868 259.416
R2774 VDPWR.n1661 VDPWR.n928 259.416
R2775 VDPWR.n2086 VDPWR.n2085 258.334
R2776 VDPWR.n1763 VDPWR.n1762 258.334
R2777 VDPWR.n2199 VDPWR.n2198 258.334
R2778 VDPWR.n1942 VDPWR.n1941 258.334
R2779 VDPWR.n1544 VDPWR.n1543 258.334
R2780 VDPWR.n766 VDPWR.n765 258.334
R2781 VDPWR.n1303 VDPWR.n1302 258.334
R2782 VDPWR.n1011 VDPWR.n950 258.334
R2783 VDPWR.n1151 VDPWR.n1150 258.334
R2784 VDPWR.n813 VDPWR.n36 254.34
R2785 VDPWR.n807 VDPWR.n36 254.34
R2786 VDPWR.n804 VDPWR.n36 254.34
R2787 VDPWR.n798 VDPWR.n36 254.34
R2788 VDPWR.n795 VDPWR.n36 254.34
R2789 VDPWR.n792 VDPWR.n36 254.34
R2790 VDPWR.n844 VDPWR.n36 254.34
R2791 VDPWR.n841 VDPWR.n36 254.34
R2792 VDPWR.n835 VDPWR.n36 254.34
R2793 VDPWR.n832 VDPWR.n36 254.34
R2794 VDPWR.n826 VDPWR.n36 254.34
R2795 VDPWR.n823 VDPWR.n36 254.34
R2796 VDPWR.n2481 VDPWR.n34 254.34
R2797 VDPWR.n810 VDPWR.n34 254.34
R2798 VDPWR.n2488 VDPWR.n34 254.34
R2799 VDPWR.n801 VDPWR.n34 254.34
R2800 VDPWR.n2495 VDPWR.n34 254.34
R2801 VDPWR.n2498 VDPWR.n34 254.34
R2802 VDPWR.n847 VDPWR.n34 254.34
R2803 VDPWR.n2460 VDPWR.n34 254.34
R2804 VDPWR.n838 VDPWR.n34 254.34
R2805 VDPWR.n2467 VDPWR.n34 254.34
R2806 VDPWR.n829 VDPWR.n34 254.34
R2807 VDPWR.n2474 VDPWR.n34 254.34
R2808 VDPWR.n1457 VDPWR.n45 254.34
R2809 VDPWR.n1366 VDPWR.n45 254.34
R2810 VDPWR.n1364 VDPWR.n45 254.34
R2811 VDPWR.n1357 VDPWR.n45 254.34
R2812 VDPWR.n1354 VDPWR.n45 254.34
R2813 VDPWR.n1348 VDPWR.n45 254.34
R2814 VDPWR.n1453 VDPWR.n43 254.34
R2815 VDPWR.n1361 VDPWR.n43 254.34
R2816 VDPWR.n1371 VDPWR.n43 254.34
R2817 VDPWR.n1360 VDPWR.n43 254.34
R2818 VDPWR.n1378 VDPWR.n43 254.34
R2819 VDPWR.n1351 VDPWR.n43 254.34
R2820 VDPWR.n2640 VDPWR.n71 254.34
R2821 VDPWR.n2640 VDPWR.n70 254.34
R2822 VDPWR.n2640 VDPWR.n69 254.34
R2823 VDPWR.n2640 VDPWR.n68 254.34
R2824 VDPWR.n2640 VDPWR.n67 254.34
R2825 VDPWR.n2640 VDPWR.n66 254.34
R2826 VDPWR.n2640 VDPWR.n59 254.34
R2827 VDPWR.n2640 VDPWR.n58 254.34
R2828 VDPWR.n2640 VDPWR.n57 254.34
R2829 VDPWR.n2640 VDPWR.n56 254.34
R2830 VDPWR.n2640 VDPWR.n55 254.34
R2831 VDPWR.n2640 VDPWR.n54 254.34
R2832 VDPWR.n2384 VDPWR.n1884 254.34
R2833 VDPWR.n2384 VDPWR.n1885 254.34
R2834 VDPWR.n2384 VDPWR.n1886 254.34
R2835 VDPWR.n2384 VDPWR.n1887 254.34
R2836 VDPWR.n2384 VDPWR.n1888 254.34
R2837 VDPWR.n2384 VDPWR.n1889 254.34
R2838 VDPWR.n2382 VDPWR.n2381 254.34
R2839 VDPWR.n2384 VDPWR.n1876 254.34
R2840 VDPWR.n2384 VDPWR.n1875 254.34
R2841 VDPWR.n2384 VDPWR.n1874 254.34
R2842 VDPWR.n2384 VDPWR.n1873 254.34
R2843 VDPWR.n2384 VDPWR.n1872 254.34
R2844 VDPWR.n2384 VDPWR.n1871 254.34
R2845 VDPWR.n2385 VDPWR.n2384 254.34
R2846 VDPWR.n2384 VDPWR.n1882 254.34
R2847 VDPWR.n2384 VDPWR.n1881 254.34
R2848 VDPWR.n2384 VDPWR.n1880 254.34
R2849 VDPWR.n2384 VDPWR.n1879 254.34
R2850 VDPWR.n1450 VDPWR.n39 254.34
R2851 VDPWR.n1444 VDPWR.n39 254.34
R2852 VDPWR.n1442 VDPWR.n39 254.34
R2853 VDPWR.n1436 VDPWR.n39 254.34
R2854 VDPWR.n1434 VDPWR.n39 254.34
R2855 VDPWR.n1428 VDPWR.n39 254.34
R2856 VDPWR.n1050 VDPWR.n50 254.34
R2857 VDPWR.n937 VDPWR.n50 254.34
R2858 VDPWR.n971 VDPWR.n50 254.34
R2859 VDPWR.n973 VDPWR.n50 254.34
R2860 VDPWR.n986 VDPWR.n50 254.34
R2861 VDPWR.n989 VDPWR.n50 254.34
R2862 VDPWR.n1685 VDPWR.n921 254.34
R2863 VDPWR.n1685 VDPWR.n920 254.34
R2864 VDPWR.n1685 VDPWR.n919 254.34
R2865 VDPWR.n1685 VDPWR.n918 254.34
R2866 VDPWR.n1685 VDPWR.n917 254.34
R2867 VDPWR.n1685 VDPWR.n916 254.34
R2868 VDPWR.n1405 VDPWR.n1235 254.34
R2869 VDPWR.n1686 VDPWR.n1685 254.34
R2870 VDPWR.n1685 VDPWR.n929 254.34
R2871 VDPWR.n1685 VDPWR.n930 254.34
R2872 VDPWR.n1685 VDPWR.n931 254.34
R2873 VDPWR.n1685 VDPWR.n932 254.34
R2874 VDPWR.n1685 VDPWR.n933 254.34
R2875 VDPWR.n1075 VDPWR.n1074 254.34
R2876 VDPWR.n1078 VDPWR.n1077 254.34
R2877 VDPWR.n1130 VDPWR.n42 254.34
R2878 VDPWR.n1194 VDPWR.n42 254.34
R2879 VDPWR.n1196 VDPWR.n42 254.34
R2880 VDPWR.n1206 VDPWR.n42 254.34
R2881 VDPWR.n1208 VDPWR.n42 254.34
R2882 VDPWR.n1219 VDPWR.n42 254.34
R2883 VDPWR.n1685 VDPWR.n927 254.34
R2884 VDPWR.n1685 VDPWR.n926 254.34
R2885 VDPWR.n1685 VDPWR.n925 254.34
R2886 VDPWR.n1685 VDPWR.n924 254.34
R2887 VDPWR.n1685 VDPWR.n923 254.34
R2888 VDPWR.n1643 VDPWR.n41 254.34
R2889 VDPWR.n1086 VDPWR.n41 254.34
R2890 VDPWR.n1650 VDPWR.n41 254.34
R2891 VDPWR.n1083 VDPWR.n41 254.34
R2892 VDPWR.n1657 VDPWR.n41 254.34
R2893 VDPWR.n1660 VDPWR.n41 254.34
R2894 VDPWR.n1089 VDPWR.n45 254.34
R2895 VDPWR.n1631 VDPWR.n45 254.34
R2896 VDPWR.n1628 VDPWR.n45 254.34
R2897 VDPWR.n1618 VDPWR.n45 254.34
R2898 VDPWR.n1616 VDPWR.n45 254.34
R2899 VDPWR.n1606 VDPWR.n45 254.34
R2900 VDPWR.n1087 VDPWR.n43 254.34
R2901 VDPWR.n1635 VDPWR.n43 254.34
R2902 VDPWR.n1624 VDPWR.n43 254.34
R2903 VDPWR.n1622 VDPWR.n43 254.34
R2904 VDPWR.n1612 VDPWR.n43 254.34
R2905 VDPWR.n1610 VDPWR.n43 254.34
R2906 VDPWR.n909 VDPWR.n45 254.34
R2907 VDPWR.n907 VDPWR.n45 254.34
R2908 VDPWR.n904 VDPWR.n45 254.34
R2909 VDPWR.n898 VDPWR.n45 254.34
R2910 VDPWR.n895 VDPWR.n45 254.34
R2911 VDPWR.n892 VDPWR.n45 254.34
R2912 VDPWR.n1714 VDPWR.n43 254.34
R2913 VDPWR.n912 VDPWR.n43 254.34
R2914 VDPWR.n1721 VDPWR.n43 254.34
R2915 VDPWR.n901 VDPWR.n43 254.34
R2916 VDPWR.n1728 VDPWR.n43 254.34
R2917 VDPWR.n1731 VDPWR.n43 254.34
R2918 VDPWR.n2320 VDPWR.n2300 254.34
R2919 VDPWR.n2384 VDPWR.n1878 254.34
R2920 VDPWR.n1867 VDPWR.n36 254.34
R2921 VDPWR.n1861 VDPWR.n36 254.34
R2922 VDPWR.n1858 VDPWR.n36 254.34
R2923 VDPWR.n1852 VDPWR.n36 254.34
R2924 VDPWR.n1849 VDPWR.n36 254.34
R2925 VDPWR.n1846 VDPWR.n36 254.34
R2926 VDPWR.n2423 VDPWR.n34 254.34
R2927 VDPWR.n1864 VDPWR.n34 254.34
R2928 VDPWR.n2430 VDPWR.n34 254.34
R2929 VDPWR.n1855 VDPWR.n34 254.34
R2930 VDPWR.n2437 VDPWR.n34 254.34
R2931 VDPWR.n2440 VDPWR.n34 254.34
R2932 VDPWR.n2640 VDPWR.n65 254.34
R2933 VDPWR.n2640 VDPWR.n63 254.34
R2934 VDPWR.n2640 VDPWR.n62 254.34
R2935 VDPWR.n2640 VDPWR.n61 254.34
R2936 VDPWR.n2640 VDPWR.n60 254.34
R2937 VDPWR.n126 VDPWR.n125 254.333
R2938 VDPWR.n139 VDPWR.n138 254.333
R2939 VDPWR.n117 VDPWR.n116 254.333
R2940 VDPWR.n150 VDPWR.n114 254.333
R2941 VDPWR.n109 VDPWR.n108 254.333
R2942 VDPWR.n164 VDPWR.n163 254.333
R2943 VDPWR.n190 VDPWR.n189 254.333
R2944 VDPWR.n196 VDPWR.n195 254.333
R2945 VDPWR.n569 VDPWR.n204 254.333
R2946 VDPWR.n206 VDPWR.n205 254.333
R2947 VDPWR.n557 VDPWR.n210 253.114
R2948 VDPWR.n2422 VDPWR.n1865 251.614
R2949 VDPWR.n1452 VDPWR.n1451 251.614
R2950 VDPWR.n2359 VDPWR.n2358 251.614
R2951 VDPWR.n2327 VDPWR.n1877 251.614
R2952 VDPWR.n2455 VDPWR.n2454 251.614
R2953 VDPWR.n2480 VDPWR.n811 251.614
R2954 VDPWR.n1713 VDPWR.n1711 251.614
R2955 VDPWR.n2387 VDPWR.n2386 251.614
R2956 VDPWR.n1642 VDPWR.n1640 251.614
R2957 VDPWR.n365 VDPWR.n364 250.349
R2958 VDPWR.n365 VDPWR.n258 250.349
R2959 VDPWR.n367 VDPWR.n257 250.349
R2960 VDPWR.n367 VDPWR.n256 250.349
R2961 VDPWR.n277 VDPWR.n255 250.349
R2962 VDPWR.n283 VDPWR.n255 250.349
R2963 VDPWR.n295 VDPWR.n293 250.349
R2964 VDPWR.n300 VDPWR.n293 250.349
R2965 VDPWR.n2544 VDPWR.n2535 250.349
R2966 VDPWR.n2559 VDPWR.n2558 250.349
R2967 VDPWR.n442 VDPWR.t64 249.731
R2968 VDPWR.n2577 VDPWR.n2574 246.25
R2969 VDPWR.n2585 VDPWR.n2574 246.25
R2970 VDPWR.n2606 VDPWR.n2596 246.25
R2971 VDPWR.n2607 VDPWR.n2606 246.25
R2972 VDPWR.n2722 VDPWR.t267 245
R2973 VDPWR.n2658 VDPWR.t278 245
R2974 VDPWR.n2667 VDPWR.t248 245
R2975 VDPWR.n2716 VDPWR.t282 245
R2976 VDPWR.n470 VDPWR.n464 241.643
R2977 VDPWR.n463 VDPWR.n458 241.643
R2978 VDPWR.n457 VDPWR.n452 241.643
R2979 VDPWR.n2614 VDPWR.n2613 241.643
R2980 VDPWR.n2608 VDPWR.t0 241.643
R2981 VDPWR.n2599 VDPWR.t0 241.643
R2982 VDPWR.n2586 VDPWR.t98 241.643
R2983 VDPWR.n2578 VDPWR.t98 241.643
R2984 VDPWR.n450 VDPWR.n255 240.625
R2985 VDPWR.n584 VDPWR.n92 237.839
R2986 VDPWR.t81 VDPWR.t18 237.839
R2987 VDPWR.t163 VDPWR.t209 236.281
R2988 VDPWR.n170 VDPWR.t59 233
R2989 VDPWR.n581 VDPWR.t124 233
R2990 VDPWR.n461 VDPWR.t202 233
R2991 VDPWR.n468 VDPWR.t204 233
R2992 VDPWR.n455 VDPWR.t198 233
R2993 VDPWR.n550 VDPWR.n215 225.534
R2994 VDPWR.n219 VDPWR.n218 225.534
R2995 VDPWR.n538 VDPWR.n222 225.534
R2996 VDPWR.n531 VDPWR.n227 225.534
R2997 VDPWR.n231 VDPWR.n230 225.534
R2998 VDPWR.n512 VDPWR.n238 225.534
R2999 VDPWR.n243 VDPWR.n242 225.534
R3000 VDPWR.n500 VDPWR.n499 225.534
R3001 VDPWR.n519 VDPWR.n234 225.534
R3002 VDPWR.t184 VDPWR.n9 218.321
R3003 VDPWR.t190 VDPWR.t177 214.054
R3004 VDPWR.t226 VDPWR.t43 214.054
R3005 VDPWR.t87 VDPWR.t158 214.054
R3006 VDPWR.t64 VDPWR.t99 214.054
R3007 VDPWR.n2664 VDPWR.n2663 210.601
R3008 VDPWR.n2662 VDPWR.n2661 210.601
R3009 VDPWR.n2665 VDPWR.n2659 210.601
R3010 VDPWR.n650 VDPWR.t63 204.458
R3011 VDPWR.n645 VDPWR.t15 204.458
R3012 VDPWR.n637 VDPWR.t27 204.458
R3013 VDPWR.n632 VDPWR.t84 204.458
R3014 VDPWR.n387 VDPWR.t44 204.458
R3015 VDPWR.n392 VDPWR.t219 204.458
R3016 VDPWR.n377 VDPWR.t40 204.458
R3017 VDPWR.n406 VDPWR.t161 204.458
R3018 VDPWR.n2719 VDPWR.n2643 204.201
R3019 VDPWR.n2718 VDPWR.n2644 204.201
R3020 VDPWR.n2720 VDPWR.n2641 204.201
R3021 VDPWR.n2668 VDPWR.t28 203.913
R3022 VDPWR.n422 VDPWR.t162 202.162
R3023 VDPWR.n2557 VDPWR.n703 197
R3024 VDPWR.n2543 VDPWR.n2536 197
R3025 VDPWR.n299 VDPWR.n294 197
R3026 VDPWR.n282 VDPWR.n274 197
R3027 VDPWR.n337 VDPWR.n336 197
R3028 VDPWR.n360 VDPWR.n259 197
R3029 VDPWR.t76 VDPWR.t153 190.27
R3030 VDPWR.t290 VDPWR.t52 190.27
R3031 VDPWR.t45 VDPWR.t105 189.062
R3032 VDPWR.t3 VDPWR.t45 189.062
R3033 VDPWR.t317 VDPWR.t220 189.062
R3034 VDPWR.t232 VDPWR.t212 189.062
R3035 VDPWR.t214 VDPWR.t216 189.062
R3036 VDPWR.t211 VDPWR.t37 189.062
R3037 VDPWR.t22 VDPWR.t32 189.062
R3038 VDPWR.t54 VDPWR.t108 189.062
R3039 VDPWR.t298 VDPWR.t101 189.062
R3040 VDPWR.n2085 VDPWR.n2067 185
R3041 VDPWR.n2083 VDPWR.n2082 185
R3042 VDPWR.n2081 VDPWR.n2069 185
R3043 VDPWR.n2080 VDPWR.n2079 185
R3044 VDPWR.n2077 VDPWR.n2070 185
R3045 VDPWR.n2075 VDPWR.n2074 185
R3046 VDPWR.n2073 VDPWR.n2072 185
R3047 VDPWR.n2033 VDPWR.n2032 185
R3048 VDPWR.n2299 VDPWR.n2298 185
R3049 VDPWR.n2087 VDPWR.n2086 185
R3050 VDPWR.n2088 VDPWR.n2066 185
R3051 VDPWR.n2090 VDPWR.n2089 185
R3052 VDPWR.n2092 VDPWR.n2064 185
R3053 VDPWR.n2094 VDPWR.n2093 185
R3054 VDPWR.n2095 VDPWR.n2063 185
R3055 VDPWR.n2097 VDPWR.n2096 185
R3056 VDPWR.n2099 VDPWR.n2062 185
R3057 VDPWR.n2102 VDPWR.n2101 185
R3058 VDPWR.n2103 VDPWR.n2061 185
R3059 VDPWR.n2105 VDPWR.n2104 185
R3060 VDPWR.n2107 VDPWR.n2060 185
R3061 VDPWR.n2110 VDPWR.n2109 185
R3062 VDPWR.n2111 VDPWR.n2059 185
R3063 VDPWR.n2113 VDPWR.n2112 185
R3064 VDPWR.n2115 VDPWR.n2058 185
R3065 VDPWR.n2118 VDPWR.n2117 185
R3066 VDPWR.n2119 VDPWR.n2057 185
R3067 VDPWR.n1762 VDPWR.n1744 185
R3068 VDPWR.n1760 VDPWR.n1759 185
R3069 VDPWR.n1758 VDPWR.n1746 185
R3070 VDPWR.n1757 VDPWR.n1756 185
R3071 VDPWR.n1754 VDPWR.n1747 185
R3072 VDPWR.n1752 VDPWR.n1751 185
R3073 VDPWR.n1750 VDPWR.n1749 185
R3074 VDPWR.n856 VDPWR.n855 185
R3075 VDPWR.n1838 VDPWR.n1837 185
R3076 VDPWR.n1764 VDPWR.n1763 185
R3077 VDPWR.n1765 VDPWR.n1743 185
R3078 VDPWR.n1767 VDPWR.n1766 185
R3079 VDPWR.n1769 VDPWR.n1741 185
R3080 VDPWR.n1771 VDPWR.n1770 185
R3081 VDPWR.n1772 VDPWR.n1740 185
R3082 VDPWR.n1774 VDPWR.n1773 185
R3083 VDPWR.n1776 VDPWR.n1739 185
R3084 VDPWR.n1779 VDPWR.n1778 185
R3085 VDPWR.n1780 VDPWR.n1738 185
R3086 VDPWR.n1782 VDPWR.n1781 185
R3087 VDPWR.n1784 VDPWR.n1737 185
R3088 VDPWR.n1787 VDPWR.n1786 185
R3089 VDPWR.n1788 VDPWR.n1736 185
R3090 VDPWR.n1790 VDPWR.n1789 185
R3091 VDPWR.n1792 VDPWR.n1735 185
R3092 VDPWR.n1795 VDPWR.n1794 185
R3093 VDPWR.n1796 VDPWR.n877 185
R3094 VDPWR.n2587 VDPWR.n2573 185
R3095 VDPWR.n2580 VDPWR.n2579 185
R3096 VDPWR.n2598 VDPWR.n2594 185
R3097 VDPWR.n2600 VDPWR.n2598 185
R3098 VDPWR.n2198 VDPWR.n2148 185
R3099 VDPWR.n2196 VDPWR.n2195 185
R3100 VDPWR.n2194 VDPWR.n2150 185
R3101 VDPWR.n2193 VDPWR.n2192 185
R3102 VDPWR.n2190 VDPWR.n2151 185
R3103 VDPWR.n2188 VDPWR.n2187 185
R3104 VDPWR.n2186 VDPWR.n2152 185
R3105 VDPWR.n2185 VDPWR.n2184 185
R3106 VDPWR.n2182 VDPWR.n2024 185
R3107 VDPWR.n2200 VDPWR.n2199 185
R3108 VDPWR.n2201 VDPWR.n2147 185
R3109 VDPWR.n2203 VDPWR.n2202 185
R3110 VDPWR.n2205 VDPWR.n2145 185
R3111 VDPWR.n2207 VDPWR.n2206 185
R3112 VDPWR.n2208 VDPWR.n2144 185
R3113 VDPWR.n2210 VDPWR.n2209 185
R3114 VDPWR.n2212 VDPWR.n2143 185
R3115 VDPWR.n2215 VDPWR.n2214 185
R3116 VDPWR.n2216 VDPWR.n2142 185
R3117 VDPWR.n2218 VDPWR.n2217 185
R3118 VDPWR.n2220 VDPWR.n2141 185
R3119 VDPWR.n2223 VDPWR.n2222 185
R3120 VDPWR.n2224 VDPWR.n2140 185
R3121 VDPWR.n2226 VDPWR.n2225 185
R3122 VDPWR.n2228 VDPWR.n2139 185
R3123 VDPWR.n2231 VDPWR.n2230 185
R3124 VDPWR.n2232 VDPWR.n2138 185
R3125 VDPWR.n1941 VDPWR.n1919 185
R3126 VDPWR.n1939 VDPWR.n1938 185
R3127 VDPWR.n1937 VDPWR.n1921 185
R3128 VDPWR.n1936 VDPWR.n1935 185
R3129 VDPWR.n1933 VDPWR.n1922 185
R3130 VDPWR.n1931 VDPWR.n1930 185
R3131 VDPWR.n1929 VDPWR.n1923 185
R3132 VDPWR.n1928 VDPWR.n1927 185
R3133 VDPWR.n1925 VDPWR.n1891 185
R3134 VDPWR.n1943 VDPWR.n1942 185
R3135 VDPWR.n1944 VDPWR.n1918 185
R3136 VDPWR.n1946 VDPWR.n1945 185
R3137 VDPWR.n1948 VDPWR.n1916 185
R3138 VDPWR.n1950 VDPWR.n1949 185
R3139 VDPWR.n1951 VDPWR.n1915 185
R3140 VDPWR.n1953 VDPWR.n1952 185
R3141 VDPWR.n1955 VDPWR.n1914 185
R3142 VDPWR.n1958 VDPWR.n1957 185
R3143 VDPWR.n1959 VDPWR.n1913 185
R3144 VDPWR.n1961 VDPWR.n1960 185
R3145 VDPWR.n1963 VDPWR.n1912 185
R3146 VDPWR.n1966 VDPWR.n1965 185
R3147 VDPWR.n1967 VDPWR.n1911 185
R3148 VDPWR.n1969 VDPWR.n1968 185
R3149 VDPWR.n1971 VDPWR.n1910 185
R3150 VDPWR.n1974 VDPWR.n1973 185
R3151 VDPWR.n1975 VDPWR.n1909 185
R3152 VDPWR.n1986 VDPWR.n1985 185
R3153 VDPWR.n1988 VDPWR.n1906 185
R3154 VDPWR.n1991 VDPWR.n1990 185
R3155 VDPWR.n1907 VDPWR.n1901 185
R3156 VDPWR.n2001 VDPWR.n2000 185
R3157 VDPWR.n2003 VDPWR.n1900 185
R3158 VDPWR.n2004 VDPWR.n1896 185
R3159 VDPWR.n2007 VDPWR.n2006 185
R3160 VDPWR.n1898 VDPWR.n1892 185
R3161 VDPWR.n1543 VDPWR.n1483 185
R3162 VDPWR.n1541 VDPWR.n1540 185
R3163 VDPWR.n1539 VDPWR.n1485 185
R3164 VDPWR.n1538 VDPWR.n1537 185
R3165 VDPWR.n1535 VDPWR.n1486 185
R3166 VDPWR.n1533 VDPWR.n1532 185
R3167 VDPWR.n1531 VDPWR.n1487 185
R3168 VDPWR.n1530 VDPWR.n1529 185
R3169 VDPWR.n1527 VDPWR.n1488 185
R3170 VDPWR.n1545 VDPWR.n1544 185
R3171 VDPWR.n1546 VDPWR.n1482 185
R3172 VDPWR.n1548 VDPWR.n1547 185
R3173 VDPWR.n1550 VDPWR.n1480 185
R3174 VDPWR.n1552 VDPWR.n1551 185
R3175 VDPWR.n1553 VDPWR.n1479 185
R3176 VDPWR.n1555 VDPWR.n1554 185
R3177 VDPWR.n1557 VDPWR.n1478 185
R3178 VDPWR.n1560 VDPWR.n1559 185
R3179 VDPWR.n1561 VDPWR.n1477 185
R3180 VDPWR.n1563 VDPWR.n1562 185
R3181 VDPWR.n1565 VDPWR.n1476 185
R3182 VDPWR.n1568 VDPWR.n1567 185
R3183 VDPWR.n1569 VDPWR.n1475 185
R3184 VDPWR.n1571 VDPWR.n1570 185
R3185 VDPWR.n1573 VDPWR.n1474 185
R3186 VDPWR.n1576 VDPWR.n1575 185
R3187 VDPWR.n1577 VDPWR.n1473 185
R3188 VDPWR.n1583 VDPWR.n1582 185
R3189 VDPWR.n1585 VDPWR.n1472 185
R3190 VDPWR.n1586 VDPWR.n1468 185
R3191 VDPWR.n1589 VDPWR.n1588 185
R3192 VDPWR.n1503 VDPWR.n1470 185
R3193 VDPWR.n1508 VDPWR.n1506 185
R3194 VDPWR.n1511 VDPWR.n1510 185
R3195 VDPWR.n1512 VDPWR.n1489 185
R3196 VDPWR.n1525 VDPWR.n1524 185
R3197 VDPWR.n767 VDPWR.n766 185
R3198 VDPWR.n769 VDPWR.n768 185
R3199 VDPWR.n771 VDPWR.n770 185
R3200 VDPWR.n773 VDPWR.n772 185
R3201 VDPWR.n775 VDPWR.n774 185
R3202 VDPWR.n777 VDPWR.n776 185
R3203 VDPWR.n779 VDPWR.n778 185
R3204 VDPWR.n781 VDPWR.n780 185
R3205 VDPWR.n782 VDPWR.n728 185
R3206 VDPWR.n765 VDPWR.n764 185
R3207 VDPWR.n763 VDPWR.n762 185
R3208 VDPWR.n761 VDPWR.n760 185
R3209 VDPWR.n759 VDPWR.n758 185
R3210 VDPWR.n757 VDPWR.n756 185
R3211 VDPWR.n755 VDPWR.n754 185
R3212 VDPWR.n753 VDPWR.n752 185
R3213 VDPWR.n751 VDPWR.n750 185
R3214 VDPWR.n749 VDPWR.n748 185
R3215 VDPWR.n747 VDPWR.n746 185
R3216 VDPWR.n745 VDPWR.n744 185
R3217 VDPWR.n743 VDPWR.n742 185
R3218 VDPWR.n741 VDPWR.n740 185
R3219 VDPWR.n739 VDPWR.n738 185
R3220 VDPWR.n737 VDPWR.n736 185
R3221 VDPWR.n735 VDPWR.n734 185
R3222 VDPWR.n733 VDPWR.n732 185
R3223 VDPWR.n731 VDPWR.n710 185
R3224 VDPWR.n1304 VDPWR.n1303 185
R3225 VDPWR.n1306 VDPWR.n1305 185
R3226 VDPWR.n1308 VDPWR.n1307 185
R3227 VDPWR.n1310 VDPWR.n1309 185
R3228 VDPWR.n1312 VDPWR.n1311 185
R3229 VDPWR.n1314 VDPWR.n1313 185
R3230 VDPWR.n1316 VDPWR.n1315 185
R3231 VDPWR.n1318 VDPWR.n1317 185
R3232 VDPWR.n1319 VDPWR.n1261 185
R3233 VDPWR.n1302 VDPWR.n1301 185
R3234 VDPWR.n1300 VDPWR.n1299 185
R3235 VDPWR.n1298 VDPWR.n1297 185
R3236 VDPWR.n1296 VDPWR.n1295 185
R3237 VDPWR.n1294 VDPWR.n1293 185
R3238 VDPWR.n1292 VDPWR.n1291 185
R3239 VDPWR.n1290 VDPWR.n1289 185
R3240 VDPWR.n1288 VDPWR.n1287 185
R3241 VDPWR.n1286 VDPWR.n1285 185
R3242 VDPWR.n1284 VDPWR.n1283 185
R3243 VDPWR.n1282 VDPWR.n1281 185
R3244 VDPWR.n1280 VDPWR.n1279 185
R3245 VDPWR.n1278 VDPWR.n1277 185
R3246 VDPWR.n1276 VDPWR.n1275 185
R3247 VDPWR.n1274 VDPWR.n1273 185
R3248 VDPWR.n1272 VDPWR.n1271 185
R3249 VDPWR.n1270 VDPWR.n1269 185
R3250 VDPWR.n1268 VDPWR.n1267 185
R3251 VDPWR.n1266 VDPWR.n1265 185
R3252 VDPWR.n1243 VDPWR.n1241 185
R3253 VDPWR.n1396 VDPWR.n1395 185
R3254 VDPWR.n1324 VDPWR.n1244 185
R3255 VDPWR.n1328 VDPWR.n1327 185
R3256 VDPWR.n1333 VDPWR.n1330 185
R3257 VDPWR.n1335 VDPWR.n1334 185
R3258 VDPWR.n1331 VDPWR.n1262 185
R3259 VDPWR.n1392 VDPWR.n1391 185
R3260 VDPWR.n2553 VDPWR.n2552 185
R3261 VDPWR.n2509 VDPWR.n711 185
R3262 VDPWR.n2515 VDPWR.n2514 185
R3263 VDPWR.n2519 VDPWR.n2518 185
R3264 VDPWR.n2517 VDPWR.n2507 185
R3265 VDPWR.n2526 VDPWR.n2525 185
R3266 VDPWR.n2528 VDPWR.n2527 185
R3267 VDPWR.n2529 VDPWR.n729 185
R3268 VDPWR.n2549 VDPWR.n2548 185
R3269 VDPWR.n2240 VDPWR.n2239 185
R3270 VDPWR.n2242 VDPWR.n2137 185
R3271 VDPWR.n2243 VDPWR.n2133 185
R3272 VDPWR.n2246 VDPWR.n2245 185
R3273 VDPWR.n2158 VDPWR.n2135 185
R3274 VDPWR.n2159 VDPWR.n2156 185
R3275 VDPWR.n2177 VDPWR.n2176 185
R3276 VDPWR.n2179 VDPWR.n2154 185
R3277 VDPWR.n2180 VDPWR.n2023 185
R3278 VDPWR.n1009 VDPWR.n950 185
R3279 VDPWR.n1008 VDPWR.n1007 185
R3280 VDPWR.n1005 VDPWR.n951 185
R3281 VDPWR.n1003 VDPWR.n1002 185
R3282 VDPWR.n1001 VDPWR.n952 185
R3283 VDPWR.n1000 VDPWR.n999 185
R3284 VDPWR.n997 VDPWR.n953 185
R3285 VDPWR.n995 VDPWR.n994 185
R3286 VDPWR.n993 VDPWR.n954 185
R3287 VDPWR.n1011 VDPWR.n1010 185
R3288 VDPWR.n1013 VDPWR.n948 185
R3289 VDPWR.n1015 VDPWR.n1014 185
R3290 VDPWR.n1016 VDPWR.n947 185
R3291 VDPWR.n1018 VDPWR.n1017 185
R3292 VDPWR.n1020 VDPWR.n945 185
R3293 VDPWR.n1022 VDPWR.n1021 185
R3294 VDPWR.n1023 VDPWR.n944 185
R3295 VDPWR.n1025 VDPWR.n1024 185
R3296 VDPWR.n1027 VDPWR.n943 185
R3297 VDPWR.n1030 VDPWR.n1029 185
R3298 VDPWR.n1031 VDPWR.n942 185
R3299 VDPWR.n1033 VDPWR.n1032 185
R3300 VDPWR.n1035 VDPWR.n941 185
R3301 VDPWR.n1038 VDPWR.n1037 185
R3302 VDPWR.n1039 VDPWR.n940 185
R3303 VDPWR.n1041 VDPWR.n1040 185
R3304 VDPWR.n1043 VDPWR.n935 185
R3305 VDPWR.n1044 VDPWR.n936 185
R3306 VDPWR.n1047 VDPWR.n1046 185
R3307 VDPWR.n967 VDPWR.n939 185
R3308 VDPWR.n968 VDPWR.n964 185
R3309 VDPWR.n977 VDPWR.n976 185
R3310 VDPWR.n979 VDPWR.n962 185
R3311 VDPWR.n980 VDPWR.n958 185
R3312 VDPWR.n983 VDPWR.n982 185
R3313 VDPWR.n960 VDPWR.n955 185
R3314 VDPWR.n280 VDPWR.n275 185
R3315 VDPWR.n281 VDPWR.n272 185
R3316 VDPWR.n338 VDPWR.n335 185
R3317 VDPWR.n332 VDPWR.n331 185
R3318 VDPWR.n1150 VDPWR.n1149 185
R3319 VDPWR.n1148 VDPWR.n1147 185
R3320 VDPWR.n1146 VDPWR.n1145 185
R3321 VDPWR.n1144 VDPWR.n1143 185
R3322 VDPWR.n1142 VDPWR.n1141 185
R3323 VDPWR.n1140 VDPWR.n1139 185
R3324 VDPWR.n1138 VDPWR.n1137 185
R3325 VDPWR.n1136 VDPWR.n1135 185
R3326 VDPWR.n1134 VDPWR.n1104 185
R3327 VDPWR.n1152 VDPWR.n1151 185
R3328 VDPWR.n1154 VDPWR.n1153 185
R3329 VDPWR.n1156 VDPWR.n1155 185
R3330 VDPWR.n1158 VDPWR.n1157 185
R3331 VDPWR.n1160 VDPWR.n1159 185
R3332 VDPWR.n1162 VDPWR.n1161 185
R3333 VDPWR.n1164 VDPWR.n1163 185
R3334 VDPWR.n1166 VDPWR.n1165 185
R3335 VDPWR.n1168 VDPWR.n1167 185
R3336 VDPWR.n1170 VDPWR.n1169 185
R3337 VDPWR.n1172 VDPWR.n1171 185
R3338 VDPWR.n1174 VDPWR.n1173 185
R3339 VDPWR.n1176 VDPWR.n1175 185
R3340 VDPWR.n1178 VDPWR.n1177 185
R3341 VDPWR.n1180 VDPWR.n1179 185
R3342 VDPWR.n1182 VDPWR.n1181 185
R3343 VDPWR.n1184 VDPWR.n1183 185
R3344 VDPWR.n1186 VDPWR.n1185 185
R3345 VDPWR.n1188 VDPWR.n1187 185
R3346 VDPWR.n1191 VDPWR.n1190 185
R3347 VDPWR.n1189 VDPWR.n1126 185
R3348 VDPWR.n1200 VDPWR.n1199 185
R3349 VDPWR.n1202 VDPWR.n1201 185
R3350 VDPWR.n1203 VDPWR.n1121 185
R3351 VDPWR.n1212 VDPWR.n1211 185
R3352 VDPWR.n1123 VDPWR.n1103 185
R3353 VDPWR.n1216 VDPWR.n1215 185
R3354 VDPWR.n1811 VDPWR.n1810 185
R3355 VDPWR.n1813 VDPWR.n876 185
R3356 VDPWR.n1814 VDPWR.n868 185
R3357 VDPWR.n1817 VDPWR.n1816 185
R3358 VDPWR.n874 VDPWR.n873 185
R3359 VDPWR.n871 VDPWR.n859 185
R3360 VDPWR.n1832 VDPWR.n1831 185
R3361 VDPWR.n1834 VDPWR.n858 185
R3362 VDPWR.n1835 VDPWR.n854 185
R3363 VDPWR.n2271 VDPWR.n2270 185
R3364 VDPWR.n2273 VDPWR.n2056 185
R3365 VDPWR.n2274 VDPWR.n2047 185
R3366 VDPWR.n2277 VDPWR.n2276 185
R3367 VDPWR.n2054 VDPWR.n2053 185
R3368 VDPWR.n2050 VDPWR.n2036 185
R3369 VDPWR.n2293 VDPWR.n2292 185
R3370 VDPWR.n2295 VDPWR.n2035 185
R3371 VDPWR.n2296 VDPWR.n2031 185
R3372 VDPWR.n2639 VDPWR.n74 175.546
R3373 VDPWR.n2635 VDPWR.n2634 175.546
R3374 VDPWR.n2631 VDPWR.n2630 175.546
R3375 VDPWR.n2412 VDPWR.n2411 175.546
R3376 VDPWR.n2414 VDPWR.n64 175.546
R3377 VDPWR.n2417 VDPWR.n64 175.546
R3378 VDPWR.n2441 VDPWR.n1843 175.546
R3379 VDPWR.n2439 VDPWR.n2438 175.546
R3380 VDPWR.n2436 VDPWR.n1845 175.546
R3381 VDPWR.n2432 VDPWR.n2431 175.546
R3382 VDPWR.n2429 VDPWR.n1856 175.546
R3383 VDPWR.n2425 VDPWR.n2424 175.546
R3384 VDPWR.n1799 VDPWR.n879 175.546
R3385 VDPWR.n1808 VDPWR.n879 175.546
R3386 VDPWR.n1808 VDPWR.n866 175.546
R3387 VDPWR.n1819 VDPWR.n866 175.546
R3388 VDPWR.n1819 VDPWR.n867 175.546
R3389 VDPWR.n867 VDPWR.n861 175.546
R3390 VDPWR.n1828 VDPWR.n861 175.546
R3391 VDPWR.n1829 VDPWR.n1828 175.546
R3392 VDPWR.n1829 VDPWR.n852 175.546
R3393 VDPWR.n2447 VDPWR.n852 175.546
R3394 VDPWR.n2447 VDPWR.n853 175.546
R3395 VDPWR.n887 VDPWR.n884 175.546
R3396 VDPWR.n894 VDPWR.n893 175.546
R3397 VDPWR.n897 VDPWR.n896 175.546
R3398 VDPWR.n903 VDPWR.n899 175.546
R3399 VDPWR.n906 VDPWR.n905 175.546
R3400 VDPWR.n910 VDPWR.n908 175.546
R3401 VDPWR.n1403 VDPWR.n1402 175.546
R3402 VDPWR.n1402 VDPWR.n1237 175.546
R3403 VDPWR.n1398 VDPWR.n1237 175.546
R3404 VDPWR.n1398 VDPWR.n1240 175.546
R3405 VDPWR.n1325 VDPWR.n1240 175.546
R3406 VDPWR.n1325 VDPWR.n1323 175.546
R3407 VDPWR.n1337 VDPWR.n1323 175.546
R3408 VDPWR.n1337 VDPWR.n1321 175.546
R3409 VDPWR.n1341 VDPWR.n1321 175.546
R3410 VDPWR.n1389 VDPWR.n1341 175.546
R3411 VDPWR.n1389 VDPWR.n1342 175.546
R3412 VDPWR.n1408 VDPWR.n1407 175.546
R3413 VDPWR.n1412 VDPWR.n1411 175.546
R3414 VDPWR.n1416 VDPWR.n1415 175.546
R3415 VDPWR.n1420 VDPWR.n1419 175.546
R3416 VDPWR.n1424 VDPWR.n1423 175.546
R3417 VDPWR.n1433 VDPWR.n1234 175.546
R3418 VDPWR.n1437 VDPWR.n1435 175.546
R3419 VDPWR.n1441 VDPWR.n1232 175.546
R3420 VDPWR.n1445 VDPWR.n1443 175.546
R3421 VDPWR.n1449 VDPWR.n1230 175.546
R3422 VDPWR.n1385 VDPWR.n1343 175.546
R3423 VDPWR.n1380 VDPWR.n1379 175.546
R3424 VDPWR.n1377 VDPWR.n1352 175.546
R3425 VDPWR.n1373 VDPWR.n1372 175.546
R3426 VDPWR.n1370 VDPWR.n1362 175.546
R3427 VDPWR.n1454 VDPWR.n1229 175.546
R3428 VDPWR.n1978 VDPWR.n788 175.546
R3429 VDPWR.n794 VDPWR.n793 175.546
R3430 VDPWR.n797 VDPWR.n796 175.546
R3431 VDPWR.n803 VDPWR.n799 175.546
R3432 VDPWR.n806 VDPWR.n805 175.546
R3433 VDPWR.n812 VDPWR.n808 175.546
R3434 VDPWR.n1982 VDPWR.n1977 175.546
R3435 VDPWR.n1982 VDPWR.n1905 175.546
R3436 VDPWR.n1993 VDPWR.n1905 175.546
R3437 VDPWR.n1993 VDPWR.n1903 175.546
R3438 VDPWR.n1997 VDPWR.n1903 175.546
R3439 VDPWR.n1998 VDPWR.n1997 175.546
R3440 VDPWR.n1998 VDPWR.n1895 175.546
R3441 VDPWR.n2009 VDPWR.n1895 175.546
R3442 VDPWR.n2009 VDPWR.n1893 175.546
R3443 VDPWR.n2013 VDPWR.n1893 175.546
R3444 VDPWR.n2013 VDPWR.n1890 175.546
R3445 VDPWR.n2379 VDPWR.n2378 175.546
R3446 VDPWR.n2375 VDPWR.n2374 175.546
R3447 VDPWR.n2371 VDPWR.n2370 175.546
R3448 VDPWR.n2367 VDPWR.n2366 175.546
R3449 VDPWR.n2363 VDPWR.n2362 175.546
R3450 VDPWR.n2256 VDPWR.n2255 175.546
R3451 VDPWR.n2255 VDPWR.n2127 175.546
R3452 VDPWR.n2251 VDPWR.n2127 175.546
R3453 VDPWR.n2251 VDPWR.n2129 175.546
R3454 VDPWR.n2166 VDPWR.n2129 175.546
R3455 VDPWR.n2167 VDPWR.n2166 175.546
R3456 VDPWR.n2167 VDPWR.n2164 175.546
R3457 VDPWR.n2172 VDPWR.n2164 175.546
R3458 VDPWR.n2172 VDPWR.n2018 175.546
R3459 VDPWR.n2357 VDPWR.n2018 175.546
R3460 VDPWR.n2358 VDPWR.n2357 175.546
R3461 VDPWR.n822 VDPWR.n817 175.546
R3462 VDPWR.n825 VDPWR.n824 175.546
R3463 VDPWR.n831 VDPWR.n827 175.546
R3464 VDPWR.n834 VDPWR.n833 175.546
R3465 VDPWR.n840 VDPWR.n836 175.546
R3466 VDPWR.n843 VDPWR.n842 175.546
R3467 VDPWR.n2236 VDPWR.n2125 175.546
R3468 VDPWR.n2237 VDPWR.n2236 175.546
R3469 VDPWR.n2237 VDPWR.n2131 175.546
R3470 VDPWR.n2248 VDPWR.n2131 175.546
R3471 VDPWR.n2248 VDPWR.n2132 175.546
R3472 VDPWR.n2161 VDPWR.n2132 175.546
R3473 VDPWR.n2162 VDPWR.n2161 175.546
R3474 VDPWR.n2174 VDPWR.n2162 175.546
R3475 VDPWR.n2174 VDPWR.n2021 175.546
R3476 VDPWR.n2355 VDPWR.n2021 175.546
R3477 VDPWR.n2355 VDPWR.n2022 175.546
R3478 VDPWR.n2348 VDPWR.n2025 175.546
R3479 VDPWR.n2346 VDPWR.n2345 175.546
R3480 VDPWR.n2342 VDPWR.n2341 175.546
R3481 VDPWR.n2338 VDPWR.n2337 175.546
R3482 VDPWR.n2334 VDPWR.n2333 175.546
R3483 VDPWR.n2330 VDPWR.n1877 175.546
R3484 VDPWR.n2261 VDPWR.n2124 175.546
R3485 VDPWR.n2266 VDPWR.n2124 175.546
R3486 VDPWR.n2266 VDPWR.n2042 175.546
R3487 VDPWR.n2281 VDPWR.n2042 175.546
R3488 VDPWR.n2282 VDPWR.n2281 175.546
R3489 VDPWR.n2283 VDPWR.n2282 175.546
R3490 VDPWR.n2283 VDPWR.n2040 175.546
R3491 VDPWR.n2288 VDPWR.n2040 175.546
R3492 VDPWR.n2288 VDPWR.n2027 175.546
R3493 VDPWR.n2326 VDPWR.n2027 175.546
R3494 VDPWR.n2327 VDPWR.n2326 175.546
R3495 VDPWR.n1607 VDPWR.n1605 175.546
R3496 VDPWR.n1615 VDPWR.n1097 175.546
R3497 VDPWR.n1619 VDPWR.n1617 175.546
R3498 VDPWR.n1627 VDPWR.n1093 175.546
R3499 VDPWR.n1632 VDPWR.n1629 175.546
R3500 VDPWR.n1630 VDPWR.n1090 175.546
R3501 VDPWR.n1801 VDPWR.n881 175.546
R3502 VDPWR.n1806 VDPWR.n881 175.546
R3503 VDPWR.n1806 VDPWR.n864 175.546
R3504 VDPWR.n1821 VDPWR.n864 175.546
R3505 VDPWR.n1822 VDPWR.n1821 175.546
R3506 VDPWR.n1822 VDPWR.n862 175.546
R3507 VDPWR.n1826 VDPWR.n862 175.546
R3508 VDPWR.n1826 VDPWR.n850 175.546
R3509 VDPWR.n2450 VDPWR.n850 175.546
R3510 VDPWR.n2450 VDPWR.n848 175.546
R3511 VDPWR.n2454 VDPWR.n848 175.546
R3512 VDPWR.n2476 VDPWR.n2475 175.546
R3513 VDPWR.n2473 VDPWR.n821 175.546
R3514 VDPWR.n2469 VDPWR.n2468 175.546
R3515 VDPWR.n2466 VDPWR.n830 175.546
R3516 VDPWR.n2462 VDPWR.n2461 175.546
R3517 VDPWR.n2459 VDPWR.n839 175.546
R3518 VDPWR.n1460 VDPWR.n1223 175.546
R3519 VDPWR.n1461 VDPWR.n1460 175.546
R3520 VDPWR.n1466 VDPWR.n1461 175.546
R3521 VDPWR.n1591 VDPWR.n1466 175.546
R3522 VDPWR.n1591 VDPWR.n1467 175.546
R3523 VDPWR.n1504 VDPWR.n1467 175.546
R3524 VDPWR.n1504 VDPWR.n1501 175.546
R3525 VDPWR.n1514 VDPWR.n1501 175.546
R3526 VDPWR.n1514 VDPWR.n1493 175.546
R3527 VDPWR.n1522 VDPWR.n1493 175.546
R3528 VDPWR.n1522 VDPWR.n819 175.546
R3529 VDPWR.n1347 VDPWR.n1344 175.546
R3530 VDPWR.n1353 VDPWR.n1349 175.546
R3531 VDPWR.n1356 VDPWR.n1355 175.546
R3532 VDPWR.n1363 VDPWR.n1358 175.546
R3533 VDPWR.n1367 VDPWR.n1365 175.546
R3534 VDPWR.n1456 VDPWR.n1227 175.546
R3535 VDPWR.n2555 VDPWR.n706 175.546
R3536 VDPWR.n2555 VDPWR.n707 175.546
R3537 VDPWR.n2512 VDPWR.n707 175.546
R3538 VDPWR.n2512 VDPWR.n2508 175.546
R3539 VDPWR.n2521 VDPWR.n2508 175.546
R3540 VDPWR.n2523 VDPWR.n2521 175.546
R3541 VDPWR.n2523 VDPWR.n2505 175.546
R3542 VDPWR.n2531 VDPWR.n2505 175.546
R3543 VDPWR.n2531 VDPWR.n784 175.546
R3544 VDPWR.n2546 VDPWR.n784 175.546
R3545 VDPWR.n2546 VDPWR.n2503 175.546
R3546 VDPWR.n2499 VDPWR.n785 175.546
R3547 VDPWR.n2497 VDPWR.n2496 175.546
R3548 VDPWR.n2494 VDPWR.n791 175.546
R3549 VDPWR.n2490 VDPWR.n2489 175.546
R3550 VDPWR.n2487 VDPWR.n802 175.546
R3551 VDPWR.n2483 VDPWR.n2482 175.546
R3552 VDPWR.n1601 VDPWR.n1459 175.546
R3553 VDPWR.n1597 VDPWR.n1459 175.546
R3554 VDPWR.n1597 VDPWR.n1463 175.546
R3555 VDPWR.n1593 VDPWR.n1463 175.546
R3556 VDPWR.n1593 VDPWR.n1465 175.546
R3557 VDPWR.n1498 VDPWR.n1465 175.546
R3558 VDPWR.n1499 VDPWR.n1498 175.546
R3559 VDPWR.n1516 VDPWR.n1499 175.546
R3560 VDPWR.n1516 VDPWR.n1495 175.546
R3561 VDPWR.n1520 VDPWR.n1495 175.546
R3562 VDPWR.n1520 VDPWR.n811 175.546
R3563 VDPWR.n1072 VDPWR.n1071 175.546
R3564 VDPWR.n1068 VDPWR.n1067 175.546
R3565 VDPWR.n1064 VDPWR.n1063 175.546
R3566 VDPWR.n1060 VDPWR.n1059 175.546
R3567 VDPWR.n1056 VDPWR.n914 175.546
R3568 VDPWR.n1051 VDPWR.n1049 175.546
R3569 VDPWR.n970 VDPWR.n966 175.546
R3570 VDPWR.n974 VDPWR.n972 175.546
R3571 VDPWR.n985 VDPWR.n957 175.546
R3572 VDPWR.n990 VDPWR.n987 175.546
R3573 VDPWR.n1732 VDPWR.n889 175.546
R3574 VDPWR.n1730 VDPWR.n1729 175.546
R3575 VDPWR.n1727 VDPWR.n891 175.546
R3576 VDPWR.n1723 VDPWR.n1722 175.546
R3577 VDPWR.n1720 VDPWR.n902 175.546
R3578 VDPWR.n1716 VDPWR.n1715 175.546
R3579 VDPWR.n1692 VDPWR.n1691 175.546
R3580 VDPWR.n1696 VDPWR.n1695 175.546
R3581 VDPWR.n1700 VDPWR.n1699 175.546
R3582 VDPWR.n1704 VDPWR.n1703 175.546
R3583 VDPWR.n1708 VDPWR.n1707 175.546
R3584 VDPWR.n2258 VDPWR.n1841 175.546
R3585 VDPWR.n1848 VDPWR.n1847 175.546
R3586 VDPWR.n1851 VDPWR.n1850 175.546
R3587 VDPWR.n1857 VDPWR.n1853 175.546
R3588 VDPWR.n1860 VDPWR.n1859 175.546
R3589 VDPWR.n1866 VDPWR.n1862 175.546
R3590 VDPWR.n2259 VDPWR.n2122 175.546
R3591 VDPWR.n2268 VDPWR.n2122 175.546
R3592 VDPWR.n2268 VDPWR.n2045 175.546
R3593 VDPWR.n2279 VDPWR.n2045 175.546
R3594 VDPWR.n2279 VDPWR.n2046 175.546
R3595 VDPWR.n2051 VDPWR.n2046 175.546
R3596 VDPWR.n2051 VDPWR.n2038 175.546
R3597 VDPWR.n2290 VDPWR.n2038 175.546
R3598 VDPWR.n2290 VDPWR.n2029 175.546
R3599 VDPWR.n2324 VDPWR.n2029 175.546
R3600 VDPWR.n2324 VDPWR.n2030 175.546
R3601 VDPWR.n2318 VDPWR.n2317 175.546
R3602 VDPWR.n2314 VDPWR.n2313 175.546
R3603 VDPWR.n2310 VDPWR.n2309 175.546
R3604 VDPWR.n2306 VDPWR.n2305 175.546
R3605 VDPWR.n2302 VDPWR.n1870 175.546
R3606 VDPWR.n2407 VDPWR.n2406 175.546
R3607 VDPWR.n2403 VDPWR.n2402 175.546
R3608 VDPWR.n2399 VDPWR.n2398 175.546
R3609 VDPWR.n2395 VDPWR.n2394 175.546
R3610 VDPWR.n2391 VDPWR.n2390 175.546
R3611 VDPWR.n1659 VDPWR.n1658 175.546
R3612 VDPWR.n1656 VDPWR.n1081 175.546
R3613 VDPWR.n1652 VDPWR.n1651 175.546
R3614 VDPWR.n1649 VDPWR.n1084 175.546
R3615 VDPWR.n1645 VDPWR.n1644 175.546
R3616 VDPWR.n1609 VDPWR.n1099 175.546
R3617 VDPWR.n1613 VDPWR.n1611 175.546
R3618 VDPWR.n1621 VDPWR.n1095 175.546
R3619 VDPWR.n1625 VDPWR.n1623 175.546
R3620 VDPWR.n1634 VDPWR.n1091 175.546
R3621 VDPWR.n1637 VDPWR.n1636 175.546
R3622 VDPWR.n1193 VDPWR.n1128 175.546
R3623 VDPWR.n1197 VDPWR.n1195 175.546
R3624 VDPWR.n1205 VDPWR.n1124 175.546
R3625 VDPWR.n1209 VDPWR.n1207 175.546
R3626 VDPWR.n1218 VDPWR.n1101 175.546
R3627 VDPWR.n1684 VDPWR.n1683 175.546
R3628 VDPWR.n1680 VDPWR.n1679 175.546
R3629 VDPWR.n1676 VDPWR.n1675 175.546
R3630 VDPWR.n1672 VDPWR.n1671 175.546
R3631 VDPWR.n1668 VDPWR.n1667 175.546
R3632 VDPWR.n1664 VDPWR.n928 175.546
R3633 VDPWR.t240 VDPWR.n273 174.089
R3634 VDPWR.n279 VDPWR.t240 174.089
R3635 VDPWR.n340 VDPWR.t256 174.089
R3636 VDPWR.t256 VDPWR.n339 174.089
R3637 VDPWR.t263 VDPWR.n362 173.506
R3638 VDPWR.n363 VDPWR.t263 173.506
R3639 VDPWR.t270 VDPWR.n290 173.506
R3640 VDPWR.n296 VDPWR.t270 173.506
R3641 VDPWR.t235 VDPWR.n39 173.084
R3642 VDPWR.t235 VDPWR.n41 173.084
R3643 VDPWR.n473 VDPWR.n472 172.888
R3644 VDPWR.t235 VDPWR.n42 172.302
R3645 VDPWR.t235 VDPWR.n50 172.302
R3646 VDPWR.n278 VDPWR.n276 166.63
R3647 VDPWR.n334 VDPWR.n333 166.63
R3648 VDPWR.t34 VDPWR.t12 166.487
R3649 VDPWR.t137 VDPWR.t39 166.487
R3650 VDPWR.t160 VDPWR.t66 166.487
R3651 VDPWR.t129 VDPWR.t120 166.487
R3652 VDPWR.n2271 VDPWR.n2057 163.333
R3653 VDPWR.n1811 VDPWR.n877 163.333
R3654 VDPWR.n2240 VDPWR.n2138 163.333
R3655 VDPWR.n1986 VDPWR.n1909 163.333
R3656 VDPWR.n1583 VDPWR.n1473 163.333
R3657 VDPWR.n2552 VDPWR.n710 163.333
R3658 VDPWR.n1267 VDPWR.n1266 163.333
R3659 VDPWR.n1044 VDPWR.n1043 163.333
R3660 VDPWR.n1187 VDPWR.n1186 163.333
R3661 VDPWR.t212 VDPWR.t285 163.281
R3662 VDPWR.n2621 VDPWR.n77 157.601
R3663 VDPWR.t150 VDPWR.n445 154.595
R3664 VDPWR.n444 VDPWR.t34 154.595
R3665 VDPWR.t120 VDPWR.n443 154.595
R3666 VDPWR.n1235 VDPWR.n916 152.643
R3667 VDPWR.n2382 VDPWR.n1889 152.643
R3668 VDPWR.n1075 VDPWR.n933 152.643
R3669 VDPWR.n2300 VDPWR.n1878 152.643
R3670 VDPWR.n79 VDPWR.t156 151.275
R3671 VDPWR.n2618 VDPWR.t29 151.153
R3672 VDPWR.n2619 VDPWR.t132 150.885
R3673 VDPWR.n79 VDPWR.t164 150.817
R3674 VDPWR.n2274 VDPWR.n2273 150
R3675 VDPWR.n2276 VDPWR.n2054 150
R3676 VDPWR.n2293 VDPWR.n2036 150
R3677 VDPWR.n2296 VDPWR.n2295 150
R3678 VDPWR.n2117 VDPWR.n2115 150
R3679 VDPWR.n2113 VDPWR.n2059 150
R3680 VDPWR.n2109 VDPWR.n2107 150
R3681 VDPWR.n2105 VDPWR.n2061 150
R3682 VDPWR.n2101 VDPWR.n2099 150
R3683 VDPWR.n2097 VDPWR.n2063 150
R3684 VDPWR.n2093 VDPWR.n2092 150
R3685 VDPWR.n2090 VDPWR.n2066 150
R3686 VDPWR.n2298 VDPWR.n2033 150
R3687 VDPWR.n2075 VDPWR.n2072 150
R3688 VDPWR.n2079 VDPWR.n2077 150
R3689 VDPWR.n2083 VDPWR.n2069 150
R3690 VDPWR.n1814 VDPWR.n1813 150
R3691 VDPWR.n1816 VDPWR.n874 150
R3692 VDPWR.n1832 VDPWR.n859 150
R3693 VDPWR.n1835 VDPWR.n1834 150
R3694 VDPWR.n1794 VDPWR.n1792 150
R3695 VDPWR.n1790 VDPWR.n1736 150
R3696 VDPWR.n1786 VDPWR.n1784 150
R3697 VDPWR.n1782 VDPWR.n1738 150
R3698 VDPWR.n1778 VDPWR.n1776 150
R3699 VDPWR.n1774 VDPWR.n1740 150
R3700 VDPWR.n1770 VDPWR.n1769 150
R3701 VDPWR.n1767 VDPWR.n1743 150
R3702 VDPWR.n1837 VDPWR.n856 150
R3703 VDPWR.n1752 VDPWR.n1749 150
R3704 VDPWR.n1756 VDPWR.n1754 150
R3705 VDPWR.n1760 VDPWR.n1746 150
R3706 VDPWR.n2243 VDPWR.n2242 150
R3707 VDPWR.n2245 VDPWR.n2135 150
R3708 VDPWR.n2177 VDPWR.n2156 150
R3709 VDPWR.n2180 VDPWR.n2179 150
R3710 VDPWR.n2230 VDPWR.n2228 150
R3711 VDPWR.n2226 VDPWR.n2140 150
R3712 VDPWR.n2222 VDPWR.n2220 150
R3713 VDPWR.n2218 VDPWR.n2142 150
R3714 VDPWR.n2214 VDPWR.n2212 150
R3715 VDPWR.n2210 VDPWR.n2144 150
R3716 VDPWR.n2206 VDPWR.n2205 150
R3717 VDPWR.n2203 VDPWR.n2147 150
R3718 VDPWR.n2184 VDPWR.n2182 150
R3719 VDPWR.n2188 VDPWR.n2152 150
R3720 VDPWR.n2192 VDPWR.n2190 150
R3721 VDPWR.n2196 VDPWR.n2150 150
R3722 VDPWR.n1990 VDPWR.n1988 150
R3723 VDPWR.n2001 VDPWR.n1901 150
R3724 VDPWR.n2004 VDPWR.n2003 150
R3725 VDPWR.n2006 VDPWR.n1898 150
R3726 VDPWR.n1973 VDPWR.n1971 150
R3727 VDPWR.n1969 VDPWR.n1911 150
R3728 VDPWR.n1965 VDPWR.n1963 150
R3729 VDPWR.n1961 VDPWR.n1913 150
R3730 VDPWR.n1957 VDPWR.n1955 150
R3731 VDPWR.n1953 VDPWR.n1915 150
R3732 VDPWR.n1949 VDPWR.n1948 150
R3733 VDPWR.n1946 VDPWR.n1918 150
R3734 VDPWR.n1927 VDPWR.n1925 150
R3735 VDPWR.n1931 VDPWR.n1923 150
R3736 VDPWR.n1935 VDPWR.n1933 150
R3737 VDPWR.n1939 VDPWR.n1921 150
R3738 VDPWR.n1586 VDPWR.n1585 150
R3739 VDPWR.n1588 VDPWR.n1470 150
R3740 VDPWR.n1510 VDPWR.n1508 150
R3741 VDPWR.n1525 VDPWR.n1489 150
R3742 VDPWR.n1575 VDPWR.n1573 150
R3743 VDPWR.n1571 VDPWR.n1475 150
R3744 VDPWR.n1567 VDPWR.n1565 150
R3745 VDPWR.n1563 VDPWR.n1477 150
R3746 VDPWR.n1559 VDPWR.n1557 150
R3747 VDPWR.n1555 VDPWR.n1479 150
R3748 VDPWR.n1551 VDPWR.n1550 150
R3749 VDPWR.n1548 VDPWR.n1482 150
R3750 VDPWR.n1529 VDPWR.n1527 150
R3751 VDPWR.n1533 VDPWR.n1487 150
R3752 VDPWR.n1537 VDPWR.n1535 150
R3753 VDPWR.n1541 VDPWR.n1485 150
R3754 VDPWR.n2514 VDPWR.n711 150
R3755 VDPWR.n2518 VDPWR.n2517 150
R3756 VDPWR.n2527 VDPWR.n2526 150
R3757 VDPWR.n2549 VDPWR.n729 150
R3758 VDPWR.n734 VDPWR.n733 150
R3759 VDPWR.n738 VDPWR.n737 150
R3760 VDPWR.n742 VDPWR.n741 150
R3761 VDPWR.n746 VDPWR.n745 150
R3762 VDPWR.n750 VDPWR.n749 150
R3763 VDPWR.n754 VDPWR.n753 150
R3764 VDPWR.n758 VDPWR.n757 150
R3765 VDPWR.n762 VDPWR.n761 150
R3766 VDPWR.n780 VDPWR.n728 150
R3767 VDPWR.n778 VDPWR.n777 150
R3768 VDPWR.n774 VDPWR.n773 150
R3769 VDPWR.n770 VDPWR.n769 150
R3770 VDPWR.n1395 VDPWR.n1243 150
R3771 VDPWR.n1327 VDPWR.n1244 150
R3772 VDPWR.n1334 VDPWR.n1333 150
R3773 VDPWR.n1392 VDPWR.n1262 150
R3774 VDPWR.n1271 VDPWR.n1270 150
R3775 VDPWR.n1275 VDPWR.n1274 150
R3776 VDPWR.n1279 VDPWR.n1278 150
R3777 VDPWR.n1283 VDPWR.n1282 150
R3778 VDPWR.n1287 VDPWR.n1286 150
R3779 VDPWR.n1291 VDPWR.n1290 150
R3780 VDPWR.n1295 VDPWR.n1294 150
R3781 VDPWR.n1299 VDPWR.n1298 150
R3782 VDPWR.n1317 VDPWR.n1261 150
R3783 VDPWR.n1315 VDPWR.n1314 150
R3784 VDPWR.n1311 VDPWR.n1310 150
R3785 VDPWR.n1307 VDPWR.n1306 150
R3786 VDPWR.n1046 VDPWR.n939 150
R3787 VDPWR.n977 VDPWR.n964 150
R3788 VDPWR.n980 VDPWR.n979 150
R3789 VDPWR.n982 VDPWR.n960 150
R3790 VDPWR.n1041 VDPWR.n940 150
R3791 VDPWR.n1037 VDPWR.n1035 150
R3792 VDPWR.n1033 VDPWR.n942 150
R3793 VDPWR.n1029 VDPWR.n1027 150
R3794 VDPWR.n1025 VDPWR.n944 150
R3795 VDPWR.n1021 VDPWR.n1020 150
R3796 VDPWR.n1018 VDPWR.n947 150
R3797 VDPWR.n1014 VDPWR.n1013 150
R3798 VDPWR.n995 VDPWR.n954 150
R3799 VDPWR.n999 VDPWR.n997 150
R3800 VDPWR.n1003 VDPWR.n952 150
R3801 VDPWR.n1007 VDPWR.n1005 150
R3802 VDPWR.n1190 VDPWR.n1189 150
R3803 VDPWR.n1201 VDPWR.n1200 150
R3804 VDPWR.n1212 VDPWR.n1121 150
R3805 VDPWR.n1215 VDPWR.n1103 150
R3806 VDPWR.n1183 VDPWR.n1182 150
R3807 VDPWR.n1179 VDPWR.n1178 150
R3808 VDPWR.n1175 VDPWR.n1174 150
R3809 VDPWR.n1171 VDPWR.n1170 150
R3810 VDPWR.n1167 VDPWR.n1166 150
R3811 VDPWR.n1163 VDPWR.n1162 150
R3812 VDPWR.n1159 VDPWR.n1158 150
R3813 VDPWR.n1155 VDPWR.n1154 150
R3814 VDPWR.n1135 VDPWR.n1104 150
R3815 VDPWR.n1139 VDPWR.n1138 150
R3816 VDPWR.n1143 VDPWR.n1142 150
R3817 VDPWR.n1147 VDPWR.n1146 150
R3818 VDPWR.t94 VDPWR.n291 146.095
R3819 VDPWR.t216 VDPWR.n255 146.095
R3820 VDPWR.t32 VDPWR.n367 146.095
R3821 VDPWR.n704 VDPWR.n44 146.041
R3822 VDPWR.n1799 VDPWR.n884 144.338
R3823 VDPWR.n1403 VDPWR.n915 144.338
R3824 VDPWR.n1978 VDPWR.n1977 144.338
R3825 VDPWR.n2125 VDPWR.n817 144.338
R3826 VDPWR.n1605 VDPWR.n1223 144.338
R3827 VDPWR.n1344 VDPWR.n706 144.338
R3828 VDPWR.n1076 VDPWR.n934 144.338
R3829 VDPWR.n2259 VDPWR.n2258 144.338
R3830 VDPWR.n1131 VDPWR.n922 144.338
R3831 VDPWR.n2534 VDPWR.n35 138.81
R3832 VDPWR.n2728 VDPWR.n17 137.243
R3833 VDPWR.n1843 VDPWR.n853 136.536
R3834 VDPWR.n1385 VDPWR.n1342 136.536
R3835 VDPWR.n2383 VDPWR.n1890 136.536
R3836 VDPWR.n2350 VDPWR.n2022 136.536
R3837 VDPWR.n2476 VDPWR.n819 136.536
R3838 VDPWR.n2503 VDPWR.n785 136.536
R3839 VDPWR.n988 VDPWR.n889 136.536
R3840 VDPWR.n2030 VDPWR.n1883 136.536
R3841 VDPWR.n1220 VDPWR.n1099 136.536
R3842 VDPWR.t16 VDPWR.n1979 135.919
R3843 VDPWR.n2713 VDPWR.t275 134.501
R3844 VDPWR.t113 VDPWR.n1386 134.474
R3845 VDPWR.n2603 VDPWR.n2595 134.268
R3846 VDPWR.n2598 VDPWR.n2595 134.268
R3847 VDPWR.n457 VDPWR.t36 133.483
R3848 VDPWR.n463 VDPWR.t201 133.483
R3849 VDPWR.n470 VDPWR.t107 133.483
R3850 VDPWR.t127 VDPWR.n470 133.483
R3851 VDPWR.n2656 VDPWR.t245 132.058
R3852 VDPWR.n379 VDPWR.t88 130.713
R3853 VDPWR.n2725 VDPWR.t30 130.314
R3854 VDPWR.n1400 VDPWR.n1399 130.136
R3855 VDPWR.n1338 VDPWR.n1322 130.136
R3856 VDPWR.n1388 VDPWR.n1387 130.136
R3857 VDPWR.n2556 VDPWR.n705 130.136
R3858 VDPWR.n2511 VDPWR.n705 130.136
R3859 VDPWR.n2511 VDPWR.n2510 130.136
R3860 VDPWR.n2510 VDPWR.n32 130.136
R3861 VDPWR.n2522 VDPWR.n2504 130.136
R3862 VDPWR.n2532 VDPWR.n2504 130.136
R3863 VDPWR.n2533 VDPWR.n2532 130.136
R3864 VDPWR.n2545 VDPWR.n2533 130.136
R3865 VDPWR.n1981 VDPWR.n1980 130.136
R3866 VDPWR.n1996 VDPWR.n1995 130.136
R3867 VDPWR.n2011 VDPWR.n2010 130.136
R3868 VDPWR.n10 VDPWR.t307 130.001
R3869 VDPWR.n11 VDPWR.t225 130.001
R3870 VDPWR.n12 VDPWR.t21 130.001
R3871 VDPWR.n13 VDPWR.t79 130.001
R3872 VDPWR.n2743 VDPWR.t293 130.001
R3873 VDPWR.n370 VDPWR.t178 130.001
R3874 VDPWR.n372 VDPWR.t130 130.001
R3875 VDPWR.n441 VDPWR.t111 130.001
R3876 VDPWR.n418 VDPWR.t100 130.001
R3877 VDPWR.n423 VDPWR.t182 130.001
R3878 VDPWR.n628 VDPWR.t126 130.001
R3879 VDPWR.n626 VDPWR.t134 130.001
R3880 VDPWR.n398 VDPWR.t13 130.001
R3881 VDPWR.n2613 VDPWR.t199 129.47
R3882 VDPWR.t220 VDPWR.t269 128.906
R3883 VDPWR.t37 VDPWR.t118 128.906
R3884 VDPWR.t108 VDPWR.t255 128.906
R3885 VDPWR.t101 VDPWR.t179 128.906
R3886 VDPWR.n466 VDPWR.t128 128.562
R3887 VDPWR.n459 VDPWR.t289 127.754
R3888 VDPWR.n453 VDPWR.t121 127.754
R3889 VDPWR.n1239 VDPWR.t312 125.797
R3890 VDPWR.n1339 VDPWR.t90 125.797
R3891 VDPWR.t235 VDPWR.n35 125.797
R3892 VDPWR.t235 VDPWR.n44 124.352
R3893 VDPWR.t155 VDPWR.t75 122.996
R3894 VDPWR.n676 VDPWR.t147 122.501
R3895 VDPWR.n683 VDPWR.t316 122.501
R3896 VDPWR.n691 VDPWR.t229 122.501
R3897 VDPWR.n585 VDPWR.t223 122.501
R3898 VDPWR.n86 VDPWR.t82 122.501
R3899 VDPWR.n93 VDPWR.t53 122.501
R3900 VDPWR.n450 VDPWR.t239 120.312
R3901 VDPWR.t296 VDPWR.n1994 120.013
R3902 VDPWR.n1894 VDPWR.t297 120.013
R3903 VDPWR.t162 VDPWR.t181 118.919
R3904 VDPWR.t222 VDPWR.t167 118.919
R3905 VDPWR.n2732 VDPWR.n16 117.558
R3906 VDPWR.t92 VDPWR.n18 111.719
R3907 VDPWR.t61 VDPWR.t235 109.287
R3908 VDPWR.t187 VDPWR.t193 108.764
R3909 VDPWR.t175 VDPWR.t145 108.764
R3910 VDPWR.t50 VDPWR.t175 108.764
R3911 VDPWR.n445 VDPWR.t190 107.028
R3912 VDPWR.t158 VDPWR.n444 107.028
R3913 VDPWR.n443 VDPWR.t183 107.028
R3914 VDPWR.n583 VDPWR.t165 107.028
R3915 VDPWR.t14 VDPWR.n2740 106.796
R3916 VDPWR.n2608 VDPWR.n2607 101.718
R3917 VDPWR.n2599 VDPWR.n2596 101.718
R3918 VDPWR.n2586 VDPWR.n2585 101.718
R3919 VDPWR.n2578 VDPWR.n2577 101.718
R3920 VDPWR.t235 VDPWR.n36 47.6173
R3921 VDPWR.t235 VDPWR.n45 47.6173
R3922 VDPWR.n2715 VDPWR.t281 100.18
R3923 VDPWR.n2723 VDPWR.t265 99.9042
R3924 VDPWR.n2726 VDPWR.t103 98.8769
R3925 VDPWR.n2705 VDPWR.n2704 97.8707
R3926 VDPWR.n2697 VDPWR.n2696 97.8707
R3927 VDPWR.n2689 VDPWR.n2688 97.8707
R3928 VDPWR.n2681 VDPWR.n2680 97.8707
R3929 VDPWR.n2655 VDPWR.n2654 97.8707
R3930 VDPWR.n2012 VDPWR.t172 96.8786
R3931 VDPWR.t12 VDPWR.t137 95.1356
R3932 VDPWR.t39 VDPWR.t173 95.1356
R3933 VDPWR.t308 VDPWR.t160 95.1356
R3934 VDPWR.t66 VDPWR.t129 95.1356
R3935 VDPWR.n270 VDPWR.n269 92.2603
R3936 VDPWR.n267 VDPWR.n266 92.2603
R3937 VDPWR.n348 VDPWR.n347 92.2603
R3938 VDPWR.n356 VDPWR.n355 92.2603
R3939 VDPWR.n311 VDPWR.n288 92.2603
R3940 VDPWR.n305 VDPWR.n304 92.2603
R3941 VDPWR.n1401 VDPWR.t89 91.0948
R3942 VDPWR.n2583 VDPWR.n2573 91.069
R3943 VDPWR.n2576 VDPWR.n2573 91.069
R3944 VDPWR.n2580 VDPWR.n2572 91.069
R3945 VDPWR.n2581 VDPWR.n2580 91.069
R3946 VDPWR.n2604 VDPWR.n2603 91.069
R3947 VDPWR.n2603 VDPWR.n2602 91.069
R3948 VDPWR.n2598 VDPWR.n2597 91.069
R3949 VDPWR.t302 VDPWR.t96 86.757
R3950 VDPWR.t49 VDPWR.t72 86.757
R3951 VDPWR.n472 VDPWR.t323 86.0829
R3952 VDPWR.n300 VDPWR.n299 84.306
R3953 VDPWR.n283 VDPWR.n282 84.306
R3954 VDPWR.n336 VDPWR.n256 84.306
R3955 VDPWR.n360 VDPWR.n258 84.306
R3956 VDPWR.n364 VDPWR.n259 84.306
R3957 VDPWR.n337 VDPWR.n257 84.306
R3958 VDPWR.n277 VDPWR.n274 84.306
R3959 VDPWR.n295 VDPWR.n294 84.306
R3960 VDPWR.n2536 VDPWR.n2535 84.306
R3961 VDPWR.n2559 VDPWR.n703 84.306
R3962 VDPWR.n472 VDPWR.t320 82.8829
R3963 VDPWR.n1401 VDPWR.t122 82.4192
R3964 VDPWR.t80 VDPWR.n40 82.4192
R3965 VDPWR.n1340 VDPWR.t60 82.4192
R3966 VDPWR.n2544 VDPWR.n2534 82.4192
R3967 VDPWR.n2671 VDPWR.t1 80.8404
R3968 VDPWR.t1 VDPWR.n2670 80.8404
R3969 VDPWR.n2715 VDPWR.n2714 78.9297
R3970 VDPWR.t281 VDPWR.t230 78.8211
R3971 VDPWR.t230 VDPWR.t300 78.7125
R3972 VDPWR.t300 VDPWR.t114 78.7125
R3973 VDPWR.t265 VDPWR.t169 78.7125
R3974 VDPWR.t131 VDPWR.t74 77.6818
R3975 VDPWR.t28 VDPWR.t17 77.6818
R3976 VDPWR.t291 VDPWR.t192 77.6818
R3977 VDPWR.t192 VDPWR.t189 77.6818
R3978 VDPWR.t189 VDPWR.t155 77.6818
R3979 VDPWR.t75 VDPWR.t154 77.6818
R3980 VDPWR.t154 VDPWR.t163 77.6818
R3981 VDPWR.n2558 VDPWR.n704 76.6354
R3982 VDPWR.n1904 VDPWR.t304 76.6354
R3983 VDPWR.t152 VDPWR.n53 76.6354
R3984 VDPWR.n2012 VDPWR.t142 76.6354
R3985 VDPWR.n74 VDPWR.n60 76.3222
R3986 VDPWR.n2634 VDPWR.n61 76.3222
R3987 VDPWR.n2630 VDPWR.n62 76.3222
R3988 VDPWR.n2412 VDPWR.n63 76.3222
R3989 VDPWR.n1865 VDPWR.n65 76.3222
R3990 VDPWR.n2440 VDPWR.n2439 76.3222
R3991 VDPWR.n2437 VDPWR.n2436 76.3222
R3992 VDPWR.n2432 VDPWR.n1855 76.3222
R3993 VDPWR.n2430 VDPWR.n2429 76.3222
R3994 VDPWR.n2425 VDPWR.n1864 76.3222
R3995 VDPWR.n2423 VDPWR.n2422 76.3222
R3996 VDPWR.n893 VDPWR.n892 76.3222
R3997 VDPWR.n896 VDPWR.n895 76.3222
R3998 VDPWR.n899 VDPWR.n898 76.3222
R3999 VDPWR.n905 VDPWR.n904 76.3222
R4000 VDPWR.n908 VDPWR.n907 76.3222
R4001 VDPWR.n909 VDPWR.n73 76.3222
R4002 VDPWR.n1407 VDPWR.n916 76.3222
R4003 VDPWR.n1411 VDPWR.n917 76.3222
R4004 VDPWR.n1415 VDPWR.n918 76.3222
R4005 VDPWR.n1419 VDPWR.n919 76.3222
R4006 VDPWR.n1423 VDPWR.n920 76.3222
R4007 VDPWR.n1427 VDPWR.n921 76.3222
R4008 VDPWR.n1428 VDPWR.n1234 76.3222
R4009 VDPWR.n1435 VDPWR.n1434 76.3222
R4010 VDPWR.n1436 VDPWR.n1232 76.3222
R4011 VDPWR.n1443 VDPWR.n1442 76.3222
R4012 VDPWR.n1444 VDPWR.n1230 76.3222
R4013 VDPWR.n1451 VDPWR.n1450 76.3222
R4014 VDPWR.n1380 VDPWR.n1351 76.3222
R4015 VDPWR.n1378 VDPWR.n1377 76.3222
R4016 VDPWR.n1373 VDPWR.n1360 76.3222
R4017 VDPWR.n1371 VDPWR.n1370 76.3222
R4018 VDPWR.n1361 VDPWR.n1229 76.3222
R4019 VDPWR.n1453 VDPWR.n1452 76.3222
R4020 VDPWR.n793 VDPWR.n792 76.3222
R4021 VDPWR.n796 VDPWR.n795 76.3222
R4022 VDPWR.n799 VDPWR.n798 76.3222
R4023 VDPWR.n805 VDPWR.n804 76.3222
R4024 VDPWR.n808 VDPWR.n807 76.3222
R4025 VDPWR.n814 VDPWR.n813 76.3222
R4026 VDPWR.n2379 VDPWR.n1889 76.3222
R4027 VDPWR.n2375 VDPWR.n1888 76.3222
R4028 VDPWR.n2371 VDPWR.n1887 76.3222
R4029 VDPWR.n2367 VDPWR.n1886 76.3222
R4030 VDPWR.n2363 VDPWR.n1885 76.3222
R4031 VDPWR.n2359 VDPWR.n1884 76.3222
R4032 VDPWR.n824 VDPWR.n823 76.3222
R4033 VDPWR.n827 VDPWR.n826 76.3222
R4034 VDPWR.n833 VDPWR.n832 76.3222
R4035 VDPWR.n836 VDPWR.n835 76.3222
R4036 VDPWR.n842 VDPWR.n841 76.3222
R4037 VDPWR.n845 VDPWR.n844 76.3222
R4038 VDPWR.n2350 VDPWR.n1871 76.3222
R4039 VDPWR.n2348 VDPWR.n1872 76.3222
R4040 VDPWR.n2345 VDPWR.n1873 76.3222
R4041 VDPWR.n2341 VDPWR.n1874 76.3222
R4042 VDPWR.n2337 VDPWR.n1875 76.3222
R4043 VDPWR.n2333 VDPWR.n1876 76.3222
R4044 VDPWR.n1606 VDPWR.n1097 76.3222
R4045 VDPWR.n1617 VDPWR.n1616 76.3222
R4046 VDPWR.n1618 VDPWR.n1093 76.3222
R4047 VDPWR.n1629 VDPWR.n1628 76.3222
R4048 VDPWR.n1631 VDPWR.n1630 76.3222
R4049 VDPWR.n1089 VDPWR.n883 76.3222
R4050 VDPWR.n2474 VDPWR.n2473 76.3222
R4051 VDPWR.n2469 VDPWR.n829 76.3222
R4052 VDPWR.n2467 VDPWR.n2466 76.3222
R4053 VDPWR.n2462 VDPWR.n838 76.3222
R4054 VDPWR.n2460 VDPWR.n2459 76.3222
R4055 VDPWR.n2455 VDPWR.n847 76.3222
R4056 VDPWR.n1349 VDPWR.n1348 76.3222
R4057 VDPWR.n1355 VDPWR.n1354 76.3222
R4058 VDPWR.n1358 VDPWR.n1357 76.3222
R4059 VDPWR.n1365 VDPWR.n1364 76.3222
R4060 VDPWR.n1366 VDPWR.n1227 76.3222
R4061 VDPWR.n1458 VDPWR.n1457 76.3222
R4062 VDPWR.n2498 VDPWR.n2497 76.3222
R4063 VDPWR.n2495 VDPWR.n2494 76.3222
R4064 VDPWR.n2490 VDPWR.n801 76.3222
R4065 VDPWR.n2488 VDPWR.n2487 76.3222
R4066 VDPWR.n2483 VDPWR.n810 76.3222
R4067 VDPWR.n2481 VDPWR.n2480 76.3222
R4068 VDPWR.n813 VDPWR.n812 76.3222
R4069 VDPWR.n807 VDPWR.n806 76.3222
R4070 VDPWR.n804 VDPWR.n803 76.3222
R4071 VDPWR.n798 VDPWR.n797 76.3222
R4072 VDPWR.n795 VDPWR.n794 76.3222
R4073 VDPWR.n792 VDPWR.n788 76.3222
R4074 VDPWR.n844 VDPWR.n843 76.3222
R4075 VDPWR.n841 VDPWR.n840 76.3222
R4076 VDPWR.n835 VDPWR.n834 76.3222
R4077 VDPWR.n832 VDPWR.n831 76.3222
R4078 VDPWR.n826 VDPWR.n825 76.3222
R4079 VDPWR.n823 VDPWR.n822 76.3222
R4080 VDPWR.n2482 VDPWR.n2481 76.3222
R4081 VDPWR.n810 VDPWR.n802 76.3222
R4082 VDPWR.n2489 VDPWR.n2488 76.3222
R4083 VDPWR.n801 VDPWR.n791 76.3222
R4084 VDPWR.n2496 VDPWR.n2495 76.3222
R4085 VDPWR.n2499 VDPWR.n2498 76.3222
R4086 VDPWR.n847 VDPWR.n839 76.3222
R4087 VDPWR.n2461 VDPWR.n2460 76.3222
R4088 VDPWR.n838 VDPWR.n830 76.3222
R4089 VDPWR.n2468 VDPWR.n2467 76.3222
R4090 VDPWR.n829 VDPWR.n821 76.3222
R4091 VDPWR.n2475 VDPWR.n2474 76.3222
R4092 VDPWR.n1457 VDPWR.n1456 76.3222
R4093 VDPWR.n1367 VDPWR.n1366 76.3222
R4094 VDPWR.n1364 VDPWR.n1363 76.3222
R4095 VDPWR.n1357 VDPWR.n1356 76.3222
R4096 VDPWR.n1354 VDPWR.n1353 76.3222
R4097 VDPWR.n1348 VDPWR.n1347 76.3222
R4098 VDPWR.n1454 VDPWR.n1453 76.3222
R4099 VDPWR.n1362 VDPWR.n1361 76.3222
R4100 VDPWR.n1372 VDPWR.n1371 76.3222
R4101 VDPWR.n1360 VDPWR.n1352 76.3222
R4102 VDPWR.n1379 VDPWR.n1378 76.3222
R4103 VDPWR.n1351 VDPWR.n1343 76.3222
R4104 VDPWR.n1072 VDPWR.n933 76.3222
R4105 VDPWR.n1068 VDPWR.n932 76.3222
R4106 VDPWR.n1064 VDPWR.n931 76.3222
R4107 VDPWR.n1060 VDPWR.n930 76.3222
R4108 VDPWR.n1056 VDPWR.n929 76.3222
R4109 VDPWR.n1687 VDPWR.n1686 76.3222
R4110 VDPWR.n1050 VDPWR.n934 76.3222
R4111 VDPWR.n1049 VDPWR.n937 76.3222
R4112 VDPWR.n971 VDPWR.n970 76.3222
R4113 VDPWR.n974 VDPWR.n973 76.3222
R4114 VDPWR.n986 VDPWR.n985 76.3222
R4115 VDPWR.n990 VDPWR.n989 76.3222
R4116 VDPWR.n1731 VDPWR.n1730 76.3222
R4117 VDPWR.n1728 VDPWR.n1727 76.3222
R4118 VDPWR.n1723 VDPWR.n901 76.3222
R4119 VDPWR.n1721 VDPWR.n1720 76.3222
R4120 VDPWR.n1716 VDPWR.n912 76.3222
R4121 VDPWR.n1714 VDPWR.n1713 76.3222
R4122 VDPWR.n1691 VDPWR.n54 76.3222
R4123 VDPWR.n1695 VDPWR.n55 76.3222
R4124 VDPWR.n1699 VDPWR.n56 76.3222
R4125 VDPWR.n1703 VDPWR.n57 76.3222
R4126 VDPWR.n1707 VDPWR.n58 76.3222
R4127 VDPWR.n1711 VDPWR.n59 76.3222
R4128 VDPWR.n1847 VDPWR.n1846 76.3222
R4129 VDPWR.n1850 VDPWR.n1849 76.3222
R4130 VDPWR.n1853 VDPWR.n1852 76.3222
R4131 VDPWR.n1859 VDPWR.n1858 76.3222
R4132 VDPWR.n1862 VDPWR.n1861 76.3222
R4133 VDPWR.n1868 VDPWR.n1867 76.3222
R4134 VDPWR.n2317 VDPWR.n1879 76.3222
R4135 VDPWR.n2313 VDPWR.n1880 76.3222
R4136 VDPWR.n2309 VDPWR.n1881 76.3222
R4137 VDPWR.n2305 VDPWR.n1882 76.3222
R4138 VDPWR.n2385 VDPWR.n1870 76.3222
R4139 VDPWR.n2407 VDPWR.n66 76.3222
R4140 VDPWR.n2403 VDPWR.n67 76.3222
R4141 VDPWR.n2399 VDPWR.n68 76.3222
R4142 VDPWR.n2395 VDPWR.n69 76.3222
R4143 VDPWR.n2391 VDPWR.n70 76.3222
R4144 VDPWR.n2387 VDPWR.n71 76.3222
R4145 VDPWR.n2390 VDPWR.n71 76.3222
R4146 VDPWR.n2394 VDPWR.n70 76.3222
R4147 VDPWR.n2398 VDPWR.n69 76.3222
R4148 VDPWR.n2402 VDPWR.n68 76.3222
R4149 VDPWR.n2406 VDPWR.n67 76.3222
R4150 VDPWR.n2409 VDPWR.n66 76.3222
R4151 VDPWR.n1708 VDPWR.n59 76.3222
R4152 VDPWR.n1704 VDPWR.n58 76.3222
R4153 VDPWR.n1700 VDPWR.n57 76.3222
R4154 VDPWR.n1696 VDPWR.n56 76.3222
R4155 VDPWR.n1692 VDPWR.n55 76.3222
R4156 VDPWR.n1688 VDPWR.n54 76.3222
R4157 VDPWR.n2362 VDPWR.n1884 76.3222
R4158 VDPWR.n2366 VDPWR.n1885 76.3222
R4159 VDPWR.n2370 VDPWR.n1886 76.3222
R4160 VDPWR.n2374 VDPWR.n1887 76.3222
R4161 VDPWR.n2378 VDPWR.n1888 76.3222
R4162 VDPWR.n2383 VDPWR.n2382 76.3222
R4163 VDPWR.n2330 VDPWR.n1876 76.3222
R4164 VDPWR.n2334 VDPWR.n1875 76.3222
R4165 VDPWR.n2338 VDPWR.n1874 76.3222
R4166 VDPWR.n2342 VDPWR.n1873 76.3222
R4167 VDPWR.n2346 VDPWR.n1872 76.3222
R4168 VDPWR.n2025 VDPWR.n1871 76.3222
R4169 VDPWR.n2386 VDPWR.n2385 76.3222
R4170 VDPWR.n2302 VDPWR.n1882 76.3222
R4171 VDPWR.n2306 VDPWR.n1881 76.3222
R4172 VDPWR.n2310 VDPWR.n1880 76.3222
R4173 VDPWR.n2314 VDPWR.n1879 76.3222
R4174 VDPWR.n2318 VDPWR.n1878 76.3222
R4175 VDPWR.n1450 VDPWR.n1449 76.3222
R4176 VDPWR.n1445 VDPWR.n1444 76.3222
R4177 VDPWR.n1442 VDPWR.n1441 76.3222
R4178 VDPWR.n1437 VDPWR.n1436 76.3222
R4179 VDPWR.n1434 VDPWR.n1433 76.3222
R4180 VDPWR.n1429 VDPWR.n1428 76.3222
R4181 VDPWR.n1051 VDPWR.n1050 76.3222
R4182 VDPWR.n966 VDPWR.n937 76.3222
R4183 VDPWR.n972 VDPWR.n971 76.3222
R4184 VDPWR.n973 VDPWR.n957 76.3222
R4185 VDPWR.n987 VDPWR.n986 76.3222
R4186 VDPWR.n989 VDPWR.n988 76.3222
R4187 VDPWR.n1424 VDPWR.n921 76.3222
R4188 VDPWR.n1420 VDPWR.n920 76.3222
R4189 VDPWR.n1416 VDPWR.n919 76.3222
R4190 VDPWR.n1412 VDPWR.n918 76.3222
R4191 VDPWR.n1408 VDPWR.n917 76.3222
R4192 VDPWR.n1235 VDPWR.n915 76.3222
R4193 VDPWR.n1686 VDPWR.n914 76.3222
R4194 VDPWR.n1059 VDPWR.n929 76.3222
R4195 VDPWR.n1063 VDPWR.n930 76.3222
R4196 VDPWR.n1067 VDPWR.n931 76.3222
R4197 VDPWR.n1071 VDPWR.n932 76.3222
R4198 VDPWR.n1076 VDPWR.n1075 76.3222
R4199 VDPWR.n1660 VDPWR.n1659 76.3222
R4200 VDPWR.n1657 VDPWR.n1656 76.3222
R4201 VDPWR.n1652 VDPWR.n1083 76.3222
R4202 VDPWR.n1650 VDPWR.n1649 76.3222
R4203 VDPWR.n1645 VDPWR.n1086 76.3222
R4204 VDPWR.n1643 VDPWR.n1642 76.3222
R4205 VDPWR.n1611 VDPWR.n1610 76.3222
R4206 VDPWR.n1612 VDPWR.n1095 76.3222
R4207 VDPWR.n1623 VDPWR.n1622 76.3222
R4208 VDPWR.n1624 VDPWR.n1091 76.3222
R4209 VDPWR.n1636 VDPWR.n1635 76.3222
R4210 VDPWR.n1640 VDPWR.n1087 76.3222
R4211 VDPWR.n1131 VDPWR.n1130 76.3222
R4212 VDPWR.n1194 VDPWR.n1193 76.3222
R4213 VDPWR.n1197 VDPWR.n1196 76.3222
R4214 VDPWR.n1206 VDPWR.n1205 76.3222
R4215 VDPWR.n1209 VDPWR.n1208 76.3222
R4216 VDPWR.n1219 VDPWR.n1218 76.3222
R4217 VDPWR.n1684 VDPWR.n1077 76.3222
R4218 VDPWR.n1683 VDPWR.n923 76.3222
R4219 VDPWR.n1679 VDPWR.n924 76.3222
R4220 VDPWR.n1675 VDPWR.n925 76.3222
R4221 VDPWR.n1671 VDPWR.n926 76.3222
R4222 VDPWR.n1667 VDPWR.n927 76.3222
R4223 VDPWR.n1077 VDPWR.n922 76.3222
R4224 VDPWR.n1130 VDPWR.n1128 76.3222
R4225 VDPWR.n1195 VDPWR.n1194 76.3222
R4226 VDPWR.n1196 VDPWR.n1124 76.3222
R4227 VDPWR.n1207 VDPWR.n1206 76.3222
R4228 VDPWR.n1208 VDPWR.n1101 76.3222
R4229 VDPWR.n1220 VDPWR.n1219 76.3222
R4230 VDPWR.n1664 VDPWR.n927 76.3222
R4231 VDPWR.n1668 VDPWR.n926 76.3222
R4232 VDPWR.n1672 VDPWR.n925 76.3222
R4233 VDPWR.n1676 VDPWR.n924 76.3222
R4234 VDPWR.n1680 VDPWR.n923 76.3222
R4235 VDPWR.n1644 VDPWR.n1643 76.3222
R4236 VDPWR.n1086 VDPWR.n1084 76.3222
R4237 VDPWR.n1651 VDPWR.n1650 76.3222
R4238 VDPWR.n1083 VDPWR.n1081 76.3222
R4239 VDPWR.n1658 VDPWR.n1657 76.3222
R4240 VDPWR.n1661 VDPWR.n1660 76.3222
R4241 VDPWR.n1090 VDPWR.n1089 76.3222
R4242 VDPWR.n1632 VDPWR.n1631 76.3222
R4243 VDPWR.n1628 VDPWR.n1627 76.3222
R4244 VDPWR.n1619 VDPWR.n1618 76.3222
R4245 VDPWR.n1616 VDPWR.n1615 76.3222
R4246 VDPWR.n1607 VDPWR.n1606 76.3222
R4247 VDPWR.n1637 VDPWR.n1087 76.3222
R4248 VDPWR.n1635 VDPWR.n1634 76.3222
R4249 VDPWR.n1625 VDPWR.n1624 76.3222
R4250 VDPWR.n1622 VDPWR.n1621 76.3222
R4251 VDPWR.n1613 VDPWR.n1612 76.3222
R4252 VDPWR.n1610 VDPWR.n1609 76.3222
R4253 VDPWR.n910 VDPWR.n909 76.3222
R4254 VDPWR.n907 VDPWR.n906 76.3222
R4255 VDPWR.n904 VDPWR.n903 76.3222
R4256 VDPWR.n898 VDPWR.n897 76.3222
R4257 VDPWR.n895 VDPWR.n894 76.3222
R4258 VDPWR.n892 VDPWR.n887 76.3222
R4259 VDPWR.n1715 VDPWR.n1714 76.3222
R4260 VDPWR.n912 VDPWR.n902 76.3222
R4261 VDPWR.n1722 VDPWR.n1721 76.3222
R4262 VDPWR.n901 VDPWR.n891 76.3222
R4263 VDPWR.n1729 VDPWR.n1728 76.3222
R4264 VDPWR.n1732 VDPWR.n1731 76.3222
R4265 VDPWR.n2300 VDPWR.n1883 76.3222
R4266 VDPWR.n1867 VDPWR.n1866 76.3222
R4267 VDPWR.n1861 VDPWR.n1860 76.3222
R4268 VDPWR.n1858 VDPWR.n1857 76.3222
R4269 VDPWR.n1852 VDPWR.n1851 76.3222
R4270 VDPWR.n1849 VDPWR.n1848 76.3222
R4271 VDPWR.n1846 VDPWR.n1841 76.3222
R4272 VDPWR.n2424 VDPWR.n2423 76.3222
R4273 VDPWR.n1864 VDPWR.n1856 76.3222
R4274 VDPWR.n2431 VDPWR.n2430 76.3222
R4275 VDPWR.n1855 VDPWR.n1845 76.3222
R4276 VDPWR.n2438 VDPWR.n2437 76.3222
R4277 VDPWR.n2441 VDPWR.n2440 76.3222
R4278 VDPWR.n2417 VDPWR.n65 76.3222
R4279 VDPWR.n2414 VDPWR.n63 76.3222
R4280 VDPWR.n2411 VDPWR.n62 76.3222
R4281 VDPWR.n2631 VDPWR.n61 76.3222
R4282 VDPWR.n2635 VDPWR.n60 76.3222
R4283 VDPWR.t8 VDPWR.t273 75.894
R4284 VDPWR.n2100 VDPWR.n2061 74.5978
R4285 VDPWR.n2101 VDPWR.n2100 74.5978
R4286 VDPWR.n1777 VDPWR.n1738 74.5978
R4287 VDPWR.n1778 VDPWR.n1777 74.5978
R4288 VDPWR.n2213 VDPWR.n2142 74.5978
R4289 VDPWR.n2214 VDPWR.n2213 74.5978
R4290 VDPWR.n1956 VDPWR.n1913 74.5978
R4291 VDPWR.n1957 VDPWR.n1956 74.5978
R4292 VDPWR.n1558 VDPWR.n1477 74.5978
R4293 VDPWR.n1559 VDPWR.n1558 74.5978
R4294 VDPWR.n746 VDPWR.n720 74.5978
R4295 VDPWR.n749 VDPWR.n720 74.5978
R4296 VDPWR.n1283 VDPWR.n1253 74.5978
R4297 VDPWR.n1286 VDPWR.n1253 74.5978
R4298 VDPWR.n1027 VDPWR.n1026 74.5978
R4299 VDPWR.n1026 VDPWR.n1025 74.5978
R4300 VDPWR.n1170 VDPWR.n1113 74.5978
R4301 VDPWR.n1167 VDPWR.n1113 74.5978
R4302 VDPWR.t52 VDPWR.t314 71.3518
R4303 VDPWR.n2665 VDPWR.n2664 70.4005
R4304 VDPWR.n2664 VDPWR.n2662 70.4005
R4305 VDPWR.n2297 VDPWR.n2296 69.3109
R4306 VDPWR.n2298 VDPWR.n2297 69.3109
R4307 VDPWR.n1836 VDPWR.n1835 69.3109
R4308 VDPWR.n1837 VDPWR.n1836 69.3109
R4309 VDPWR.n2181 VDPWR.n2180 69.3109
R4310 VDPWR.n2182 VDPWR.n2181 69.3109
R4311 VDPWR.n1924 VDPWR.n1898 69.3109
R4312 VDPWR.n1925 VDPWR.n1924 69.3109
R4313 VDPWR.n1526 VDPWR.n1525 69.3109
R4314 VDPWR.n1527 VDPWR.n1526 69.3109
R4315 VDPWR.n2550 VDPWR.n2549 69.3109
R4316 VDPWR.n2550 VDPWR.n728 69.3109
R4317 VDPWR.n1393 VDPWR.n1392 69.3109
R4318 VDPWR.n1393 VDPWR.n1261 69.3109
R4319 VDPWR.n960 VDPWR.n959 69.3109
R4320 VDPWR.n959 VDPWR.n954 69.3109
R4321 VDPWR.n1215 VDPWR.n1214 69.3109
R4322 VDPWR.n1214 VDPWR.n1104 69.3109
R4323 VDPWR.n2622 VDPWR.n2621 69.0412
R4324 VDPWR.t10 VDPWR.n292 68.7505
R4325 VDPWR.t196 VDPWR.n368 68.7505
R4326 VDPWR.t261 VDPWR.n366 68.7505
R4327 VDPWR.t235 VDPWR.n53 67.9598
R4328 VDPWR.n622 VDPWR.n10 66.69
R4329 VDPWR.n657 VDPWR.n11 66.69
R4330 VDPWR.n663 VDPWR.n12 66.69
R4331 VDPWR.n670 VDPWR.n13 66.69
R4332 VDPWR.n2744 VDPWR.n2743 66.69
R4333 VDPWR.n384 VDPWR.n370 66.69
R4334 VDPWR.n410 VDPWR.n372 66.69
R4335 VDPWR.n441 VDPWR.n440 66.69
R4336 VDPWR.n434 VDPWR.n418 66.69
R4337 VDPWR.n428 VDPWR.n423 66.69
R4338 VDPWR.n2719 VDPWR.n2718 66.5605
R4339 VDPWR.n2720 VDPWR.n2719 66.5605
R4340 VDPWR.n2719 VDPWR.n2642 65.9634
R4341 VDPWR.n692 VDPWR.n691 65.9579
R4342 VDPWR.n677 VDPWR.n676 65.9579
R4343 VDPWR.n684 VDPWR.n683 65.9579
R4344 VDPWR.n2084 VDPWR.t236 65.8183
R4345 VDPWR.n2078 VDPWR.t236 65.8183
R4346 VDPWR.n2076 VDPWR.t236 65.8183
R4347 VDPWR.n2071 VDPWR.t236 65.8183
R4348 VDPWR.n2068 VDPWR.t236 65.8183
R4349 VDPWR.n2091 VDPWR.t236 65.8183
R4350 VDPWR.n2065 VDPWR.t236 65.8183
R4351 VDPWR.n2098 VDPWR.t236 65.8183
R4352 VDPWR.n2106 VDPWR.t236 65.8183
R4353 VDPWR.n2108 VDPWR.t236 65.8183
R4354 VDPWR.n2114 VDPWR.t236 65.8183
R4355 VDPWR.n2116 VDPWR.t236 65.8183
R4356 VDPWR.n1761 VDPWR.t243 65.8183
R4357 VDPWR.n1755 VDPWR.t243 65.8183
R4358 VDPWR.n1753 VDPWR.t243 65.8183
R4359 VDPWR.n1748 VDPWR.t243 65.8183
R4360 VDPWR.n1745 VDPWR.t243 65.8183
R4361 VDPWR.n1768 VDPWR.t243 65.8183
R4362 VDPWR.n1742 VDPWR.t243 65.8183
R4363 VDPWR.n1775 VDPWR.t243 65.8183
R4364 VDPWR.n1783 VDPWR.t243 65.8183
R4365 VDPWR.n1785 VDPWR.t243 65.8183
R4366 VDPWR.n1791 VDPWR.t243 65.8183
R4367 VDPWR.n1793 VDPWR.t243 65.8183
R4368 VDPWR.n2197 VDPWR.t259 65.8183
R4369 VDPWR.n2191 VDPWR.t259 65.8183
R4370 VDPWR.n2189 VDPWR.t259 65.8183
R4371 VDPWR.n2183 VDPWR.t259 65.8183
R4372 VDPWR.n2149 VDPWR.t259 65.8183
R4373 VDPWR.n2204 VDPWR.t259 65.8183
R4374 VDPWR.n2146 VDPWR.t259 65.8183
R4375 VDPWR.n2211 VDPWR.t259 65.8183
R4376 VDPWR.n2219 VDPWR.t259 65.8183
R4377 VDPWR.n2221 VDPWR.t259 65.8183
R4378 VDPWR.n2227 VDPWR.t259 65.8183
R4379 VDPWR.n2229 VDPWR.t259 65.8183
R4380 VDPWR.n1940 VDPWR.t279 65.8183
R4381 VDPWR.n1934 VDPWR.t279 65.8183
R4382 VDPWR.n1932 VDPWR.t279 65.8183
R4383 VDPWR.n1926 VDPWR.t279 65.8183
R4384 VDPWR.n1920 VDPWR.t279 65.8183
R4385 VDPWR.n1947 VDPWR.t279 65.8183
R4386 VDPWR.n1917 VDPWR.t279 65.8183
R4387 VDPWR.n1954 VDPWR.t279 65.8183
R4388 VDPWR.n1962 VDPWR.t279 65.8183
R4389 VDPWR.n1964 VDPWR.t279 65.8183
R4390 VDPWR.n1970 VDPWR.t279 65.8183
R4391 VDPWR.n1972 VDPWR.t279 65.8183
R4392 VDPWR.n1987 VDPWR.t279 65.8183
R4393 VDPWR.n1989 VDPWR.t279 65.8183
R4394 VDPWR.n2002 VDPWR.t279 65.8183
R4395 VDPWR.n2005 VDPWR.t279 65.8183
R4396 VDPWR.n1542 VDPWR.t288 65.8183
R4397 VDPWR.n1536 VDPWR.t288 65.8183
R4398 VDPWR.n1534 VDPWR.t288 65.8183
R4399 VDPWR.n1528 VDPWR.t288 65.8183
R4400 VDPWR.n1484 VDPWR.t288 65.8183
R4401 VDPWR.n1549 VDPWR.t288 65.8183
R4402 VDPWR.n1481 VDPWR.t288 65.8183
R4403 VDPWR.n1556 VDPWR.t288 65.8183
R4404 VDPWR.n1564 VDPWR.t288 65.8183
R4405 VDPWR.n1566 VDPWR.t288 65.8183
R4406 VDPWR.n1572 VDPWR.t288 65.8183
R4407 VDPWR.n1574 VDPWR.t288 65.8183
R4408 VDPWR.n1584 VDPWR.t288 65.8183
R4409 VDPWR.n1587 VDPWR.t288 65.8183
R4410 VDPWR.n1507 VDPWR.t288 65.8183
R4411 VDPWR.n1509 VDPWR.t288 65.8183
R4412 VDPWR.t234 VDPWR.n719 65.8183
R4413 VDPWR.t234 VDPWR.n717 65.8183
R4414 VDPWR.t234 VDPWR.n715 65.8183
R4415 VDPWR.t234 VDPWR.n713 65.8183
R4416 VDPWR.t234 VDPWR.n721 65.8183
R4417 VDPWR.t234 VDPWR.n722 65.8183
R4418 VDPWR.t234 VDPWR.n723 65.8183
R4419 VDPWR.t234 VDPWR.n724 65.8183
R4420 VDPWR.t234 VDPWR.n718 65.8183
R4421 VDPWR.t234 VDPWR.n716 65.8183
R4422 VDPWR.t234 VDPWR.n714 65.8183
R4423 VDPWR.t234 VDPWR.n712 65.8183
R4424 VDPWR.t258 VDPWR.n1252 65.8183
R4425 VDPWR.t258 VDPWR.n1250 65.8183
R4426 VDPWR.t258 VDPWR.n1248 65.8183
R4427 VDPWR.t258 VDPWR.n1246 65.8183
R4428 VDPWR.t258 VDPWR.n1254 65.8183
R4429 VDPWR.t258 VDPWR.n1255 65.8183
R4430 VDPWR.t258 VDPWR.n1256 65.8183
R4431 VDPWR.t258 VDPWR.n1257 65.8183
R4432 VDPWR.t258 VDPWR.n1251 65.8183
R4433 VDPWR.t258 VDPWR.n1249 65.8183
R4434 VDPWR.t258 VDPWR.n1247 65.8183
R4435 VDPWR.t258 VDPWR.n1245 65.8183
R4436 VDPWR.t258 VDPWR.n1258 65.8183
R4437 VDPWR.n1394 VDPWR.t258 65.8183
R4438 VDPWR.t258 VDPWR.n1259 65.8183
R4439 VDPWR.t258 VDPWR.n1260 65.8183
R4440 VDPWR.n2551 VDPWR.t234 65.8183
R4441 VDPWR.t234 VDPWR.n725 65.8183
R4442 VDPWR.t234 VDPWR.n726 65.8183
R4443 VDPWR.t234 VDPWR.n727 65.8183
R4444 VDPWR.n2241 VDPWR.t259 65.8183
R4445 VDPWR.n2244 VDPWR.t259 65.8183
R4446 VDPWR.n2155 VDPWR.t259 65.8183
R4447 VDPWR.n2178 VDPWR.t259 65.8183
R4448 VDPWR.n1006 VDPWR.t242 65.8183
R4449 VDPWR.n1004 VDPWR.t242 65.8183
R4450 VDPWR.n998 VDPWR.t242 65.8183
R4451 VDPWR.n996 VDPWR.t242 65.8183
R4452 VDPWR.n1012 VDPWR.t242 65.8183
R4453 VDPWR.n949 VDPWR.t242 65.8183
R4454 VDPWR.n1019 VDPWR.t242 65.8183
R4455 VDPWR.n946 VDPWR.t242 65.8183
R4456 VDPWR.n1028 VDPWR.t242 65.8183
R4457 VDPWR.n1034 VDPWR.t242 65.8183
R4458 VDPWR.n1036 VDPWR.t242 65.8183
R4459 VDPWR.n1042 VDPWR.t242 65.8183
R4460 VDPWR.n1045 VDPWR.t242 65.8183
R4461 VDPWR.n963 VDPWR.t242 65.8183
R4462 VDPWR.n978 VDPWR.t242 65.8183
R4463 VDPWR.n981 VDPWR.t242 65.8183
R4464 VDPWR.t237 VDPWR.n1112 65.8183
R4465 VDPWR.t237 VDPWR.n1110 65.8183
R4466 VDPWR.t237 VDPWR.n1108 65.8183
R4467 VDPWR.t237 VDPWR.n1106 65.8183
R4468 VDPWR.t237 VDPWR.n1114 65.8183
R4469 VDPWR.t237 VDPWR.n1115 65.8183
R4470 VDPWR.t237 VDPWR.n1116 65.8183
R4471 VDPWR.t237 VDPWR.n1117 65.8183
R4472 VDPWR.t237 VDPWR.n1111 65.8183
R4473 VDPWR.t237 VDPWR.n1109 65.8183
R4474 VDPWR.t237 VDPWR.n1107 65.8183
R4475 VDPWR.t237 VDPWR.n1105 65.8183
R4476 VDPWR.t237 VDPWR.n1118 65.8183
R4477 VDPWR.t237 VDPWR.n1119 65.8183
R4478 VDPWR.t237 VDPWR.n1120 65.8183
R4479 VDPWR.t237 VDPWR.n1213 65.8183
R4480 VDPWR.n1812 VDPWR.t243 65.8183
R4481 VDPWR.n1815 VDPWR.t243 65.8183
R4482 VDPWR.n870 VDPWR.t243 65.8183
R4483 VDPWR.n1833 VDPWR.t243 65.8183
R4484 VDPWR.n2272 VDPWR.t236 65.8183
R4485 VDPWR.n2275 VDPWR.t236 65.8183
R4486 VDPWR.n2049 VDPWR.t236 65.8183
R4487 VDPWR.n2294 VDPWR.t236 65.8183
R4488 VDPWR.n586 VDPWR.n585 65.3889
R4489 VDPWR.n599 VDPWR.n86 65.3889
R4490 VDPWR.n93 VDPWR.n81 65.3889
R4491 VDPWR.t235 VDPWR.n40 62.176
R4492 VDPWR.t235 VDPWR.n32 62.176
R4493 VDPWR.n629 VDPWR.n628 60.8005
R4494 VDPWR.n643 VDPWR.n626 60.8005
R4495 VDPWR.n380 VDPWR.n379 60.8005
R4496 VDPWR.n399 VDPWR.n398 60.8005
R4497 VDPWR.n171 VDPWR.n170 60.8005
R4498 VDPWR.n581 VDPWR.n580 60.8005
R4499 VDPWR.t269 VDPWR.t68 60.1567
R4500 VDPWR.t239 VDPWR.t211 60.1567
R4501 VDPWR.t118 VDPWR.t310 60.1567
R4502 VDPWR.t143 VDPWR.t298 60.1567
R4503 VDPWR.t179 VDPWR.t5 60.1567
R4504 VDPWR.n2643 VDPWR.t301 60.0005
R4505 VDPWR.n2643 VDPWR.t115 60.0005
R4506 VDPWR.n2663 VDPWR.t41 60.0005
R4507 VDPWR.n2663 VDPWR.t313 60.0005
R4508 VDPWR.n2661 VDPWR.t195 60.0005
R4509 VDPWR.n2661 VDPWR.t277 60.0005
R4510 VDPWR.n2659 VDPWR.t249 60.0005
R4511 VDPWR.n2659 VDPWR.t299 60.0005
R4512 VDPWR.n2644 VDPWR.t283 60.0005
R4513 VDPWR.n2644 VDPWR.t231 60.0005
R4514 VDPWR.n2641 VDPWR.t170 60.0005
R4515 VDPWR.n2641 VDPWR.t266 60.0005
R4516 VDPWR.t287 VDPWR.n272 60.0005
R4517 VDPWR.n275 VDPWR.t287 60.0005
R4518 VDPWR.t253 VDPWR.n331 60.0005
R4519 VDPWR.n335 VDPWR.t253 60.0005
R4520 VDPWR.n422 VDPWR.t58 59.46
R4521 VDPWR.t123 VDPWR.n94 59.46
R4522 VDPWR.n2522 VDPWR.t135 59.2841
R4523 VDPWR.n1924 VDPWR.t279 57.8461
R4524 VDPWR.n1526 VDPWR.t288 57.8461
R4525 VDPWR.t258 VDPWR.n1393 57.8461
R4526 VDPWR.t234 VDPWR.n2550 57.8461
R4527 VDPWR.n2181 VDPWR.t259 57.8461
R4528 VDPWR.n959 VDPWR.t242 57.8461
R4529 VDPWR.n1214 VDPWR.t237 57.8461
R4530 VDPWR.n1836 VDPWR.t243 57.8461
R4531 VDPWR.n2297 VDPWR.t236 57.8461
R4532 VDPWR.t235 VDPWR.t205 57.8382
R4533 VDPWR.t235 VDPWR.t207 57.8382
R4534 VDPWR.t114 VDPWR.t235 57.5208
R4535 VDPWR.n2100 VDPWR.t236 55.2026
R4536 VDPWR.n1777 VDPWR.t243 55.2026
R4537 VDPWR.n2213 VDPWR.t259 55.2026
R4538 VDPWR.n1956 VDPWR.t279 55.2026
R4539 VDPWR.n1558 VDPWR.t288 55.2026
R4540 VDPWR.t234 VDPWR.n720 55.2026
R4541 VDPWR.t258 VDPWR.n1253 55.2026
R4542 VDPWR.n1026 VDPWR.t242 55.2026
R4543 VDPWR.t237 VDPWR.n1113 55.2026
R4544 VDPWR.n2724 VDPWR.n2723 54.4934
R4545 VDPWR.n2664 VDPWR.n2652 54.4005
R4546 VDPWR.n2558 VDPWR.n2556 53.5003
R4547 VDPWR.n1994 VDPWR.t304 53.5003
R4548 VDPWR.n1894 VDPWR.t152 53.5003
R4549 VDPWR.t142 VDPWR.n52 53.5003
R4550 VDPWR.n2272 VDPWR.n2271 53.3664
R4551 VDPWR.n2275 VDPWR.n2274 53.3664
R4552 VDPWR.n2054 VDPWR.n2049 53.3664
R4553 VDPWR.n2294 VDPWR.n2293 53.3664
R4554 VDPWR.n2116 VDPWR.n2057 53.3664
R4555 VDPWR.n2115 VDPWR.n2114 53.3664
R4556 VDPWR.n2108 VDPWR.n2059 53.3664
R4557 VDPWR.n2107 VDPWR.n2106 53.3664
R4558 VDPWR.n2098 VDPWR.n2097 53.3664
R4559 VDPWR.n2093 VDPWR.n2065 53.3664
R4560 VDPWR.n2091 VDPWR.n2090 53.3664
R4561 VDPWR.n2086 VDPWR.n2068 53.3664
R4562 VDPWR.n2071 VDPWR.n2033 53.3664
R4563 VDPWR.n2076 VDPWR.n2075 53.3664
R4564 VDPWR.n2079 VDPWR.n2078 53.3664
R4565 VDPWR.n2084 VDPWR.n2083 53.3664
R4566 VDPWR.n2085 VDPWR.n2084 53.3664
R4567 VDPWR.n2078 VDPWR.n2069 53.3664
R4568 VDPWR.n2077 VDPWR.n2076 53.3664
R4569 VDPWR.n2072 VDPWR.n2071 53.3664
R4570 VDPWR.n2068 VDPWR.n2066 53.3664
R4571 VDPWR.n2092 VDPWR.n2091 53.3664
R4572 VDPWR.n2065 VDPWR.n2063 53.3664
R4573 VDPWR.n2099 VDPWR.n2098 53.3664
R4574 VDPWR.n2106 VDPWR.n2105 53.3664
R4575 VDPWR.n2109 VDPWR.n2108 53.3664
R4576 VDPWR.n2114 VDPWR.n2113 53.3664
R4577 VDPWR.n2117 VDPWR.n2116 53.3664
R4578 VDPWR.n1812 VDPWR.n1811 53.3664
R4579 VDPWR.n1815 VDPWR.n1814 53.3664
R4580 VDPWR.n874 VDPWR.n870 53.3664
R4581 VDPWR.n1833 VDPWR.n1832 53.3664
R4582 VDPWR.n1793 VDPWR.n877 53.3664
R4583 VDPWR.n1792 VDPWR.n1791 53.3664
R4584 VDPWR.n1785 VDPWR.n1736 53.3664
R4585 VDPWR.n1784 VDPWR.n1783 53.3664
R4586 VDPWR.n1775 VDPWR.n1774 53.3664
R4587 VDPWR.n1770 VDPWR.n1742 53.3664
R4588 VDPWR.n1768 VDPWR.n1767 53.3664
R4589 VDPWR.n1763 VDPWR.n1745 53.3664
R4590 VDPWR.n1748 VDPWR.n856 53.3664
R4591 VDPWR.n1753 VDPWR.n1752 53.3664
R4592 VDPWR.n1756 VDPWR.n1755 53.3664
R4593 VDPWR.n1761 VDPWR.n1760 53.3664
R4594 VDPWR.n1762 VDPWR.n1761 53.3664
R4595 VDPWR.n1755 VDPWR.n1746 53.3664
R4596 VDPWR.n1754 VDPWR.n1753 53.3664
R4597 VDPWR.n1749 VDPWR.n1748 53.3664
R4598 VDPWR.n1745 VDPWR.n1743 53.3664
R4599 VDPWR.n1769 VDPWR.n1768 53.3664
R4600 VDPWR.n1742 VDPWR.n1740 53.3664
R4601 VDPWR.n1776 VDPWR.n1775 53.3664
R4602 VDPWR.n1783 VDPWR.n1782 53.3664
R4603 VDPWR.n1786 VDPWR.n1785 53.3664
R4604 VDPWR.n1791 VDPWR.n1790 53.3664
R4605 VDPWR.n1794 VDPWR.n1793 53.3664
R4606 VDPWR.n2241 VDPWR.n2240 53.3664
R4607 VDPWR.n2244 VDPWR.n2243 53.3664
R4608 VDPWR.n2155 VDPWR.n2135 53.3664
R4609 VDPWR.n2178 VDPWR.n2177 53.3664
R4610 VDPWR.n2229 VDPWR.n2138 53.3664
R4611 VDPWR.n2228 VDPWR.n2227 53.3664
R4612 VDPWR.n2221 VDPWR.n2140 53.3664
R4613 VDPWR.n2220 VDPWR.n2219 53.3664
R4614 VDPWR.n2211 VDPWR.n2210 53.3664
R4615 VDPWR.n2206 VDPWR.n2146 53.3664
R4616 VDPWR.n2204 VDPWR.n2203 53.3664
R4617 VDPWR.n2199 VDPWR.n2149 53.3664
R4618 VDPWR.n2184 VDPWR.n2183 53.3664
R4619 VDPWR.n2189 VDPWR.n2188 53.3664
R4620 VDPWR.n2192 VDPWR.n2191 53.3664
R4621 VDPWR.n2197 VDPWR.n2196 53.3664
R4622 VDPWR.n2198 VDPWR.n2197 53.3664
R4623 VDPWR.n2191 VDPWR.n2150 53.3664
R4624 VDPWR.n2190 VDPWR.n2189 53.3664
R4625 VDPWR.n2183 VDPWR.n2152 53.3664
R4626 VDPWR.n2149 VDPWR.n2147 53.3664
R4627 VDPWR.n2205 VDPWR.n2204 53.3664
R4628 VDPWR.n2146 VDPWR.n2144 53.3664
R4629 VDPWR.n2212 VDPWR.n2211 53.3664
R4630 VDPWR.n2219 VDPWR.n2218 53.3664
R4631 VDPWR.n2222 VDPWR.n2221 53.3664
R4632 VDPWR.n2227 VDPWR.n2226 53.3664
R4633 VDPWR.n2230 VDPWR.n2229 53.3664
R4634 VDPWR.n1987 VDPWR.n1986 53.3664
R4635 VDPWR.n1990 VDPWR.n1989 53.3664
R4636 VDPWR.n2002 VDPWR.n2001 53.3664
R4637 VDPWR.n2005 VDPWR.n2004 53.3664
R4638 VDPWR.n1972 VDPWR.n1909 53.3664
R4639 VDPWR.n1971 VDPWR.n1970 53.3664
R4640 VDPWR.n1964 VDPWR.n1911 53.3664
R4641 VDPWR.n1963 VDPWR.n1962 53.3664
R4642 VDPWR.n1954 VDPWR.n1953 53.3664
R4643 VDPWR.n1949 VDPWR.n1917 53.3664
R4644 VDPWR.n1947 VDPWR.n1946 53.3664
R4645 VDPWR.n1942 VDPWR.n1920 53.3664
R4646 VDPWR.n1927 VDPWR.n1926 53.3664
R4647 VDPWR.n1932 VDPWR.n1931 53.3664
R4648 VDPWR.n1935 VDPWR.n1934 53.3664
R4649 VDPWR.n1940 VDPWR.n1939 53.3664
R4650 VDPWR.n1941 VDPWR.n1940 53.3664
R4651 VDPWR.n1934 VDPWR.n1921 53.3664
R4652 VDPWR.n1933 VDPWR.n1932 53.3664
R4653 VDPWR.n1926 VDPWR.n1923 53.3664
R4654 VDPWR.n1920 VDPWR.n1918 53.3664
R4655 VDPWR.n1948 VDPWR.n1947 53.3664
R4656 VDPWR.n1917 VDPWR.n1915 53.3664
R4657 VDPWR.n1955 VDPWR.n1954 53.3664
R4658 VDPWR.n1962 VDPWR.n1961 53.3664
R4659 VDPWR.n1965 VDPWR.n1964 53.3664
R4660 VDPWR.n1970 VDPWR.n1969 53.3664
R4661 VDPWR.n1973 VDPWR.n1972 53.3664
R4662 VDPWR.n1988 VDPWR.n1987 53.3664
R4663 VDPWR.n1989 VDPWR.n1901 53.3664
R4664 VDPWR.n2003 VDPWR.n2002 53.3664
R4665 VDPWR.n2006 VDPWR.n2005 53.3664
R4666 VDPWR.n1584 VDPWR.n1583 53.3664
R4667 VDPWR.n1587 VDPWR.n1586 53.3664
R4668 VDPWR.n1507 VDPWR.n1470 53.3664
R4669 VDPWR.n1510 VDPWR.n1509 53.3664
R4670 VDPWR.n1574 VDPWR.n1473 53.3664
R4671 VDPWR.n1573 VDPWR.n1572 53.3664
R4672 VDPWR.n1566 VDPWR.n1475 53.3664
R4673 VDPWR.n1565 VDPWR.n1564 53.3664
R4674 VDPWR.n1556 VDPWR.n1555 53.3664
R4675 VDPWR.n1551 VDPWR.n1481 53.3664
R4676 VDPWR.n1549 VDPWR.n1548 53.3664
R4677 VDPWR.n1544 VDPWR.n1484 53.3664
R4678 VDPWR.n1529 VDPWR.n1528 53.3664
R4679 VDPWR.n1534 VDPWR.n1533 53.3664
R4680 VDPWR.n1537 VDPWR.n1536 53.3664
R4681 VDPWR.n1542 VDPWR.n1541 53.3664
R4682 VDPWR.n1543 VDPWR.n1542 53.3664
R4683 VDPWR.n1536 VDPWR.n1485 53.3664
R4684 VDPWR.n1535 VDPWR.n1534 53.3664
R4685 VDPWR.n1528 VDPWR.n1487 53.3664
R4686 VDPWR.n1484 VDPWR.n1482 53.3664
R4687 VDPWR.n1550 VDPWR.n1549 53.3664
R4688 VDPWR.n1481 VDPWR.n1479 53.3664
R4689 VDPWR.n1557 VDPWR.n1556 53.3664
R4690 VDPWR.n1564 VDPWR.n1563 53.3664
R4691 VDPWR.n1567 VDPWR.n1566 53.3664
R4692 VDPWR.n1572 VDPWR.n1571 53.3664
R4693 VDPWR.n1575 VDPWR.n1574 53.3664
R4694 VDPWR.n1585 VDPWR.n1584 53.3664
R4695 VDPWR.n1588 VDPWR.n1587 53.3664
R4696 VDPWR.n1508 VDPWR.n1507 53.3664
R4697 VDPWR.n1509 VDPWR.n1489 53.3664
R4698 VDPWR.n2552 VDPWR.n2551 53.3664
R4699 VDPWR.n2514 VDPWR.n725 53.3664
R4700 VDPWR.n2517 VDPWR.n726 53.3664
R4701 VDPWR.n2527 VDPWR.n727 53.3664
R4702 VDPWR.n712 VDPWR.n710 53.3664
R4703 VDPWR.n734 VDPWR.n714 53.3664
R4704 VDPWR.n738 VDPWR.n716 53.3664
R4705 VDPWR.n742 VDPWR.n718 53.3664
R4706 VDPWR.n753 VDPWR.n724 53.3664
R4707 VDPWR.n757 VDPWR.n723 53.3664
R4708 VDPWR.n761 VDPWR.n722 53.3664
R4709 VDPWR.n765 VDPWR.n721 53.3664
R4710 VDPWR.n780 VDPWR.n713 53.3664
R4711 VDPWR.n777 VDPWR.n715 53.3664
R4712 VDPWR.n773 VDPWR.n717 53.3664
R4713 VDPWR.n769 VDPWR.n719 53.3664
R4714 VDPWR.n766 VDPWR.n719 53.3664
R4715 VDPWR.n770 VDPWR.n717 53.3664
R4716 VDPWR.n774 VDPWR.n715 53.3664
R4717 VDPWR.n778 VDPWR.n713 53.3664
R4718 VDPWR.n762 VDPWR.n721 53.3664
R4719 VDPWR.n758 VDPWR.n722 53.3664
R4720 VDPWR.n754 VDPWR.n723 53.3664
R4721 VDPWR.n750 VDPWR.n724 53.3664
R4722 VDPWR.n745 VDPWR.n718 53.3664
R4723 VDPWR.n741 VDPWR.n716 53.3664
R4724 VDPWR.n737 VDPWR.n714 53.3664
R4725 VDPWR.n733 VDPWR.n712 53.3664
R4726 VDPWR.n1266 VDPWR.n1258 53.3664
R4727 VDPWR.n1395 VDPWR.n1394 53.3664
R4728 VDPWR.n1327 VDPWR.n1259 53.3664
R4729 VDPWR.n1334 VDPWR.n1260 53.3664
R4730 VDPWR.n1267 VDPWR.n1245 53.3664
R4731 VDPWR.n1271 VDPWR.n1247 53.3664
R4732 VDPWR.n1275 VDPWR.n1249 53.3664
R4733 VDPWR.n1279 VDPWR.n1251 53.3664
R4734 VDPWR.n1290 VDPWR.n1257 53.3664
R4735 VDPWR.n1294 VDPWR.n1256 53.3664
R4736 VDPWR.n1298 VDPWR.n1255 53.3664
R4737 VDPWR.n1302 VDPWR.n1254 53.3664
R4738 VDPWR.n1317 VDPWR.n1246 53.3664
R4739 VDPWR.n1314 VDPWR.n1248 53.3664
R4740 VDPWR.n1310 VDPWR.n1250 53.3664
R4741 VDPWR.n1306 VDPWR.n1252 53.3664
R4742 VDPWR.n1303 VDPWR.n1252 53.3664
R4743 VDPWR.n1307 VDPWR.n1250 53.3664
R4744 VDPWR.n1311 VDPWR.n1248 53.3664
R4745 VDPWR.n1315 VDPWR.n1246 53.3664
R4746 VDPWR.n1299 VDPWR.n1254 53.3664
R4747 VDPWR.n1295 VDPWR.n1255 53.3664
R4748 VDPWR.n1291 VDPWR.n1256 53.3664
R4749 VDPWR.n1287 VDPWR.n1257 53.3664
R4750 VDPWR.n1282 VDPWR.n1251 53.3664
R4751 VDPWR.n1278 VDPWR.n1249 53.3664
R4752 VDPWR.n1274 VDPWR.n1247 53.3664
R4753 VDPWR.n1270 VDPWR.n1245 53.3664
R4754 VDPWR.n1258 VDPWR.n1243 53.3664
R4755 VDPWR.n1394 VDPWR.n1244 53.3664
R4756 VDPWR.n1333 VDPWR.n1259 53.3664
R4757 VDPWR.n1262 VDPWR.n1260 53.3664
R4758 VDPWR.n2551 VDPWR.n711 53.3664
R4759 VDPWR.n2518 VDPWR.n725 53.3664
R4760 VDPWR.n2526 VDPWR.n726 53.3664
R4761 VDPWR.n729 VDPWR.n727 53.3664
R4762 VDPWR.n2242 VDPWR.n2241 53.3664
R4763 VDPWR.n2245 VDPWR.n2244 53.3664
R4764 VDPWR.n2156 VDPWR.n2155 53.3664
R4765 VDPWR.n2179 VDPWR.n2178 53.3664
R4766 VDPWR.n1045 VDPWR.n1044 53.3664
R4767 VDPWR.n963 VDPWR.n939 53.3664
R4768 VDPWR.n978 VDPWR.n977 53.3664
R4769 VDPWR.n981 VDPWR.n980 53.3664
R4770 VDPWR.n1043 VDPWR.n1042 53.3664
R4771 VDPWR.n1036 VDPWR.n940 53.3664
R4772 VDPWR.n1035 VDPWR.n1034 53.3664
R4773 VDPWR.n1028 VDPWR.n942 53.3664
R4774 VDPWR.n1021 VDPWR.n946 53.3664
R4775 VDPWR.n1019 VDPWR.n1018 53.3664
R4776 VDPWR.n1014 VDPWR.n949 53.3664
R4777 VDPWR.n1012 VDPWR.n1011 53.3664
R4778 VDPWR.n996 VDPWR.n995 53.3664
R4779 VDPWR.n999 VDPWR.n998 53.3664
R4780 VDPWR.n1004 VDPWR.n1003 53.3664
R4781 VDPWR.n1007 VDPWR.n1006 53.3664
R4782 VDPWR.n1006 VDPWR.n950 53.3664
R4783 VDPWR.n1005 VDPWR.n1004 53.3664
R4784 VDPWR.n998 VDPWR.n952 53.3664
R4785 VDPWR.n997 VDPWR.n996 53.3664
R4786 VDPWR.n1013 VDPWR.n1012 53.3664
R4787 VDPWR.n949 VDPWR.n947 53.3664
R4788 VDPWR.n1020 VDPWR.n1019 53.3664
R4789 VDPWR.n946 VDPWR.n944 53.3664
R4790 VDPWR.n1029 VDPWR.n1028 53.3664
R4791 VDPWR.n1034 VDPWR.n1033 53.3664
R4792 VDPWR.n1037 VDPWR.n1036 53.3664
R4793 VDPWR.n1042 VDPWR.n1041 53.3664
R4794 VDPWR.n1046 VDPWR.n1045 53.3664
R4795 VDPWR.n964 VDPWR.n963 53.3664
R4796 VDPWR.n979 VDPWR.n978 53.3664
R4797 VDPWR.n982 VDPWR.n981 53.3664
R4798 VDPWR.n1187 VDPWR.n1118 53.3664
R4799 VDPWR.n1189 VDPWR.n1119 53.3664
R4800 VDPWR.n1201 VDPWR.n1120 53.3664
R4801 VDPWR.n1213 VDPWR.n1212 53.3664
R4802 VDPWR.n1186 VDPWR.n1105 53.3664
R4803 VDPWR.n1182 VDPWR.n1107 53.3664
R4804 VDPWR.n1178 VDPWR.n1109 53.3664
R4805 VDPWR.n1174 VDPWR.n1111 53.3664
R4806 VDPWR.n1163 VDPWR.n1117 53.3664
R4807 VDPWR.n1159 VDPWR.n1116 53.3664
R4808 VDPWR.n1155 VDPWR.n1115 53.3664
R4809 VDPWR.n1151 VDPWR.n1114 53.3664
R4810 VDPWR.n1135 VDPWR.n1106 53.3664
R4811 VDPWR.n1139 VDPWR.n1108 53.3664
R4812 VDPWR.n1143 VDPWR.n1110 53.3664
R4813 VDPWR.n1147 VDPWR.n1112 53.3664
R4814 VDPWR.n1150 VDPWR.n1112 53.3664
R4815 VDPWR.n1146 VDPWR.n1110 53.3664
R4816 VDPWR.n1142 VDPWR.n1108 53.3664
R4817 VDPWR.n1138 VDPWR.n1106 53.3664
R4818 VDPWR.n1154 VDPWR.n1114 53.3664
R4819 VDPWR.n1158 VDPWR.n1115 53.3664
R4820 VDPWR.n1162 VDPWR.n1116 53.3664
R4821 VDPWR.n1166 VDPWR.n1117 53.3664
R4822 VDPWR.n1171 VDPWR.n1111 53.3664
R4823 VDPWR.n1175 VDPWR.n1109 53.3664
R4824 VDPWR.n1179 VDPWR.n1107 53.3664
R4825 VDPWR.n1183 VDPWR.n1105 53.3664
R4826 VDPWR.n1190 VDPWR.n1118 53.3664
R4827 VDPWR.n1200 VDPWR.n1119 53.3664
R4828 VDPWR.n1121 VDPWR.n1120 53.3664
R4829 VDPWR.n1213 VDPWR.n1103 53.3664
R4830 VDPWR.n1813 VDPWR.n1812 53.3664
R4831 VDPWR.n1816 VDPWR.n1815 53.3664
R4832 VDPWR.n870 VDPWR.n859 53.3664
R4833 VDPWR.n1834 VDPWR.n1833 53.3664
R4834 VDPWR.n2273 VDPWR.n2272 53.3664
R4835 VDPWR.n2276 VDPWR.n2275 53.3664
R4836 VDPWR.n2049 VDPWR.n2036 53.3664
R4837 VDPWR.n2295 VDPWR.n2294 53.3664
R4838 VDPWR.n123 VDPWR.t25 48.0005
R4839 VDPWR.n123 VDPWR.t151 48.0005
R4840 VDPWR.n125 VDPWR.t191 48.0005
R4841 VDPWR.n125 VDPWR.t227 48.0005
R4842 VDPWR.n138 VDPWR.t159 48.0005
R4843 VDPWR.n138 VDPWR.t35 48.0005
R4844 VDPWR.n116 VDPWR.t138 48.0005
R4845 VDPWR.n116 VDPWR.t174 48.0005
R4846 VDPWR.n114 VDPWR.t309 48.0005
R4847 VDPWR.n114 VDPWR.t67 48.0005
R4848 VDPWR.n108 VDPWR.t57 48.0005
R4849 VDPWR.n108 VDPWR.t65 48.0005
R4850 VDPWR.n163 VDPWR.t86 48.0005
R4851 VDPWR.n163 VDPWR.t295 48.0005
R4852 VDPWR.n189 VDPWR.t166 48.0005
R4853 VDPWR.n189 VDPWR.t48 48.0005
R4854 VDPWR.n195 VDPWR.t19 48.0005
R4855 VDPWR.n195 VDPWR.t77 48.0005
R4856 VDPWR.n204 VDPWR.t106 48.0005
R4857 VDPWR.n204 VDPWR.t46 48.0005
R4858 VDPWR.n205 VDPWR.t4 48.0005
R4859 VDPWR.n205 VDPWR.t95 48.0005
R4860 VDPWR.n210 VDPWR.t221 48.0005
R4861 VDPWR.n210 VDPWR.t69 48.0005
R4862 VDPWR.n215 VDPWR.t233 48.0005
R4863 VDPWR.n215 VDPWR.t213 48.0005
R4864 VDPWR.n218 VDPWR.t215 48.0005
R4865 VDPWR.n218 VDPWR.t217 48.0005
R4866 VDPWR.n222 VDPWR.t38 48.0005
R4867 VDPWR.n222 VDPWR.t311 48.0005
R4868 VDPWR.n227 VDPWR.t23 48.0005
R4869 VDPWR.n227 VDPWR.t33 48.0005
R4870 VDPWR.n230 VDPWR.t55 48.0005
R4871 VDPWR.n230 VDPWR.t109 48.0005
R4872 VDPWR.n238 VDPWR.t93 48.0005
R4873 VDPWR.n238 VDPWR.t194 48.0005
R4874 VDPWR.n242 VDPWR.t188 48.0005
R4875 VDPWR.n242 VDPWR.t104 48.0005
R4876 VDPWR.n499 VDPWR.t176 48.0005
R4877 VDPWR.n499 VDPWR.t51 48.0005
R4878 VDPWR.n234 VDPWR.t102 48.0005
R4879 VDPWR.n234 VDPWR.t6 48.0005
R4880 VDPWR.t122 VDPWR.n38 47.7166
R4881 VDPWR.n1239 VDPWR.t80 47.7166
R4882 VDPWR.t60 VDPWR.n1339 47.7166
R4883 VDPWR.n2545 VDPWR.n2544 47.7166
R4884 VDPWR.t177 VDPWR.t226 47.5681
R4885 VDPWR.t203 VDPWR.t148 47.5681
R4886 VDPWR.t235 VDPWR.n34 47.5454
R4887 VDPWR.t235 VDPWR.n43 47.5454
R4888 VDPWR.n48 VDPWR.n47 47.0176
R4889 VDPWR.t193 VDPWR.n18 44.4949
R4890 VDPWR.n447 VDPWR.t24 44.2319
R4891 VDPWR.n291 VDPWR.t3 42.9693
R4892 VDPWR.n293 VDPWR.t317 42.9693
R4893 VDPWR.n367 VDPWR.t54 42.9693
R4894 VDPWR.n365 VDPWR.t92 42.9693
R4895 VDPWR.t17 VDPWR.t235 42.7252
R4896 VDPWR.n2676 VDPWR.n2675 39.5025
R4897 VDPWR.n2709 VDPWR.n2642 39.4985
R4898 VDPWR.n2669 VDPWR.t8 39.4651
R4899 VDPWR.t89 VDPWR.n1400 39.0409
R4900 VDPWR.n1322 VDPWR.t98 39.0409
R4901 VDPWR.n1388 VDPWR.t302 39.0409
R4902 VDPWR.n1386 VDPWR.t71 39.0409
R4903 VDPWR.n1979 VDPWR.t171 37.595
R4904 VDPWR.n2725 VDPWR.n19 36.8449
R4905 VDPWR.n446 VDPWR.t150 35.6762
R4906 VDPWR.n448 VDPWR.t99 35.6762
R4907 VDPWR.n461 VDPWR.n460 35.6576
R4908 VDPWR.n483 VDPWR.n251 35.6576
R4909 VDPWR.n455 VDPWR.n454 35.6576
R4910 VDPWR.n493 VDPWR.n247 35.6576
R4911 VDPWR.t235 VDPWR.t74 34.9571
R4912 VDPWR.t235 VDPWR.n38 34.7031
R4913 VDPWR.t235 VDPWR.n37 34.4319
R4914 VDPWR.n468 VDPWR.n467 34.3278
R4915 VDPWR.n465 VDPWR.n254 34.3278
R4916 VDPWR.t235 VDPWR.n51 33.9847
R4917 VDPWR.n1981 VDPWR.t49 33.2572
R4918 VDPWR.n1996 VDPWR.t0 33.2572
R4919 VDPWR.t172 VDPWR.n2011 33.2572
R4920 VDPWR.n2588 VDPWR.n2587 33.0535
R4921 VDPWR.n2610 VDPWR.n2609 32.3962
R4922 VDPWR.n2731 VDPWR.n2730 32.257
R4923 VDPWR.n601 VDPWR.n600 32.0005
R4924 VDPWR.n601 VDPWR.n83 32.0005
R4925 VDPWR.n605 VDPWR.n83 32.0005
R4926 VDPWR.n606 VDPWR.n605 32.0005
R4927 VDPWR.n607 VDPWR.n606 32.0005
R4928 VDPWR.n2677 VDPWR.n2676 32.0005
R4929 VDPWR.n2683 VDPWR.n2652 32.0005
R4930 VDPWR.n2684 VDPWR.n2683 32.0005
R4931 VDPWR.n2685 VDPWR.n2684 32.0005
R4932 VDPWR.n2685 VDPWR.n2650 32.0005
R4933 VDPWR.n2691 VDPWR.n2650 32.0005
R4934 VDPWR.n2692 VDPWR.n2691 32.0005
R4935 VDPWR.n2693 VDPWR.n2692 32.0005
R4936 VDPWR.n2693 VDPWR.n2648 32.0005
R4937 VDPWR.n2699 VDPWR.n2648 32.0005
R4938 VDPWR.n2700 VDPWR.n2699 32.0005
R4939 VDPWR.n2701 VDPWR.n2700 32.0005
R4940 VDPWR.n2701 VDPWR.n2646 32.0005
R4941 VDPWR.n2707 VDPWR.n2646 32.0005
R4942 VDPWR.n2708 VDPWR.n2707 32.0005
R4943 VDPWR.n2709 VDPWR.n2708 32.0005
R4944 VDPWR.n656 VDPWR.n655 32.0005
R4945 VDPWR.n657 VDPWR.n656 32.0005
R4946 VDPWR.n661 VDPWR.n620 32.0005
R4947 VDPWR.n662 VDPWR.n661 32.0005
R4948 VDPWR.n664 VDPWR.n662 32.0005
R4949 VDPWR.n668 VDPWR.n618 32.0005
R4950 VDPWR.n669 VDPWR.n668 32.0005
R4951 VDPWR.n674 VDPWR.n616 32.0005
R4952 VDPWR.n675 VDPWR.n674 32.0005
R4953 VDPWR.n677 VDPWR.n675 32.0005
R4954 VDPWR.n681 VDPWR.n614 32.0005
R4955 VDPWR.n682 VDPWR.n681 32.0005
R4956 VDPWR.n688 VDPWR.n612 32.0005
R4957 VDPWR.n689 VDPWR.n688 32.0005
R4958 VDPWR.n651 VDPWR.n622 32.0005
R4959 VDPWR.n649 VDPWR.n624 32.0005
R4960 VDPWR.n644 VDPWR.n643 32.0005
R4961 VDPWR.n638 VDPWR.n629 32.0005
R4962 VDPWR.n636 VDPWR.n631 32.0005
R4963 VDPWR.n2744 VDPWR.n4 32.0005
R4964 VDPWR.n386 VDPWR.n384 32.0005
R4965 VDPWR.n388 VDPWR.n382 32.0005
R4966 VDPWR.n394 VDPWR.n393 32.0005
R4967 VDPWR.n400 VDPWR.n399 32.0005
R4968 VDPWR.n405 VDPWR.n404 32.0005
R4969 VDPWR.n410 VDPWR.n375 32.0005
R4970 VDPWR.n412 VDPWR.n411 32.0005
R4971 VDPWR.n412 VDPWR.n373 32.0005
R4972 VDPWR.n440 VDPWR.n373 32.0005
R4973 VDPWR.n439 VDPWR.n416 32.0005
R4974 VDPWR.n435 VDPWR.n416 32.0005
R4975 VDPWR.n433 VDPWR.n432 32.0005
R4976 VDPWR.n432 VDPWR.n419 32.0005
R4977 VDPWR.n428 VDPWR.n427 32.0005
R4978 VDPWR.n427 VDPWR.n426 32.0005
R4979 VDPWR.n426 VDPWR.n90 32.0005
R4980 VDPWR.n586 VDPWR.n90 32.0005
R4981 VDPWR.n588 VDPWR.n587 32.0005
R4982 VDPWR.n588 VDPWR.n88 32.0005
R4983 VDPWR.n593 VDPWR.n88 32.0005
R4984 VDPWR.n594 VDPWR.n593 32.0005
R4985 VDPWR.n595 VDPWR.n594 32.0005
R4986 VDPWR.n595 VDPWR.n85 32.0005
R4987 VDPWR.n128 VDPWR.n127 32.0005
R4988 VDPWR.n128 VDPWR.n121 32.0005
R4989 VDPWR.n132 VDPWR.n121 32.0005
R4990 VDPWR.n134 VDPWR.n133 32.0005
R4991 VDPWR.n134 VDPWR.n119 32.0005
R4992 VDPWR.n139 VDPWR.n119 32.0005
R4993 VDPWR.n141 VDPWR.n140 32.0005
R4994 VDPWR.n145 VDPWR.n144 32.0005
R4995 VDPWR.n146 VDPWR.n145 32.0005
R4996 VDPWR.n146 VDPWR.n113 32.0005
R4997 VDPWR.n151 VDPWR.n150 32.0005
R4998 VDPWR.n152 VDPWR.n151 32.0005
R4999 VDPWR.n152 VDPWR.n111 32.0005
R5000 VDPWR.n156 VDPWR.n111 32.0005
R5001 VDPWR.n157 VDPWR.n156 32.0005
R5002 VDPWR.n158 VDPWR.n157 32.0005
R5003 VDPWR.n162 VDPWR.n161 32.0005
R5004 VDPWR.n164 VDPWR.n106 32.0005
R5005 VDPWR.n168 VDPWR.n106 32.0005
R5006 VDPWR.n169 VDPWR.n168 32.0005
R5007 VDPWR.n172 VDPWR.n169 32.0005
R5008 VDPWR.n176 VDPWR.n104 32.0005
R5009 VDPWR.n177 VDPWR.n176 32.0005
R5010 VDPWR.n178 VDPWR.n177 32.0005
R5011 VDPWR.n183 VDPWR.n182 32.0005
R5012 VDPWR.n184 VDPWR.n183 32.0005
R5013 VDPWR.n188 VDPWR.n187 32.0005
R5014 VDPWR.n194 VDPWR.n98 32.0005
R5015 VDPWR.n198 VDPWR.n197 32.0005
R5016 VDPWR.n198 VDPWR.n95 32.0005
R5017 VDPWR.n579 VDPWR.n96 32.0005
R5018 VDPWR.n575 VDPWR.n96 32.0005
R5019 VDPWR.n575 VDPWR.n574 32.0005
R5020 VDPWR.n574 VDPWR.n573 32.0005
R5021 VDPWR.n573 VDPWR.n202 32.0005
R5022 VDPWR.n569 VDPWR.n202 32.0005
R5023 VDPWR.n568 VDPWR.n567 32.0005
R5024 VDPWR.n564 VDPWR.n563 32.0005
R5025 VDPWR.n563 VDPWR.n562 32.0005
R5026 VDPWR.n562 VDPWR.n208 32.0005
R5027 VDPWR.n558 VDPWR.n208 32.0005
R5028 VDPWR.n556 VDPWR.n211 32.0005
R5029 VDPWR.n552 VDPWR.n551 32.0005
R5030 VDPWR.n551 VDPWR.n550 32.0005
R5031 VDPWR.n549 VDPWR.n216 32.0005
R5032 VDPWR.n545 VDPWR.n544 32.0005
R5033 VDPWR.n544 VDPWR.n543 32.0005
R5034 VDPWR.n543 VDPWR.n220 32.0005
R5035 VDPWR.n539 VDPWR.n220 32.0005
R5036 VDPWR.n537 VDPWR.n223 32.0005
R5037 VDPWR.n533 VDPWR.n532 32.0005
R5038 VDPWR.n532 VDPWR.n531 32.0005
R5039 VDPWR.n530 VDPWR.n228 32.0005
R5040 VDPWR.n526 VDPWR.n525 32.0005
R5041 VDPWR.n525 VDPWR.n524 32.0005
R5042 VDPWR.n524 VDPWR.n232 32.0005
R5043 VDPWR.n520 VDPWR.n232 32.0005
R5044 VDPWR.n511 VDPWR.n240 32.0005
R5045 VDPWR.n507 VDPWR.n506 32.0005
R5046 VDPWR.n506 VDPWR.n505 32.0005
R5047 VDPWR.n505 VDPWR.n244 32.0005
R5048 VDPWR.n501 VDPWR.n244 32.0005
R5049 VDPWR.n482 VDPWR.n481 32.0005
R5050 VDPWR.n481 VDPWR.n252 32.0005
R5051 VDPWR.n477 VDPWR.n252 32.0005
R5052 VDPWR.n477 VDPWR.n476 32.0005
R5053 VDPWR.n476 VDPWR.n475 32.0005
R5054 VDPWR.n489 VDPWR.n246 32.0005
R5055 VDPWR.n489 VDPWR.n488 32.0005
R5056 VDPWR.n488 VDPWR.n487 32.0005
R5057 VDPWR.n487 VDPWR.n249 32.0005
R5058 VDPWR.n483 VDPWR.n249 32.0005
R5059 VDPWR.n495 VDPWR.n494 32.0005
R5060 VDPWR.n494 VDPWR.n493 32.0005
R5061 VDPWR.n518 VDPWR.n235 32.0005
R5062 VDPWR.n514 VDPWR.n513 32.0005
R5063 VDPWR.n513 VDPWR.n512 32.0005
R5064 VDPWR.n318 VDPWR.n317 32.0005
R5065 VDPWR.n319 VDPWR.n318 32.0005
R5066 VDPWR.n323 VDPWR.n270 32.0005
R5067 VDPWR.n324 VDPWR.n323 32.0005
R5068 VDPWR.n325 VDPWR.n324 32.0005
R5069 VDPWR.n330 VDPWR.n329 32.0005
R5070 VDPWR.n346 VDPWR.n264 32.0005
R5071 VDPWR.n348 VDPWR.n346 32.0005
R5072 VDPWR.n349 VDPWR.n262 32.0005
R5073 VDPWR.n353 VDPWR.n262 32.0005
R5074 VDPWR.n354 VDPWR.n353 32.0005
R5075 VDPWR.n313 VDPWR.n312 32.0005
R5076 VDPWR.n313 VDPWR.n285 32.0005
R5077 VDPWR.n306 VDPWR.n289 32.0005
R5078 VDPWR.n310 VDPWR.n289 32.0005
R5079 VDPWR.n495 VDPWR.n80 29.4625
R5080 VDPWR.n2613 VDPWR.t131 29.131
R5081 VDPWR.n285 VDPWR.n284 29.0291
R5082 VDPWR.n342 VDPWR.n341 29.0291
R5083 VDPWR.t235 VDPWR.t98 28.9193
R5084 VDPWR.t71 VDPWR.t205 28.9193
R5085 VDPWR.t171 VDPWR.t207 28.9193
R5086 VDPWR.t235 VDPWR.t0 28.9193
R5087 VDPWR.t235 VDPWR.n52 28.9193
R5088 VDPWR.n670 VDPWR.n616 28.8005
R5089 VDPWR.n684 VDPWR.n682 28.8005
R5090 VDPWR.n178 VDPWR.n102 28.8005
R5091 VDPWR.n190 VDPWR.n188 28.8005
R5092 VDPWR.n558 VDPWR.n557 28.8005
R5093 VDPWR.n538 VDPWR.n537 28.8005
R5094 VDPWR.n519 VDPWR.n518 28.8005
R5095 VDPWR.n2087 VDPWR.n2067 27.5561
R5096 VDPWR.n1764 VDPWR.n1744 27.5561
R5097 VDPWR.n2200 VDPWR.n2148 27.5561
R5098 VDPWR.n1943 VDPWR.n1919 27.5561
R5099 VDPWR.n1545 VDPWR.n1483 27.5561
R5100 VDPWR.n767 VDPWR.n764 27.5561
R5101 VDPWR.n1304 VDPWR.n1301 27.5561
R5102 VDPWR.n1010 VDPWR.n1009 27.5561
R5103 VDPWR.n1152 VDPWR.n1149 27.5561
R5104 VDPWR.n2717 VDPWR.n2716 27.2005
R5105 VDPWR.n2722 VDPWR.n2721 27.2005
R5106 VDPWR.n2103 VDPWR.n2102 26.6672
R5107 VDPWR.n1780 VDPWR.n1779 26.6672
R5108 VDPWR.n2216 VDPWR.n2215 26.6672
R5109 VDPWR.n1959 VDPWR.n1958 26.6672
R5110 VDPWR.n1561 VDPWR.n1560 26.6672
R5111 VDPWR.n748 VDPWR.n747 26.6672
R5112 VDPWR.n1285 VDPWR.n1284 26.6672
R5113 VDPWR.n1024 VDPWR.n943 26.6672
R5114 VDPWR.n1169 VDPWR.n1168 26.6672
R5115 VDPWR.t116 VDPWR.t232 25.7817
R5116 VDPWR.t285 VDPWR.t214 25.7817
R5117 VDPWR.t251 VDPWR.t22 25.7817
R5118 VDPWR.n600 VDPWR.n599 25.6005
R5119 VDPWR.n2660 VDPWR.n2658 25.6005
R5120 VDPWR.n2667 VDPWR.n2666 25.6005
R5121 VDPWR.n692 VDPWR.n689 25.6005
R5122 VDPWR.n651 VDPWR.n650 25.6005
R5123 VDPWR.n645 VDPWR.n624 25.6005
R5124 VDPWR.n650 VDPWR.n649 25.6005
R5125 VDPWR.n645 VDPWR.n644 25.6005
R5126 VDPWR.n638 VDPWR.n637 25.6005
R5127 VDPWR.n632 VDPWR.n631 25.6005
R5128 VDPWR.n637 VDPWR.n636 25.6005
R5129 VDPWR.n632 VDPWR.n4 25.6005
R5130 VDPWR.n387 VDPWR.n386 25.6005
R5131 VDPWR.n388 VDPWR.n387 25.6005
R5132 VDPWR.n392 VDPWR.n382 25.6005
R5133 VDPWR.n393 VDPWR.n392 25.6005
R5134 VDPWR.n400 VDPWR.n377 25.6005
R5135 VDPWR.n404 VDPWR.n377 25.6005
R5136 VDPWR.n406 VDPWR.n405 25.6005
R5137 VDPWR.n406 VDPWR.n375 25.6005
R5138 VDPWR.n599 VDPWR.n85 25.6005
R5139 VDPWR.n475 VDPWR.n254 25.6005
R5140 VDPWR.n342 VDPWR.n330 25.6005
R5141 VDPWR.n306 VDPWR.n305 25.6005
R5142 VDPWR.n311 VDPWR.n310 25.6005
R5143 VDPWR.n2609 VDPWR.n2595 25.3679
R5144 VDPWR.n2713 VDPWR.n2712 24.8279
R5145 VDPWR.t145 VDPWR.n451 24.7196
R5146 VDPWR.n2704 VDPWR.t186 24.0005
R5147 VDPWR.n2704 VDPWR.t274 24.0005
R5148 VDPWR.n2696 VDPWR.t139 24.0005
R5149 VDPWR.n2696 VDPWR.t305 24.0005
R5150 VDPWR.n2688 VDPWR.t97 24.0005
R5151 VDPWR.n2688 VDPWR.t2 24.0005
R5152 VDPWR.n2680 VDPWR.t157 24.0005
R5153 VDPWR.n2680 VDPWR.t91 24.0005
R5154 VDPWR.n2654 VDPWR.t246 24.0005
R5155 VDPWR.n2654 VDPWR.t185 24.0005
R5156 VDPWR.t47 VDPWR.t81 23.7843
R5157 VDPWR.n498 VDPWR.n497 23.1805
R5158 VDPWR.n2674 VDPWR.n2673 22.4005
R5159 VDPWR.n670 VDPWR.n669 22.4005
R5160 VDPWR.n684 VDPWR.n612 22.4005
R5161 VDPWR.n127 VDPWR.n126 22.4005
R5162 VDPWR.n182 VDPWR.n102 22.4005
R5163 VDPWR.n190 VDPWR.n98 22.4005
R5164 VDPWR.n557 VDPWR.n556 22.4005
R5165 VDPWR.n539 VDPWR.n538 22.4005
R5166 VDPWR.n520 VDPWR.n519 22.4005
R5167 VDPWR.n501 VDPWR.n500 22.4005
R5168 VDPWR.t169 VDPWR.t235 21.1922
R5169 VDPWR.n358 VDPWR.n357 20.9665
R5170 VDPWR.n303 VDPWR.n302 19.3316
R5171 VDPWR.n607 VDPWR.n81 19.2005
R5172 VDPWR.n2677 VDPWR.n2652 19.2005
R5173 VDPWR.n655 VDPWR.n622 19.2005
R5174 VDPWR.n657 VDPWR.n620 19.2005
R5175 VDPWR.n677 VDPWR.n614 19.2005
R5176 VDPWR.n642 VDPWR.n629 19.2005
R5177 VDPWR.n643 VDPWR.n642 19.2005
R5178 VDPWR.n399 VDPWR.n397 19.2005
R5179 VDPWR.n411 VDPWR.n410 19.2005
R5180 VDPWR.n440 VDPWR.n439 19.2005
R5181 VDPWR.n428 VDPWR.n419 19.2005
R5182 VDPWR.n587 VDPWR.n586 19.2005
R5183 VDPWR.n133 VDPWR.n132 19.2005
R5184 VDPWR.n140 VDPWR.n139 19.2005
R5185 VDPWR.n150 VDPWR.n113 19.2005
R5186 VDPWR.n164 VDPWR.n162 19.2005
R5187 VDPWR.n569 VDPWR.n568 19.2005
R5188 VDPWR.n550 VDPWR.n549 19.2005
R5189 VDPWR.n531 VDPWR.n530 19.2005
R5190 VDPWR.n512 VDPWR.n511 19.2005
R5191 VDPWR.n325 VDPWR.n267 19.2005
R5192 VDPWR.n329 VDPWR.n267 19.2005
R5193 VDPWR.n1430 VDPWR.n1426 17.5843
R5194 VDPWR.n1689 VDPWR.n913 17.5843
R5195 VDPWR.n1663 VDPWR.n1662 17.5843
R5196 VDPWR.n2360 VDPWR.n2017 17.0672
R5197 VDPWR.n2329 VDPWR.n2328 17.0672
R5198 VDPWR.n2388 VDPWR.n1869 17.0672
R5199 VDPWR.n2628 VDPWR.n2627 16.9605
R5200 VDPWR.n1840 VDPWR.n846 16.7235
R5201 VDPWR.n1604 VDPWR.n1603 16.7235
R5202 VDPWR.n2478 VDPWR.n2477 16.7235
R5203 VDPWR.n886 VDPWR.n882 16.7235
R5204 VDPWR.n610 VDPWR.n80 16.0525
R5205 VDPWR.n2299 VDPWR.n2032 16.0005
R5206 VDPWR.n2073 VDPWR.n2032 16.0005
R5207 VDPWR.n2074 VDPWR.n2073 16.0005
R5208 VDPWR.n2074 VDPWR.n2070 16.0005
R5209 VDPWR.n2080 VDPWR.n2070 16.0005
R5210 VDPWR.n2081 VDPWR.n2080 16.0005
R5211 VDPWR.n2082 VDPWR.n2081 16.0005
R5212 VDPWR.n2082 VDPWR.n2067 16.0005
R5213 VDPWR.n2102 VDPWR.n2062 16.0005
R5214 VDPWR.n2096 VDPWR.n2062 16.0005
R5215 VDPWR.n2096 VDPWR.n2095 16.0005
R5216 VDPWR.n2095 VDPWR.n2094 16.0005
R5217 VDPWR.n2094 VDPWR.n2064 16.0005
R5218 VDPWR.n2089 VDPWR.n2064 16.0005
R5219 VDPWR.n2089 VDPWR.n2088 16.0005
R5220 VDPWR.n2088 VDPWR.n2087 16.0005
R5221 VDPWR.n2119 VDPWR.n2118 16.0005
R5222 VDPWR.n2118 VDPWR.n2058 16.0005
R5223 VDPWR.n2112 VDPWR.n2058 16.0005
R5224 VDPWR.n2112 VDPWR.n2111 16.0005
R5225 VDPWR.n2111 VDPWR.n2110 16.0005
R5226 VDPWR.n2110 VDPWR.n2060 16.0005
R5227 VDPWR.n2104 VDPWR.n2060 16.0005
R5228 VDPWR.n2104 VDPWR.n2103 16.0005
R5229 VDPWR.n1838 VDPWR.n855 16.0005
R5230 VDPWR.n1750 VDPWR.n855 16.0005
R5231 VDPWR.n1751 VDPWR.n1750 16.0005
R5232 VDPWR.n1751 VDPWR.n1747 16.0005
R5233 VDPWR.n1757 VDPWR.n1747 16.0005
R5234 VDPWR.n1758 VDPWR.n1757 16.0005
R5235 VDPWR.n1759 VDPWR.n1758 16.0005
R5236 VDPWR.n1759 VDPWR.n1744 16.0005
R5237 VDPWR.n1779 VDPWR.n1739 16.0005
R5238 VDPWR.n1773 VDPWR.n1739 16.0005
R5239 VDPWR.n1773 VDPWR.n1772 16.0005
R5240 VDPWR.n1772 VDPWR.n1771 16.0005
R5241 VDPWR.n1771 VDPWR.n1741 16.0005
R5242 VDPWR.n1766 VDPWR.n1741 16.0005
R5243 VDPWR.n1766 VDPWR.n1765 16.0005
R5244 VDPWR.n1765 VDPWR.n1764 16.0005
R5245 VDPWR.n1796 VDPWR.n1795 16.0005
R5246 VDPWR.n1795 VDPWR.n1735 16.0005
R5247 VDPWR.n1789 VDPWR.n1735 16.0005
R5248 VDPWR.n1789 VDPWR.n1788 16.0005
R5249 VDPWR.n1788 VDPWR.n1787 16.0005
R5250 VDPWR.n1787 VDPWR.n1737 16.0005
R5251 VDPWR.n1781 VDPWR.n1737 16.0005
R5252 VDPWR.n1781 VDPWR.n1780 16.0005
R5253 VDPWR.n2185 VDPWR.n2024 16.0005
R5254 VDPWR.n2186 VDPWR.n2185 16.0005
R5255 VDPWR.n2187 VDPWR.n2186 16.0005
R5256 VDPWR.n2187 VDPWR.n2151 16.0005
R5257 VDPWR.n2193 VDPWR.n2151 16.0005
R5258 VDPWR.n2194 VDPWR.n2193 16.0005
R5259 VDPWR.n2195 VDPWR.n2194 16.0005
R5260 VDPWR.n2195 VDPWR.n2148 16.0005
R5261 VDPWR.n2215 VDPWR.n2143 16.0005
R5262 VDPWR.n2209 VDPWR.n2143 16.0005
R5263 VDPWR.n2209 VDPWR.n2208 16.0005
R5264 VDPWR.n2208 VDPWR.n2207 16.0005
R5265 VDPWR.n2207 VDPWR.n2145 16.0005
R5266 VDPWR.n2202 VDPWR.n2145 16.0005
R5267 VDPWR.n2202 VDPWR.n2201 16.0005
R5268 VDPWR.n2201 VDPWR.n2200 16.0005
R5269 VDPWR.n2232 VDPWR.n2231 16.0005
R5270 VDPWR.n2231 VDPWR.n2139 16.0005
R5271 VDPWR.n2225 VDPWR.n2139 16.0005
R5272 VDPWR.n2225 VDPWR.n2224 16.0005
R5273 VDPWR.n2224 VDPWR.n2223 16.0005
R5274 VDPWR.n2223 VDPWR.n2141 16.0005
R5275 VDPWR.n2217 VDPWR.n2141 16.0005
R5276 VDPWR.n2217 VDPWR.n2216 16.0005
R5277 VDPWR.n1928 VDPWR.n1891 16.0005
R5278 VDPWR.n1929 VDPWR.n1928 16.0005
R5279 VDPWR.n1930 VDPWR.n1929 16.0005
R5280 VDPWR.n1930 VDPWR.n1922 16.0005
R5281 VDPWR.n1936 VDPWR.n1922 16.0005
R5282 VDPWR.n1937 VDPWR.n1936 16.0005
R5283 VDPWR.n1938 VDPWR.n1937 16.0005
R5284 VDPWR.n1938 VDPWR.n1919 16.0005
R5285 VDPWR.n1958 VDPWR.n1914 16.0005
R5286 VDPWR.n1952 VDPWR.n1914 16.0005
R5287 VDPWR.n1952 VDPWR.n1951 16.0005
R5288 VDPWR.n1951 VDPWR.n1950 16.0005
R5289 VDPWR.n1950 VDPWR.n1916 16.0005
R5290 VDPWR.n1945 VDPWR.n1916 16.0005
R5291 VDPWR.n1945 VDPWR.n1944 16.0005
R5292 VDPWR.n1944 VDPWR.n1943 16.0005
R5293 VDPWR.n1975 VDPWR.n1974 16.0005
R5294 VDPWR.n1974 VDPWR.n1910 16.0005
R5295 VDPWR.n1968 VDPWR.n1910 16.0005
R5296 VDPWR.n1968 VDPWR.n1967 16.0005
R5297 VDPWR.n1967 VDPWR.n1966 16.0005
R5298 VDPWR.n1966 VDPWR.n1912 16.0005
R5299 VDPWR.n1960 VDPWR.n1912 16.0005
R5300 VDPWR.n1960 VDPWR.n1959 16.0005
R5301 VDPWR.n1530 VDPWR.n1488 16.0005
R5302 VDPWR.n1531 VDPWR.n1530 16.0005
R5303 VDPWR.n1532 VDPWR.n1531 16.0005
R5304 VDPWR.n1532 VDPWR.n1486 16.0005
R5305 VDPWR.n1538 VDPWR.n1486 16.0005
R5306 VDPWR.n1539 VDPWR.n1538 16.0005
R5307 VDPWR.n1540 VDPWR.n1539 16.0005
R5308 VDPWR.n1540 VDPWR.n1483 16.0005
R5309 VDPWR.n1560 VDPWR.n1478 16.0005
R5310 VDPWR.n1554 VDPWR.n1478 16.0005
R5311 VDPWR.n1554 VDPWR.n1553 16.0005
R5312 VDPWR.n1553 VDPWR.n1552 16.0005
R5313 VDPWR.n1552 VDPWR.n1480 16.0005
R5314 VDPWR.n1547 VDPWR.n1480 16.0005
R5315 VDPWR.n1547 VDPWR.n1546 16.0005
R5316 VDPWR.n1546 VDPWR.n1545 16.0005
R5317 VDPWR.n1577 VDPWR.n1576 16.0005
R5318 VDPWR.n1576 VDPWR.n1474 16.0005
R5319 VDPWR.n1570 VDPWR.n1474 16.0005
R5320 VDPWR.n1570 VDPWR.n1569 16.0005
R5321 VDPWR.n1569 VDPWR.n1568 16.0005
R5322 VDPWR.n1568 VDPWR.n1476 16.0005
R5323 VDPWR.n1562 VDPWR.n1476 16.0005
R5324 VDPWR.n1562 VDPWR.n1561 16.0005
R5325 VDPWR.n782 VDPWR.n781 16.0005
R5326 VDPWR.n781 VDPWR.n779 16.0005
R5327 VDPWR.n779 VDPWR.n776 16.0005
R5328 VDPWR.n776 VDPWR.n775 16.0005
R5329 VDPWR.n775 VDPWR.n772 16.0005
R5330 VDPWR.n772 VDPWR.n771 16.0005
R5331 VDPWR.n771 VDPWR.n768 16.0005
R5332 VDPWR.n768 VDPWR.n767 16.0005
R5333 VDPWR.n751 VDPWR.n748 16.0005
R5334 VDPWR.n752 VDPWR.n751 16.0005
R5335 VDPWR.n755 VDPWR.n752 16.0005
R5336 VDPWR.n756 VDPWR.n755 16.0005
R5337 VDPWR.n759 VDPWR.n756 16.0005
R5338 VDPWR.n760 VDPWR.n759 16.0005
R5339 VDPWR.n763 VDPWR.n760 16.0005
R5340 VDPWR.n764 VDPWR.n763 16.0005
R5341 VDPWR.n732 VDPWR.n731 16.0005
R5342 VDPWR.n735 VDPWR.n732 16.0005
R5343 VDPWR.n736 VDPWR.n735 16.0005
R5344 VDPWR.n739 VDPWR.n736 16.0005
R5345 VDPWR.n740 VDPWR.n739 16.0005
R5346 VDPWR.n743 VDPWR.n740 16.0005
R5347 VDPWR.n744 VDPWR.n743 16.0005
R5348 VDPWR.n747 VDPWR.n744 16.0005
R5349 VDPWR.n1319 VDPWR.n1318 16.0005
R5350 VDPWR.n1318 VDPWR.n1316 16.0005
R5351 VDPWR.n1316 VDPWR.n1313 16.0005
R5352 VDPWR.n1313 VDPWR.n1312 16.0005
R5353 VDPWR.n1312 VDPWR.n1309 16.0005
R5354 VDPWR.n1309 VDPWR.n1308 16.0005
R5355 VDPWR.n1308 VDPWR.n1305 16.0005
R5356 VDPWR.n1305 VDPWR.n1304 16.0005
R5357 VDPWR.n1288 VDPWR.n1285 16.0005
R5358 VDPWR.n1289 VDPWR.n1288 16.0005
R5359 VDPWR.n1292 VDPWR.n1289 16.0005
R5360 VDPWR.n1293 VDPWR.n1292 16.0005
R5361 VDPWR.n1296 VDPWR.n1293 16.0005
R5362 VDPWR.n1297 VDPWR.n1296 16.0005
R5363 VDPWR.n1300 VDPWR.n1297 16.0005
R5364 VDPWR.n1301 VDPWR.n1300 16.0005
R5365 VDPWR.n1269 VDPWR.n1268 16.0005
R5366 VDPWR.n1272 VDPWR.n1269 16.0005
R5367 VDPWR.n1273 VDPWR.n1272 16.0005
R5368 VDPWR.n1276 VDPWR.n1273 16.0005
R5369 VDPWR.n1277 VDPWR.n1276 16.0005
R5370 VDPWR.n1280 VDPWR.n1277 16.0005
R5371 VDPWR.n1281 VDPWR.n1280 16.0005
R5372 VDPWR.n1284 VDPWR.n1281 16.0005
R5373 VDPWR.n994 VDPWR.n993 16.0005
R5374 VDPWR.n994 VDPWR.n953 16.0005
R5375 VDPWR.n1000 VDPWR.n953 16.0005
R5376 VDPWR.n1001 VDPWR.n1000 16.0005
R5377 VDPWR.n1002 VDPWR.n1001 16.0005
R5378 VDPWR.n1002 VDPWR.n951 16.0005
R5379 VDPWR.n1008 VDPWR.n951 16.0005
R5380 VDPWR.n1009 VDPWR.n1008 16.0005
R5381 VDPWR.n1024 VDPWR.n1023 16.0005
R5382 VDPWR.n1023 VDPWR.n1022 16.0005
R5383 VDPWR.n1022 VDPWR.n945 16.0005
R5384 VDPWR.n1017 VDPWR.n945 16.0005
R5385 VDPWR.n1017 VDPWR.n1016 16.0005
R5386 VDPWR.n1016 VDPWR.n1015 16.0005
R5387 VDPWR.n1015 VDPWR.n948 16.0005
R5388 VDPWR.n1010 VDPWR.n948 16.0005
R5389 VDPWR.n1040 VDPWR.n935 16.0005
R5390 VDPWR.n1040 VDPWR.n1039 16.0005
R5391 VDPWR.n1039 VDPWR.n1038 16.0005
R5392 VDPWR.n1038 VDPWR.n941 16.0005
R5393 VDPWR.n1032 VDPWR.n941 16.0005
R5394 VDPWR.n1032 VDPWR.n1031 16.0005
R5395 VDPWR.n1031 VDPWR.n1030 16.0005
R5396 VDPWR.n1030 VDPWR.n943 16.0005
R5397 VDPWR.n397 VDPWR.n380 16.0005
R5398 VDPWR.n197 VDPWR.n196 16.0005
R5399 VDPWR.n213 VDPWR.n211 16.0005
R5400 VDPWR.n225 VDPWR.n223 16.0005
R5401 VDPWR.n237 VDPWR.n235 16.0005
R5402 VDPWR.n1136 VDPWR.n1134 16.0005
R5403 VDPWR.n1137 VDPWR.n1136 16.0005
R5404 VDPWR.n1140 VDPWR.n1137 16.0005
R5405 VDPWR.n1141 VDPWR.n1140 16.0005
R5406 VDPWR.n1144 VDPWR.n1141 16.0005
R5407 VDPWR.n1145 VDPWR.n1144 16.0005
R5408 VDPWR.n1148 VDPWR.n1145 16.0005
R5409 VDPWR.n1149 VDPWR.n1148 16.0005
R5410 VDPWR.n1168 VDPWR.n1165 16.0005
R5411 VDPWR.n1165 VDPWR.n1164 16.0005
R5412 VDPWR.n1164 VDPWR.n1161 16.0005
R5413 VDPWR.n1161 VDPWR.n1160 16.0005
R5414 VDPWR.n1160 VDPWR.n1157 16.0005
R5415 VDPWR.n1157 VDPWR.n1156 16.0005
R5416 VDPWR.n1156 VDPWR.n1153 16.0005
R5417 VDPWR.n1153 VDPWR.n1152 16.0005
R5418 VDPWR.n1185 VDPWR.n1184 16.0005
R5419 VDPWR.n1184 VDPWR.n1181 16.0005
R5420 VDPWR.n1181 VDPWR.n1180 16.0005
R5421 VDPWR.n1180 VDPWR.n1177 16.0005
R5422 VDPWR.n1177 VDPWR.n1176 16.0005
R5423 VDPWR.n1176 VDPWR.n1173 16.0005
R5424 VDPWR.n1173 VDPWR.n1172 16.0005
R5425 VDPWR.n1172 VDPWR.n1169 16.0005
R5426 VDPWR.n302 VDPWR.n301 15.6449
R5427 VDPWR.n359 VDPWR.n358 15.6449
R5428 VDPWR.n2640 VDPWR.n72 15.105
R5429 VDPWR.n269 VDPWR.t241 15.0005
R5430 VDPWR.n269 VDPWR.t119 15.0005
R5431 VDPWR.n266 VDPWR.t197 15.0005
R5432 VDPWR.n266 VDPWR.t252 15.0005
R5433 VDPWR.n347 VDPWR.t257 15.0005
R5434 VDPWR.n347 VDPWR.t144 15.0005
R5435 VDPWR.n355 VDPWR.t180 15.0005
R5436 VDPWR.n355 VDPWR.t262 15.0005
R5437 VDPWR.n288 VDPWR.t117 15.0005
R5438 VDPWR.n288 VDPWR.t286 15.0005
R5439 VDPWR.n304 VDPWR.t271 15.0005
R5440 VDPWR.n304 VDPWR.t11 15.0005
R5441 VDPWR.n2718 VDPWR.n2717 14.0805
R5442 VDPWR.n2721 VDPWR.n2720 14.0805
R5443 VDPWR.n2746 VDPWR.n2 13.0271
R5444 VDPWR.n2561 VDPWR.n702 12.8005
R5445 VDPWR.n2561 VDPWR.n2560 12.8005
R5446 VDPWR.n2542 VDPWR.n2541 12.8005
R5447 VDPWR.n2541 VDPWR.n2538 12.8005
R5448 VDPWR.n664 VDPWR.n663 12.8005
R5449 VDPWR.n144 VDPWR.n117 12.8005
R5450 VDPWR.n158 VDPWR.n109 12.8005
R5451 VDPWR.n184 VDPWR.n100 12.8005
R5452 VDPWR.n580 VDPWR.n95 12.8005
R5453 VDPWR.n564 VDPWR.n206 12.8005
R5454 VDPWR.n545 VDPWR.n219 12.8005
R5455 VDPWR.n526 VDPWR.n231 12.8005
R5456 VDPWR.n507 VDPWR.n243 12.8005
R5457 VDPWR.n483 VDPWR.n482 12.8005
R5458 VDPWR.n493 VDPWR.n246 12.8005
R5459 VDPWR.n342 VDPWR.n264 12.8005
R5460 VDPWR.n356 VDPWR.n354 12.8005
R5461 VDPWR.n312 VDPWR.n311 12.8005
R5462 VDPWR.n2627 VDPWR.n78 12.8005
R5463 VDPWR.n2623 VDPWR.n78 12.8005
R5464 VDPWR.n2746 VDPWR.n2745 11.9273
R5465 VDPWR.t56 VDPWR.n442 11.8924
R5466 VDPWR.n448 VDPWR.t85 11.8924
R5467 VDPWR.n421 VDPWR.t294 11.8924
R5468 VDPWR.n2380 VDPWR.n2377 11.6369
R5469 VDPWR.n2377 VDPWR.n2376 11.6369
R5470 VDPWR.n2376 VDPWR.n2373 11.6369
R5471 VDPWR.n2373 VDPWR.n2372 11.6369
R5472 VDPWR.n2372 VDPWR.n2369 11.6369
R5473 VDPWR.n2369 VDPWR.n2368 11.6369
R5474 VDPWR.n2368 VDPWR.n2365 11.6369
R5475 VDPWR.n2365 VDPWR.n2364 11.6369
R5476 VDPWR.n2364 VDPWR.n2361 11.6369
R5477 VDPWR.n2361 VDPWR.n2360 11.6369
R5478 VDPWR.n1409 VDPWR.n1406 11.6369
R5479 VDPWR.n1410 VDPWR.n1409 11.6369
R5480 VDPWR.n1413 VDPWR.n1410 11.6369
R5481 VDPWR.n1414 VDPWR.n1413 11.6369
R5482 VDPWR.n1417 VDPWR.n1414 11.6369
R5483 VDPWR.n1418 VDPWR.n1417 11.6369
R5484 VDPWR.n1421 VDPWR.n1418 11.6369
R5485 VDPWR.n1422 VDPWR.n1421 11.6369
R5486 VDPWR.n1425 VDPWR.n1422 11.6369
R5487 VDPWR.n1426 VDPWR.n1425 11.6369
R5488 VDPWR.n1431 VDPWR.n1430 11.6369
R5489 VDPWR.n1432 VDPWR.n1431 11.6369
R5490 VDPWR.n1432 VDPWR.n1233 11.6369
R5491 VDPWR.n1438 VDPWR.n1233 11.6369
R5492 VDPWR.n1439 VDPWR.n1438 11.6369
R5493 VDPWR.n1440 VDPWR.n1439 11.6369
R5494 VDPWR.n1440 VDPWR.n1231 11.6369
R5495 VDPWR.n1446 VDPWR.n1231 11.6369
R5496 VDPWR.n1447 VDPWR.n1446 11.6369
R5497 VDPWR.n1448 VDPWR.n1447 11.6369
R5498 VDPWR.n1448 VDPWR.n1224 11.6369
R5499 VDPWR.n1602 VDPWR.n1226 11.6369
R5500 VDPWR.n1596 VDPWR.n1226 11.6369
R5501 VDPWR.n1596 VDPWR.n1595 11.6369
R5502 VDPWR.n1595 VDPWR.n1594 11.6369
R5503 VDPWR.n1594 VDPWR.n1464 11.6369
R5504 VDPWR.n1497 VDPWR.n1464 11.6369
R5505 VDPWR.n1497 VDPWR.n1496 11.6369
R5506 VDPWR.n1517 VDPWR.n1496 11.6369
R5507 VDPWR.n1518 VDPWR.n1517 11.6369
R5508 VDPWR.n1519 VDPWR.n1518 11.6369
R5509 VDPWR.n1519 VDPWR.n815 11.6369
R5510 VDPWR.n2254 VDPWR.n816 11.6369
R5511 VDPWR.n2254 VDPWR.n2253 11.6369
R5512 VDPWR.n2253 VDPWR.n2252 11.6369
R5513 VDPWR.n2252 VDPWR.n2128 11.6369
R5514 VDPWR.n2165 VDPWR.n2128 11.6369
R5515 VDPWR.n2168 VDPWR.n2165 11.6369
R5516 VDPWR.n2169 VDPWR.n2168 11.6369
R5517 VDPWR.n2171 VDPWR.n2169 11.6369
R5518 VDPWR.n2171 VDPWR.n2170 11.6369
R5519 VDPWR.n2170 VDPWR.n2019 11.6369
R5520 VDPWR.n2019 VDPWR.n2017 11.6369
R5521 VDPWR.n2349 VDPWR.n2347 11.6369
R5522 VDPWR.n2347 VDPWR.n2344 11.6369
R5523 VDPWR.n2344 VDPWR.n2343 11.6369
R5524 VDPWR.n2343 VDPWR.n2340 11.6369
R5525 VDPWR.n2340 VDPWR.n2339 11.6369
R5526 VDPWR.n2339 VDPWR.n2336 11.6369
R5527 VDPWR.n2336 VDPWR.n2335 11.6369
R5528 VDPWR.n2335 VDPWR.n2332 11.6369
R5529 VDPWR.n2332 VDPWR.n2331 11.6369
R5530 VDPWR.n2331 VDPWR.n2329 11.6369
R5531 VDPWR.n2263 VDPWR.n2262 11.6369
R5532 VDPWR.n2265 VDPWR.n2263 11.6369
R5533 VDPWR.n2265 VDPWR.n2264 11.6369
R5534 VDPWR.n2264 VDPWR.n2043 11.6369
R5535 VDPWR.n2043 VDPWR.n2041 11.6369
R5536 VDPWR.n2284 VDPWR.n2041 11.6369
R5537 VDPWR.n2285 VDPWR.n2284 11.6369
R5538 VDPWR.n2287 VDPWR.n2285 11.6369
R5539 VDPWR.n2287 VDPWR.n2286 11.6369
R5540 VDPWR.n2286 VDPWR.n2026 11.6369
R5541 VDPWR.n2328 VDPWR.n2026 11.6369
R5542 VDPWR.n1073 VDPWR.n1070 11.6369
R5543 VDPWR.n1070 VDPWR.n1069 11.6369
R5544 VDPWR.n1069 VDPWR.n1066 11.6369
R5545 VDPWR.n1066 VDPWR.n1065 11.6369
R5546 VDPWR.n1065 VDPWR.n1062 11.6369
R5547 VDPWR.n1062 VDPWR.n1061 11.6369
R5548 VDPWR.n1061 VDPWR.n1058 11.6369
R5549 VDPWR.n1058 VDPWR.n1057 11.6369
R5550 VDPWR.n1057 VDPWR.n1055 11.6369
R5551 VDPWR.n1055 VDPWR.n913 11.6369
R5552 VDPWR.n1690 VDPWR.n1689 11.6369
R5553 VDPWR.n1693 VDPWR.n1690 11.6369
R5554 VDPWR.n1694 VDPWR.n1693 11.6369
R5555 VDPWR.n1697 VDPWR.n1694 11.6369
R5556 VDPWR.n1698 VDPWR.n1697 11.6369
R5557 VDPWR.n1701 VDPWR.n1698 11.6369
R5558 VDPWR.n1702 VDPWR.n1701 11.6369
R5559 VDPWR.n1705 VDPWR.n1702 11.6369
R5560 VDPWR.n1706 VDPWR.n1705 11.6369
R5561 VDPWR.n1709 VDPWR.n1706 11.6369
R5562 VDPWR.n1710 VDPWR.n1709 11.6369
R5563 VDPWR.n2319 VDPWR.n2316 11.6369
R5564 VDPWR.n2316 VDPWR.n2315 11.6369
R5565 VDPWR.n2315 VDPWR.n2312 11.6369
R5566 VDPWR.n2312 VDPWR.n2311 11.6369
R5567 VDPWR.n2311 VDPWR.n2308 11.6369
R5568 VDPWR.n2308 VDPWR.n2307 11.6369
R5569 VDPWR.n2307 VDPWR.n2304 11.6369
R5570 VDPWR.n2304 VDPWR.n2303 11.6369
R5571 VDPWR.n2303 VDPWR.n2301 11.6369
R5572 VDPWR.n2301 VDPWR.n1869 11.6369
R5573 VDPWR.n2410 VDPWR.n2408 11.6369
R5574 VDPWR.n2408 VDPWR.n2405 11.6369
R5575 VDPWR.n2405 VDPWR.n2404 11.6369
R5576 VDPWR.n2404 VDPWR.n2401 11.6369
R5577 VDPWR.n2401 VDPWR.n2400 11.6369
R5578 VDPWR.n2400 VDPWR.n2397 11.6369
R5579 VDPWR.n2397 VDPWR.n2396 11.6369
R5580 VDPWR.n2396 VDPWR.n2393 11.6369
R5581 VDPWR.n2393 VDPWR.n2392 11.6369
R5582 VDPWR.n2392 VDPWR.n2389 11.6369
R5583 VDPWR.n2389 VDPWR.n2388 11.6369
R5584 VDPWR.n1682 VDPWR.n1681 11.6369
R5585 VDPWR.n1681 VDPWR.n1678 11.6369
R5586 VDPWR.n1678 VDPWR.n1677 11.6369
R5587 VDPWR.n1677 VDPWR.n1674 11.6369
R5588 VDPWR.n1674 VDPWR.n1673 11.6369
R5589 VDPWR.n1673 VDPWR.n1670 11.6369
R5590 VDPWR.n1670 VDPWR.n1669 11.6369
R5591 VDPWR.n1669 VDPWR.n1666 11.6369
R5592 VDPWR.n1666 VDPWR.n1665 11.6369
R5593 VDPWR.n1665 VDPWR.n1663 11.6369
R5594 VDPWR.n1662 VDPWR.n1079 11.6369
R5595 VDPWR.n1080 VDPWR.n1079 11.6369
R5596 VDPWR.n1655 VDPWR.n1080 11.6369
R5597 VDPWR.n1655 VDPWR.n1654 11.6369
R5598 VDPWR.n1654 VDPWR.n1653 11.6369
R5599 VDPWR.n1653 VDPWR.n1082 11.6369
R5600 VDPWR.n1648 VDPWR.n1082 11.6369
R5601 VDPWR.n1648 VDPWR.n1647 11.6369
R5602 VDPWR.n1647 VDPWR.n1646 11.6369
R5603 VDPWR.n1646 VDPWR.n1085 11.6369
R5604 VDPWR.n1641 VDPWR.n1085 11.6369
R5605 VDPWR.n1803 VDPWR.n1802 11.6369
R5606 VDPWR.n1805 VDPWR.n1803 11.6369
R5607 VDPWR.n1805 VDPWR.n1804 11.6369
R5608 VDPWR.n1804 VDPWR.n863 11.6369
R5609 VDPWR.n1823 VDPWR.n863 11.6369
R5610 VDPWR.n1824 VDPWR.n1823 11.6369
R5611 VDPWR.n1825 VDPWR.n1824 11.6369
R5612 VDPWR.n1825 VDPWR.n849 11.6369
R5613 VDPWR.n2451 VDPWR.n849 11.6369
R5614 VDPWR.n2452 VDPWR.n2451 11.6369
R5615 VDPWR.n2453 VDPWR.n2452 11.6369
R5616 VDPWR.n2638 VDPWR.n2637 11.6369
R5617 VDPWR.n2637 VDPWR.n2636 11.6369
R5618 VDPWR.n2636 VDPWR.n2633 11.6369
R5619 VDPWR.n2633 VDPWR.n2632 11.6369
R5620 VDPWR.n2632 VDPWR.n2629 11.6369
R5621 VDPWR.n2413 VDPWR.n76 11.6369
R5622 VDPWR.n2415 VDPWR.n2413 11.6369
R5623 VDPWR.n2416 VDPWR.n2415 11.6369
R5624 VDPWR.n2418 VDPWR.n2416 11.6369
R5625 VDPWR.n2419 VDPWR.n2418 11.6369
R5626 VDPWR.n2729 VDPWR.n2728 11.4715
R5627 VDPWR.n1980 VDPWR.t16 10.1221
R5628 VDPWR.n1904 VDPWR.t72 10.1221
R5629 VDPWR.n1995 VDPWR.t296 10.1221
R5630 VDPWR.n2010 VDPWR.t297 10.1221
R5631 VDPWR.n2726 VDPWR.t187 9.88814
R5632 VDPWR.n2675 VDPWR.n2674 9.79932
R5633 VDPWR.n2598 VDPWR.t200 9.6005
R5634 VDPWR.n2603 VDPWR.t208 9.6005
R5635 VDPWR.n2580 VDPWR.t210 9.6005
R5636 VDPWR.n2573 VDPWR.t206 9.6005
R5637 VDPWR.n435 VDPWR.n434 9.6005
R5638 VDPWR.n434 VDPWR.n433 9.6005
R5639 VDPWR.n172 VDPWR.n171 9.6005
R5640 VDPWR.n171 VDPWR.n104 9.6005
R5641 VDPWR.n2712 VDPWR.n2711 9.58175
R5642 VDPWR.n694 VDPWR.n693 9.40114
R5643 VDPWR.n2563 VDPWR.n702 9.36264
R5644 VDPWR.n2542 VDPWR.n2537 9.36264
R5645 VDPWR.n2627 VDPWR.n2626 9.36264
R5646 VDPWR.n2562 VDPWR.n2561 9.3005
R5647 VDPWR.n2560 VDPWR.n701 9.3005
R5648 VDPWR.n2541 VDPWR.n2540 9.3005
R5649 VDPWR.n2539 VDPWR.n2538 9.3005
R5650 VDPWR.n2678 VDPWR.n2677 9.3005
R5651 VDPWR.n2676 VDPWR.n2653 9.3005
R5652 VDPWR.n2679 VDPWR.n2652 9.3005
R5653 VDPWR.n2710 VDPWR.n2709 9.3005
R5654 VDPWR.n2708 VDPWR.n2645 9.3005
R5655 VDPWR.n2707 VDPWR.n2706 9.3005
R5656 VDPWR.n2703 VDPWR.n2646 9.3005
R5657 VDPWR.n2702 VDPWR.n2701 9.3005
R5658 VDPWR.n2700 VDPWR.n2647 9.3005
R5659 VDPWR.n2699 VDPWR.n2698 9.3005
R5660 VDPWR.n2695 VDPWR.n2648 9.3005
R5661 VDPWR.n2694 VDPWR.n2693 9.3005
R5662 VDPWR.n2692 VDPWR.n2649 9.3005
R5663 VDPWR.n2691 VDPWR.n2690 9.3005
R5664 VDPWR.n2687 VDPWR.n2650 9.3005
R5665 VDPWR.n2686 VDPWR.n2685 9.3005
R5666 VDPWR.n2684 VDPWR.n2651 9.3005
R5667 VDPWR.n2683 VDPWR.n2682 9.3005
R5668 VDPWR.n642 VDPWR.n641 9.3005
R5669 VDPWR.n689 VDPWR.n611 9.3005
R5670 VDPWR.n688 VDPWR.n687 9.3005
R5671 VDPWR.n686 VDPWR.n612 9.3005
R5672 VDPWR.n685 VDPWR.n684 9.3005
R5673 VDPWR.n682 VDPWR.n613 9.3005
R5674 VDPWR.n681 VDPWR.n680 9.3005
R5675 VDPWR.n679 VDPWR.n614 9.3005
R5676 VDPWR.n678 VDPWR.n677 9.3005
R5677 VDPWR.n675 VDPWR.n615 9.3005
R5678 VDPWR.n674 VDPWR.n673 9.3005
R5679 VDPWR.n672 VDPWR.n616 9.3005
R5680 VDPWR.n671 VDPWR.n670 9.3005
R5681 VDPWR.n669 VDPWR.n617 9.3005
R5682 VDPWR.n668 VDPWR.n667 9.3005
R5683 VDPWR.n666 VDPWR.n618 9.3005
R5684 VDPWR.n665 VDPWR.n664 9.3005
R5685 VDPWR.n662 VDPWR.n619 9.3005
R5686 VDPWR.n661 VDPWR.n660 9.3005
R5687 VDPWR.n659 VDPWR.n620 9.3005
R5688 VDPWR.n658 VDPWR.n657 9.3005
R5689 VDPWR.n656 VDPWR.n621 9.3005
R5690 VDPWR.n655 VDPWR.n654 9.3005
R5691 VDPWR.n653 VDPWR.n622 9.3005
R5692 VDPWR.n652 VDPWR.n651 9.3005
R5693 VDPWR.n650 VDPWR.n623 9.3005
R5694 VDPWR.n649 VDPWR.n648 9.3005
R5695 VDPWR.n647 VDPWR.n624 9.3005
R5696 VDPWR.n646 VDPWR.n645 9.3005
R5697 VDPWR.n644 VDPWR.n625 9.3005
R5698 VDPWR.n643 VDPWR.n627 9.3005
R5699 VDPWR.n640 VDPWR.n629 9.3005
R5700 VDPWR.n639 VDPWR.n638 9.3005
R5701 VDPWR.n637 VDPWR.n630 9.3005
R5702 VDPWR.n636 VDPWR.n635 9.3005
R5703 VDPWR.n634 VDPWR.n631 9.3005
R5704 VDPWR.n633 VDPWR.n632 9.3005
R5705 VDPWR.n4 VDPWR.n3 9.3005
R5706 VDPWR.n496 VDPWR.n495 9.3005
R5707 VDPWR.n494 VDPWR.n245 9.3005
R5708 VDPWR.n493 VDPWR.n492 9.3005
R5709 VDPWR.n475 VDPWR.n474 9.3005
R5710 VDPWR.n476 VDPWR.n253 9.3005
R5711 VDPWR.n478 VDPWR.n477 9.3005
R5712 VDPWR.n479 VDPWR.n252 9.3005
R5713 VDPWR.n481 VDPWR.n480 9.3005
R5714 VDPWR.n482 VDPWR.n250 9.3005
R5715 VDPWR.n484 VDPWR.n483 9.3005
R5716 VDPWR.n485 VDPWR.n249 9.3005
R5717 VDPWR.n487 VDPWR.n486 9.3005
R5718 VDPWR.n488 VDPWR.n248 9.3005
R5719 VDPWR.n490 VDPWR.n489 9.3005
R5720 VDPWR.n491 VDPWR.n246 9.3005
R5721 VDPWR.n502 VDPWR.n501 9.3005
R5722 VDPWR.n503 VDPWR.n244 9.3005
R5723 VDPWR.n505 VDPWR.n504 9.3005
R5724 VDPWR.n506 VDPWR.n241 9.3005
R5725 VDPWR.n508 VDPWR.n507 9.3005
R5726 VDPWR.n509 VDPWR.n240 9.3005
R5727 VDPWR.n511 VDPWR.n510 9.3005
R5728 VDPWR.n521 VDPWR.n520 9.3005
R5729 VDPWR.n522 VDPWR.n232 9.3005
R5730 VDPWR.n524 VDPWR.n523 9.3005
R5731 VDPWR.n525 VDPWR.n229 9.3005
R5732 VDPWR.n527 VDPWR.n526 9.3005
R5733 VDPWR.n528 VDPWR.n228 9.3005
R5734 VDPWR.n530 VDPWR.n529 9.3005
R5735 VDPWR.n531 VDPWR.n226 9.3005
R5736 VDPWR.n532 VDPWR.n224 9.3005
R5737 VDPWR.n534 VDPWR.n533 9.3005
R5738 VDPWR.n535 VDPWR.n223 9.3005
R5739 VDPWR.n537 VDPWR.n536 9.3005
R5740 VDPWR.n538 VDPWR.n221 9.3005
R5741 VDPWR.n540 VDPWR.n539 9.3005
R5742 VDPWR.n541 VDPWR.n220 9.3005
R5743 VDPWR.n543 VDPWR.n542 9.3005
R5744 VDPWR.n544 VDPWR.n217 9.3005
R5745 VDPWR.n546 VDPWR.n545 9.3005
R5746 VDPWR.n547 VDPWR.n216 9.3005
R5747 VDPWR.n549 VDPWR.n548 9.3005
R5748 VDPWR.n550 VDPWR.n214 9.3005
R5749 VDPWR.n551 VDPWR.n212 9.3005
R5750 VDPWR.n553 VDPWR.n552 9.3005
R5751 VDPWR.n554 VDPWR.n211 9.3005
R5752 VDPWR.n556 VDPWR.n555 9.3005
R5753 VDPWR.n557 VDPWR.n209 9.3005
R5754 VDPWR.n559 VDPWR.n558 9.3005
R5755 VDPWR.n560 VDPWR.n208 9.3005
R5756 VDPWR.n562 VDPWR.n561 9.3005
R5757 VDPWR.n563 VDPWR.n207 9.3005
R5758 VDPWR.n565 VDPWR.n564 9.3005
R5759 VDPWR.n567 VDPWR.n566 9.3005
R5760 VDPWR.n568 VDPWR.n203 9.3005
R5761 VDPWR.n570 VDPWR.n569 9.3005
R5762 VDPWR.n571 VDPWR.n202 9.3005
R5763 VDPWR.n573 VDPWR.n572 9.3005
R5764 VDPWR.n574 VDPWR.n201 9.3005
R5765 VDPWR.n576 VDPWR.n575 9.3005
R5766 VDPWR.n577 VDPWR.n96 9.3005
R5767 VDPWR.n579 VDPWR.n578 9.3005
R5768 VDPWR.n200 VDPWR.n95 9.3005
R5769 VDPWR.n199 VDPWR.n198 9.3005
R5770 VDPWR.n197 VDPWR.n97 9.3005
R5771 VDPWR.n194 VDPWR.n193 9.3005
R5772 VDPWR.n192 VDPWR.n98 9.3005
R5773 VDPWR.n191 VDPWR.n190 9.3005
R5774 VDPWR.n188 VDPWR.n99 9.3005
R5775 VDPWR.n187 VDPWR.n186 9.3005
R5776 VDPWR.n185 VDPWR.n184 9.3005
R5777 VDPWR.n183 VDPWR.n101 9.3005
R5778 VDPWR.n182 VDPWR.n181 9.3005
R5779 VDPWR.n180 VDPWR.n102 9.3005
R5780 VDPWR.n179 VDPWR.n178 9.3005
R5781 VDPWR.n177 VDPWR.n103 9.3005
R5782 VDPWR.n176 VDPWR.n175 9.3005
R5783 VDPWR.n174 VDPWR.n104 9.3005
R5784 VDPWR.n173 VDPWR.n172 9.3005
R5785 VDPWR.n169 VDPWR.n105 9.3005
R5786 VDPWR.n168 VDPWR.n167 9.3005
R5787 VDPWR.n166 VDPWR.n106 9.3005
R5788 VDPWR.n165 VDPWR.n164 9.3005
R5789 VDPWR.n162 VDPWR.n107 9.3005
R5790 VDPWR.n161 VDPWR.n160 9.3005
R5791 VDPWR.n159 VDPWR.n158 9.3005
R5792 VDPWR.n157 VDPWR.n110 9.3005
R5793 VDPWR.n156 VDPWR.n155 9.3005
R5794 VDPWR.n154 VDPWR.n111 9.3005
R5795 VDPWR.n153 VDPWR.n152 9.3005
R5796 VDPWR.n151 VDPWR.n112 9.3005
R5797 VDPWR.n150 VDPWR.n149 9.3005
R5798 VDPWR.n148 VDPWR.n113 9.3005
R5799 VDPWR.n147 VDPWR.n146 9.3005
R5800 VDPWR.n145 VDPWR.n115 9.3005
R5801 VDPWR.n144 VDPWR.n143 9.3005
R5802 VDPWR.n142 VDPWR.n141 9.3005
R5803 VDPWR.n140 VDPWR.n118 9.3005
R5804 VDPWR.n139 VDPWR.n137 9.3005
R5805 VDPWR.n136 VDPWR.n119 9.3005
R5806 VDPWR.n135 VDPWR.n134 9.3005
R5807 VDPWR.n133 VDPWR.n120 9.3005
R5808 VDPWR.n132 VDPWR.n131 9.3005
R5809 VDPWR.n130 VDPWR.n121 9.3005
R5810 VDPWR.n129 VDPWR.n128 9.3005
R5811 VDPWR.n127 VDPWR.n122 9.3005
R5812 VDPWR.n519 VDPWR.n233 9.3005
R5813 VDPWR.n516 VDPWR.n235 9.3005
R5814 VDPWR.n518 VDPWR.n517 9.3005
R5815 VDPWR.n512 VDPWR.n239 9.3005
R5816 VDPWR.n513 VDPWR.n236 9.3005
R5817 VDPWR.n515 VDPWR.n514 9.3005
R5818 VDPWR.n354 VDPWR.n261 9.3005
R5819 VDPWR.n353 VDPWR.n352 9.3005
R5820 VDPWR.n351 VDPWR.n262 9.3005
R5821 VDPWR.n350 VDPWR.n349 9.3005
R5822 VDPWR.n348 VDPWR.n263 9.3005
R5823 VDPWR.n346 VDPWR.n345 9.3005
R5824 VDPWR.n344 VDPWR.n264 9.3005
R5825 VDPWR.n343 VDPWR.n342 9.3005
R5826 VDPWR.n330 VDPWR.n265 9.3005
R5827 VDPWR.n329 VDPWR.n328 9.3005
R5828 VDPWR.n327 VDPWR.n267 9.3005
R5829 VDPWR.n326 VDPWR.n325 9.3005
R5830 VDPWR.n324 VDPWR.n268 9.3005
R5831 VDPWR.n323 VDPWR.n322 9.3005
R5832 VDPWR.n321 VDPWR.n270 9.3005
R5833 VDPWR.n320 VDPWR.n319 9.3005
R5834 VDPWR.n318 VDPWR.n271 9.3005
R5835 VDPWR.n317 VDPWR.n316 9.3005
R5836 VDPWR.n315 VDPWR.n285 9.3005
R5837 VDPWR.n314 VDPWR.n313 9.3005
R5838 VDPWR.n312 VDPWR.n286 9.3005
R5839 VDPWR.n311 VDPWR.n287 9.3005
R5840 VDPWR.n310 VDPWR.n309 9.3005
R5841 VDPWR.n308 VDPWR.n289 9.3005
R5842 VDPWR.n307 VDPWR.n306 9.3005
R5843 VDPWR.n2625 VDPWR.n78 9.3005
R5844 VDPWR.n2624 VDPWR.n2623 9.3005
R5845 VDPWR.n608 VDPWR.n607 9.3005
R5846 VDPWR.n606 VDPWR.n82 9.3005
R5847 VDPWR.n605 VDPWR.n604 9.3005
R5848 VDPWR.n603 VDPWR.n83 9.3005
R5849 VDPWR.n602 VDPWR.n601 9.3005
R5850 VDPWR.n600 VDPWR.n84 9.3005
R5851 VDPWR.n599 VDPWR.n598 9.3005
R5852 VDPWR.n597 VDPWR.n85 9.3005
R5853 VDPWR.n596 VDPWR.n595 9.3005
R5854 VDPWR.n594 VDPWR.n87 9.3005
R5855 VDPWR.n593 VDPWR.n592 9.3005
R5856 VDPWR.n590 VDPWR.n88 9.3005
R5857 VDPWR.n589 VDPWR.n588 9.3005
R5858 VDPWR.n587 VDPWR.n89 9.3005
R5859 VDPWR.n586 VDPWR.n91 9.3005
R5860 VDPWR.n424 VDPWR.n90 9.3005
R5861 VDPWR.n426 VDPWR.n425 9.3005
R5862 VDPWR.n427 VDPWR.n420 9.3005
R5863 VDPWR.n429 VDPWR.n428 9.3005
R5864 VDPWR.n430 VDPWR.n419 9.3005
R5865 VDPWR.n432 VDPWR.n431 9.3005
R5866 VDPWR.n433 VDPWR.n417 9.3005
R5867 VDPWR.n436 VDPWR.n435 9.3005
R5868 VDPWR.n437 VDPWR.n416 9.3005
R5869 VDPWR.n439 VDPWR.n438 9.3005
R5870 VDPWR.n440 VDPWR.n415 9.3005
R5871 VDPWR.n414 VDPWR.n373 9.3005
R5872 VDPWR.n413 VDPWR.n412 9.3005
R5873 VDPWR.n411 VDPWR.n374 9.3005
R5874 VDPWR.n410 VDPWR.n409 9.3005
R5875 VDPWR.n408 VDPWR.n375 9.3005
R5876 VDPWR.n407 VDPWR.n406 9.3005
R5877 VDPWR.n405 VDPWR.n376 9.3005
R5878 VDPWR.n404 VDPWR.n403 9.3005
R5879 VDPWR.n402 VDPWR.n377 9.3005
R5880 VDPWR.n401 VDPWR.n400 9.3005
R5881 VDPWR.n399 VDPWR.n378 9.3005
R5882 VDPWR.n397 VDPWR.n396 9.3005
R5883 VDPWR.n395 VDPWR.n394 9.3005
R5884 VDPWR.n393 VDPWR.n381 9.3005
R5885 VDPWR.n392 VDPWR.n391 9.3005
R5886 VDPWR.n390 VDPWR.n382 9.3005
R5887 VDPWR.n389 VDPWR.n388 9.3005
R5888 VDPWR.n387 VDPWR.n383 9.3005
R5889 VDPWR.n386 VDPWR.n385 9.3005
R5890 VDPWR.n2714 VDPWR.t235 9.10772
R5891 VDPWR.t235 VDPWR.t135 8.67615
R5892 VDPWR.n8 VDPWR.n5 8.50653
R5893 VDPWR.n610 VDPWR.n609 8.31939
R5894 VDPWR.t235 VDPWR.n2640 7.60149
R5895 VDPWR.n609 VDPWR.n81 7.56834
R5896 VDPWR.n500 VDPWR.n498 7.37605
R5897 VDPWR.n693 VDPWR.n692 7.22808
R5898 VDPWR.n298 VDPWR.n297 7.11161
R5899 VDPWR.n361 VDPWR.n260 7.11161
R5900 VDPWR.n126 VDPWR.n124 7.07105
R5901 VDPWR.n2745 VDPWR.n2744 6.86155
R5902 VDPWR.n384 VDPWR.n2 6.86155
R5903 VDPWR.n473 VDPWR.n254 6.86152
R5904 VDPWR.n1603 VDPWR.n1602 6.72373
R5905 VDPWR.n2478 VDPWR.n816 6.72373
R5906 VDPWR.n2262 VDPWR.n846 6.72373
R5907 VDPWR.n2420 VDPWR.n2410 6.72373
R5908 VDPWR.n1802 VDPWR.n882 6.72373
R5909 VDPWR.n2638 VDPWR.n75 6.72373
R5910 VDPWR.n357 VDPWR.n356 6.69883
R5911 VDPWR.n2662 VDPWR.n2660 6.4005
R5912 VDPWR.n2666 VDPWR.n2665 6.4005
R5913 VDPWR.n663 VDPWR.n618 6.4005
R5914 VDPWR.n141 VDPWR.n117 6.4005
R5915 VDPWR.n161 VDPWR.n109 6.4005
R5916 VDPWR.n187 VDPWR.n100 6.4005
R5917 VDPWR.n580 VDPWR.n579 6.4005
R5918 VDPWR.n567 VDPWR.n206 6.4005
R5919 VDPWR.n219 VDPWR.n216 6.4005
R5920 VDPWR.n231 VDPWR.n228 6.4005
R5921 VDPWR.n243 VDPWR.n240 6.4005
R5922 VDPWR.n317 VDPWR.n285 6.4005
R5923 VDPWR.n319 VDPWR.n270 6.4005
R5924 VDPWR.n349 VDPWR.n348 6.4005
R5925 VDPWR.n2617 VDPWR.n2616 6.36829
R5926 VDPWR.n1603 VDPWR.n1224 6.20656
R5927 VDPWR.n2478 VDPWR.n815 6.20656
R5928 VDPWR.n1710 VDPWR.n75 6.20656
R5929 VDPWR.n1641 VDPWR.n882 6.20656
R5930 VDPWR.n2453 VDPWR.n846 6.20656
R5931 VDPWR.n2420 VDPWR.n2419 6.20656
R5932 VDPWR.n2628 VDPWR.n76 6.07727
R5933 VDPWR.t1 VDPWR.n2669 6.07198
R5934 VDPWR.n305 VDPWR.n303 5.97271
R5935 VDPWR.n2609 VDPWR.n2594 5.81868
R5936 VDPWR.n628 VDPWR.n6 5.68939
R5937 VDPWR.n626 VDPWR.n6 5.68939
R5938 VDPWR.n398 VDPWR.n371 5.68939
R5939 VDPWR.n2618 VDPWR.n2617 5.6447
R5940 VDPWR.n2629 VDPWR.n2628 5.5601
R5941 VDPWR.n2120 VDPWR.n2119 5.51161
R5942 VDPWR.n1797 VDPWR.n1796 5.51161
R5943 VDPWR.n2234 VDPWR.n2232 5.51161
R5944 VDPWR.n1976 VDPWR.n1975 5.51161
R5945 VDPWR.n1579 VDPWR.n1577 5.51161
R5946 VDPWR.n731 VDPWR.n708 5.51161
R5947 VDPWR.n1268 VDPWR.n1236 5.51161
R5948 VDPWR.n1053 VDPWR.n935 5.51161
R5949 VDPWR.n1185 VDPWR.n1133 5.51161
R5950 VDPWR.n2755 VDPWR.n2746 5.19967
R5951 VDPWR.n1405 VDPWR.n1404 5.1717
R5952 VDPWR.n1074 VDPWR.n1054 5.1717
R5953 VDPWR.n1132 VDPWR.n1078 5.1717
R5954 VDPWR.n379 VDPWR.n371 4.97828
R5955 VDPWR.n2381 VDPWR.n2016 4.9157
R5956 VDPWR.n2352 VDPWR.n2351 4.9157
R5957 VDPWR.n2321 VDPWR.n2320 4.9157
R5958 VDPWR.n2673 VDPWR.n2656 4.88834
R5959 VDPWR.n281 VDPWR.n280 4.57193
R5960 VDPWR.n338 VDPWR.n332 4.57193
R5961 VDPWR.n2539 VDPWR.n699 4.5005
R5962 VDPWR.n2564 VDPWR.n701 4.5005
R5963 VDPWR.n2567 VDPWR.n700 4.5005
R5964 VDPWR.n2569 VDPWR.n2568 4.5005
R5965 VDPWR.n2568 VDPWR.n2567 4.5005
R5966 VDPWR.n2591 VDPWR.n2590 4.5005
R5967 VDPWR.n2624 VDPWR.n2620 4.5005
R5968 VDPWR.n459 VDPWR.n251 4.49344
R5969 VDPWR.n460 VDPWR.n459 4.49344
R5970 VDPWR.n453 VDPWR.n247 4.49344
R5971 VDPWR.n454 VDPWR.n453 4.49344
R5972 VDPWR.n2617 VDPWR.n2611 4.42387
R5973 VDPWR.n301 VDPWR.n290 4.36399
R5974 VDPWR.n362 VDPWR.n359 4.36399
R5975 VDPWR.n1399 VDPWR.t312 4.33832
R5976 VDPWR.t90 VDPWR.n1338 4.33832
R5977 VDPWR.n1340 VDPWR.t96 4.33832
R5978 VDPWR.n1387 VDPWR.t113 4.33832
R5979 VDPWR.n1382 VDPWR.n1381 4.26717
R5980 VDPWR.n1381 VDPWR.n1350 4.26717
R5981 VDPWR.n1376 VDPWR.n1350 4.26717
R5982 VDPWR.n1376 VDPWR.n1375 4.26717
R5983 VDPWR.n1375 VDPWR.n1374 4.26717
R5984 VDPWR.n1374 VDPWR.n1359 4.26717
R5985 VDPWR.n1369 VDPWR.n1359 4.26717
R5986 VDPWR.n1369 VDPWR.n1368 4.26717
R5987 VDPWR.n1368 VDPWR.n1228 4.26717
R5988 VDPWR.n1455 VDPWR.n1228 4.26717
R5989 VDPWR.n1455 VDPWR.n1225 4.26717
R5990 VDPWR.n2500 VDPWR.n789 4.26717
R5991 VDPWR.n790 VDPWR.n789 4.26717
R5992 VDPWR.n2493 VDPWR.n790 4.26717
R5993 VDPWR.n2493 VDPWR.n2492 4.26717
R5994 VDPWR.n2492 VDPWR.n2491 4.26717
R5995 VDPWR.n2491 VDPWR.n800 4.26717
R5996 VDPWR.n2486 VDPWR.n800 4.26717
R5997 VDPWR.n2486 VDPWR.n2485 4.26717
R5998 VDPWR.n2485 VDPWR.n2484 4.26717
R5999 VDPWR.n2484 VDPWR.n809 4.26717
R6000 VDPWR.n2479 VDPWR.n809 4.26717
R6001 VDPWR.n2472 VDPWR.n820 4.26717
R6002 VDPWR.n2472 VDPWR.n2471 4.26717
R6003 VDPWR.n2471 VDPWR.n2470 4.26717
R6004 VDPWR.n2470 VDPWR.n828 4.26717
R6005 VDPWR.n2465 VDPWR.n828 4.26717
R6006 VDPWR.n2465 VDPWR.n2464 4.26717
R6007 VDPWR.n2464 VDPWR.n2463 4.26717
R6008 VDPWR.n2463 VDPWR.n837 4.26717
R6009 VDPWR.n2458 VDPWR.n837 4.26717
R6010 VDPWR.n2458 VDPWR.n2457 4.26717
R6011 VDPWR.n2457 VDPWR.n2456 4.26717
R6012 VDPWR.n1608 VDPWR.n1098 4.26717
R6013 VDPWR.n1614 VDPWR.n1098 4.26717
R6014 VDPWR.n1614 VDPWR.n1096 4.26717
R6015 VDPWR.n1620 VDPWR.n1096 4.26717
R6016 VDPWR.n1620 VDPWR.n1094 4.26717
R6017 VDPWR.n1626 VDPWR.n1094 4.26717
R6018 VDPWR.n1626 VDPWR.n1092 4.26717
R6019 VDPWR.n1633 VDPWR.n1092 4.26717
R6020 VDPWR.n1633 VDPWR.n1088 4.26717
R6021 VDPWR.n1638 VDPWR.n1088 4.26717
R6022 VDPWR.n1639 VDPWR.n1638 4.26717
R6023 VDPWR.n1733 VDPWR.n888 4.26717
R6024 VDPWR.n890 VDPWR.n888 4.26717
R6025 VDPWR.n1726 VDPWR.n890 4.26717
R6026 VDPWR.n1726 VDPWR.n1725 4.26717
R6027 VDPWR.n1725 VDPWR.n1724 4.26717
R6028 VDPWR.n1724 VDPWR.n900 4.26717
R6029 VDPWR.n1719 VDPWR.n900 4.26717
R6030 VDPWR.n1719 VDPWR.n1718 4.26717
R6031 VDPWR.n1718 VDPWR.n1717 4.26717
R6032 VDPWR.n1717 VDPWR.n911 4.26717
R6033 VDPWR.n1712 VDPWR.n911 4.26717
R6034 VDPWR.n2442 VDPWR.n1842 4.26717
R6035 VDPWR.n1844 VDPWR.n1842 4.26717
R6036 VDPWR.n2435 VDPWR.n1844 4.26717
R6037 VDPWR.n2435 VDPWR.n2434 4.26717
R6038 VDPWR.n2434 VDPWR.n2433 4.26717
R6039 VDPWR.n2433 VDPWR.n1854 4.26717
R6040 VDPWR.n2428 VDPWR.n1854 4.26717
R6041 VDPWR.n2428 VDPWR.n2427 4.26717
R6042 VDPWR.n2427 VDPWR.n2426 4.26717
R6043 VDPWR.n2426 VDPWR.n1863 4.26717
R6044 VDPWR.n2421 VDPWR.n1863 4.26717
R6045 VDPWR VDPWR.n2756 4.1224
R6046 VDPWR.n1603 VDPWR.n1225 3.98272
R6047 VDPWR.n2479 VDPWR.n2478 3.98272
R6048 VDPWR.n2456 VDPWR.n846 3.98272
R6049 VDPWR.n1639 VDPWR.n882 3.98272
R6050 VDPWR.n1712 VDPWR.n75 3.98272
R6051 VDPWR.n2421 VDPWR.n2420 3.98272
R6052 VDPWR.n462 VDPWR.n461 3.8278
R6053 VDPWR.n469 VDPWR.n468 3.8278
R6054 VDPWR.n456 VDPWR.n455 3.8278
R6055 VDPWR.n1985 VDPWR.n1984 3.7893
R6056 VDPWR.n1992 VDPWR.n1906 3.7893
R6057 VDPWR.n1991 VDPWR.n1908 3.7893
R6058 VDPWR.n1907 VDPWR.n1902 3.7893
R6059 VDPWR.n2000 VDPWR.n1999 3.7893
R6060 VDPWR.n1900 VDPWR.n1899 3.7893
R6061 VDPWR.n2008 VDPWR.n1896 3.7893
R6062 VDPWR.n2007 VDPWR.n1897 3.7893
R6063 VDPWR.n2014 VDPWR.n1892 3.7893
R6064 VDPWR.n1582 VDPWR.n1581 3.7893
R6065 VDPWR.n1472 VDPWR.n1471 3.7893
R6066 VDPWR.n1590 VDPWR.n1468 3.7893
R6067 VDPWR.n1589 VDPWR.n1469 3.7893
R6068 VDPWR.n1505 VDPWR.n1503 3.7893
R6069 VDPWR.n1506 VDPWR.n1502 3.7893
R6070 VDPWR.n1513 VDPWR.n1511 3.7893
R6071 VDPWR.n1512 VDPWR.n1490 3.7893
R6072 VDPWR.n1524 VDPWR.n1523 3.7893
R6073 VDPWR.n1265 VDPWR.n1264 3.7893
R6074 VDPWR.n1397 VDPWR.n1241 3.7893
R6075 VDPWR.n1396 VDPWR.n1242 3.7893
R6076 VDPWR.n1326 VDPWR.n1324 3.7893
R6077 VDPWR.n1329 VDPWR.n1328 3.7893
R6078 VDPWR.n1336 VDPWR.n1330 3.7893
R6079 VDPWR.n1335 VDPWR.n1332 3.7893
R6080 VDPWR.n1331 VDPWR.n1263 3.7893
R6081 VDPWR.n1391 VDPWR.n1390 3.7893
R6082 VDPWR.n2553 VDPWR.n709 3.7893
R6083 VDPWR.n2513 VDPWR.n2509 3.7893
R6084 VDPWR.n2516 VDPWR.n2515 3.7893
R6085 VDPWR.n2520 VDPWR.n2519 3.7893
R6086 VDPWR.n2524 VDPWR.n2507 3.7893
R6087 VDPWR.n2525 VDPWR.n2506 3.7893
R6088 VDPWR.n2530 VDPWR.n2528 3.7893
R6089 VDPWR.n2529 VDPWR.n730 3.7893
R6090 VDPWR.n2548 VDPWR.n2547 3.7893
R6091 VDPWR.n2239 VDPWR.n2238 3.7893
R6092 VDPWR.n2137 VDPWR.n2136 3.7893
R6093 VDPWR.n2247 VDPWR.n2133 3.7893
R6094 VDPWR.n2246 VDPWR.n2134 3.7893
R6095 VDPWR.n2160 VDPWR.n2158 3.7893
R6096 VDPWR.n2159 VDPWR.n2157 3.7893
R6097 VDPWR.n2176 VDPWR.n2175 3.7893
R6098 VDPWR.n2154 VDPWR.n2153 3.7893
R6099 VDPWR.n2354 VDPWR.n2023 3.7893
R6100 VDPWR.n1048 VDPWR.n936 3.7893
R6101 VDPWR.n1047 VDPWR.n938 3.7893
R6102 VDPWR.n969 VDPWR.n967 3.7893
R6103 VDPWR.n968 VDPWR.n965 3.7893
R6104 VDPWR.n976 VDPWR.n975 3.7893
R6105 VDPWR.n962 VDPWR.n961 3.7893
R6106 VDPWR.n984 VDPWR.n958 3.7893
R6107 VDPWR.n983 VDPWR.n956 3.7893
R6108 VDPWR.n991 VDPWR.n955 3.7893
R6109 VDPWR.n1192 VDPWR.n1188 3.7893
R6110 VDPWR.n1191 VDPWR.n1127 3.7893
R6111 VDPWR.n1198 VDPWR.n1126 3.7893
R6112 VDPWR.n1199 VDPWR.n1125 3.7893
R6113 VDPWR.n1204 VDPWR.n1202 3.7893
R6114 VDPWR.n1203 VDPWR.n1122 3.7893
R6115 VDPWR.n1211 VDPWR.n1210 3.7893
R6116 VDPWR.n1123 VDPWR.n1102 3.7893
R6117 VDPWR.n1217 VDPWR.n1216 3.7893
R6118 VDPWR.n1810 VDPWR.n1809 3.7893
R6119 VDPWR.n876 VDPWR.n875 3.7893
R6120 VDPWR.n1818 VDPWR.n868 3.7893
R6121 VDPWR.n1817 VDPWR.n869 3.7893
R6122 VDPWR.n873 VDPWR.n872 3.7893
R6123 VDPWR.n871 VDPWR.n860 3.7893
R6124 VDPWR.n1831 VDPWR.n1830 3.7893
R6125 VDPWR.n858 VDPWR.n857 3.7893
R6126 VDPWR.n2446 VDPWR.n854 3.7893
R6127 VDPWR.n2270 VDPWR.n2269 3.7893
R6128 VDPWR.n2056 VDPWR.n2055 3.7893
R6129 VDPWR.n2278 VDPWR.n2047 3.7893
R6130 VDPWR.n2277 VDPWR.n2048 3.7893
R6131 VDPWR.n2053 VDPWR.n2052 3.7893
R6132 VDPWR.n2050 VDPWR.n2037 3.7893
R6133 VDPWR.n2292 VDPWR.n2291 3.7893
R6134 VDPWR.n2035 VDPWR.n2034 3.7893
R6135 VDPWR.n2323 VDPWR.n2031 3.7893
R6136 VDPWR.n2751 VDPWR.n2748 3.4105
R6137 VDPWR.n2753 VDPWR.n2748 3.4105
R6138 VDPWR.n2755 VDPWR.n2748 3.4105
R6139 VDPWR.n2754 VDPWR.n2753 3.4105
R6140 VDPWR.n2755 VDPWR.n2754 3.4105
R6141 VDPWR.n2753 VDPWR.n2747 3.4105
R6142 VDPWR.n2755 VDPWR.n2747 3.4105
R6143 VDPWR.n2756 VDPWR.n2755 3.4105
R6144 VDPWR.n394 VDPWR.n380 3.2005
R6145 VDPWR.n196 VDPWR.n194 3.2005
R6146 VDPWR.n552 VDPWR.n213 3.2005
R6147 VDPWR.n533 VDPWR.n225 3.2005
R6148 VDPWR.n514 VDPWR.n237 3.2005
R6149 VDPWR.t199 VDPWR.n51 3.13108
R6150 VDPWR.t273 VDPWR.t61 3.03624
R6151 VDPWR.n2611 VDPWR.n2610 2.986
R6152 VDPWR.n466 VDPWR.n465 2.8779
R6153 VDPWR.n467 VDPWR.n466 2.8779
R6154 VDPWR.n2579 VDPWR.n2576 2.86505
R6155 VDPWR.n2581 VDPWR.n2575 2.86505
R6156 VDPWR.n2583 VDPWR.n2582 2.86505
R6157 VDPWR.n2584 VDPWR.n2572 2.86505
R6158 VDPWR.n2584 VDPWR.n2583 2.86505
R6159 VDPWR.n2576 VDPWR.n2575 2.86505
R6160 VDPWR.n2587 VDPWR.n2572 2.86505
R6161 VDPWR.n2582 VDPWR.n2581 2.86505
R6162 VDPWR.n2602 VDPWR.n2600 2.86505
R6163 VDPWR.n2601 VDPWR.n2597 2.86505
R6164 VDPWR.n2605 VDPWR.n2604 2.86505
R6165 VDPWR.n2604 VDPWR.n2594 2.86505
R6166 VDPWR.n2602 VDPWR.n2601 2.86505
R6167 VDPWR.n2605 VDPWR.n2597 2.86505
R6168 VDPWR.n284 VDPWR.n273 2.82018
R6169 VDPWR.n279 VDPWR.n278 2.82018
R6170 VDPWR.n341 VDPWR.n340 2.82018
R6171 VDPWR.n339 VDPWR.n334 2.82018
R6172 VDPWR.t209 VDPWR.n37 2.68393
R6173 VDPWR.n2501 VDPWR.n786 2.6629
R6174 VDPWR.n2016 VDPWR.n2015 2.6629
R6175 VDPWR.n1578 VDPWR.n1222 2.6629
R6176 VDPWR.n1492 VDPWR.n1491 2.6629
R6177 VDPWR.n1345 VDPWR.n1320 2.6629
R6178 VDPWR.n1383 VDPWR.n1346 2.6629
R6179 VDPWR.n2502 VDPWR.n783 2.6629
R6180 VDPWR.n2233 VDPWR.n818 2.6629
R6181 VDPWR.n2353 VDPWR.n2352 2.6629
R6182 VDPWR.n992 VDPWR.n885 2.6629
R6183 VDPWR.n1221 VDPWR.n1100 2.6629
R6184 VDPWR.n1798 VDPWR.n1734 2.6629
R6185 VDPWR.n2445 VDPWR.n2444 2.6629
R6186 VDPWR.n2443 VDPWR.n1839 2.6629
R6187 VDPWR.n2322 VDPWR.n2321 2.6629
R6188 VDPWR.n297 VDPWR.n296 2.6474
R6189 VDPWR.n298 VDPWR.n290 2.6474
R6190 VDPWR.n363 VDPWR.n260 2.6474
R6191 VDPWR.n362 VDPWR.n361 2.6474
R6192 VDPWR.n1976 VDPWR.n786 2.4581
R6193 VDPWR.n1579 VDPWR.n1578 2.4581
R6194 VDPWR.n1491 VDPWR.n818 2.4581
R6195 VDPWR.n1404 VDPWR.n1236 2.4581
R6196 VDPWR.n1383 VDPWR.n1345 2.4581
R6197 VDPWR.n1346 VDPWR.n708 2.4581
R6198 VDPWR.n2502 VDPWR.n2501 2.4581
R6199 VDPWR.n2234 VDPWR.n2233 2.4581
R6200 VDPWR.n1054 VDPWR.n1053 2.4581
R6201 VDPWR.n1734 VDPWR.n885 2.4581
R6202 VDPWR.n1133 VDPWR.n1132 2.4581
R6203 VDPWR.n1222 VDPWR.n1221 2.4581
R6204 VDPWR.n1798 VDPWR.n1797 2.4581
R6205 VDPWR.n2444 VDPWR.n2443 2.4581
R6206 VDPWR.n2120 VDPWR.n1839 2.4581
R6207 VDPWR.n2616 VDPWR.n2615 2.44675
R6208 VDPWR.n2616 VDPWR.n2612 2.44675
R6209 VDPWR.n2611 VDPWR.n694 2.31324
R6210 VDPWR.n2571 VDPWR.n695 2.26187
R6211 VDPWR.n2569 VDPWR.n697 2.24063
R6212 VDPWR.n698 VDPWR.n696 2.24063
R6213 VDPWR.n2592 VDPWR.n2570 2.24063
R6214 VDPWR.n2593 VDPWR.n695 2.24063
R6215 VDPWR.n2566 VDPWR.n2565 2.24063
R6216 VDPWR.n2589 VDPWR.n2588 2.24063
R6217 VDPWR.n2537 VDPWR.n699 2.22018
R6218 VDPWR.n2564 VDPWR.n2563 2.22018
R6219 VDPWR.n2626 VDPWR.n2620 2.22018
R6220 VDPWR.n1383 VDPWR.n1382 2.18124
R6221 VDPWR.n2501 VDPWR.n2500 2.18124
R6222 VDPWR.n820 VDPWR.n818 2.18124
R6223 VDPWR.n1608 VDPWR.n1222 2.18124
R6224 VDPWR.n1734 VDPWR.n1733 2.18124
R6225 VDPWR.n2443 VDPWR.n2442 2.18124
R6226 VDPWR.n1983 VDPWR.n1976 2.1509
R6227 VDPWR.n1580 VDPWR.n1579 2.1509
R6228 VDPWR.n1238 VDPWR.n1236 2.1509
R6229 VDPWR.n2554 VDPWR.n708 2.1509
R6230 VDPWR.n2235 VDPWR.n2234 2.1509
R6231 VDPWR.n1053 VDPWR.n1052 2.1509
R6232 VDPWR.n1133 VDPWR.n1129 2.1509
R6233 VDPWR.n1797 VDPWR.n878 2.1509
R6234 VDPWR.n2121 VDPWR.n2120 2.1509
R6235 VDPWR.n2322 VDPWR.n2299 2.13383
R6236 VDPWR.n2445 VDPWR.n1838 2.13383
R6237 VDPWR.n2353 VDPWR.n2024 2.13383
R6238 VDPWR.n2015 VDPWR.n1891 2.13383
R6239 VDPWR.n1492 VDPWR.n1488 2.13383
R6240 VDPWR.n783 VDPWR.n782 2.13383
R6241 VDPWR.n1320 VDPWR.n1319 2.13383
R6242 VDPWR.n993 VDPWR.n992 2.13383
R6243 VDPWR.n1134 VDPWR.n1100 2.13383
R6244 VDPWR.n1384 VDPWR.n1383 2.08643
R6245 VDPWR.n2501 VDPWR.n787 2.08643
R6246 VDPWR.n2477 VDPWR.n818 2.08643
R6247 VDPWR.n1604 VDPWR.n1222 2.08643
R6248 VDPWR.n1734 VDPWR.n886 2.08643
R6249 VDPWR.n2443 VDPWR.n1840 2.08643
R6250 VDPWR.n2015 VDPWR.n2014 1.9461
R6251 VDPWR.n1523 VDPWR.n1492 1.9461
R6252 VDPWR.n1390 VDPWR.n1320 1.9461
R6253 VDPWR.n2547 VDPWR.n783 1.9461
R6254 VDPWR.n2354 VDPWR.n2353 1.9461
R6255 VDPWR.n992 VDPWR.n991 1.9461
R6256 VDPWR.n1217 VDPWR.n1100 1.9461
R6257 VDPWR.n2446 VDPWR.n2445 1.9461
R6258 VDPWR.n2323 VDPWR.n2322 1.9461
R6259 VDPWR.n280 VDPWR.n279 1.71099
R6260 VDPWR.n281 VDPWR.n273 1.71099
R6261 VDPWR.n339 VDPWR.n338 1.71099
R6262 VDPWR.n340 VDPWR.n332 1.71099
R6263 VDPWR.n2750 VDPWR.n2749 1.70307
R6264 VDPWR.n2752 VDPWR.n2751 1.70307
R6265 VDPWR.n2756 VDPWR.n1 1.70307
R6266 VDPWR.n2749 VDPWR.n0 1.70307
R6267 VDPWR.n2381 VDPWR.n2380 1.52512
R6268 VDPWR.n2351 VDPWR.n2349 1.52512
R6269 VDPWR.n2320 VDPWR.n2319 1.52512
R6270 VDPWR.n1406 VDPWR.n1405 1.42272
R6271 VDPWR.n1074 VDPWR.n1073 1.42272
R6272 VDPWR.n1682 VDPWR.n1078 1.42272
R6273 VDPWR.n2384 VDPWR.n51 1.28415
R6274 VDPWR.n2620 VDPWR.n79 1.20883
R6275 VDPWR.n2620 VDPWR.n2619 1.14633
R6276 VDPWR.n1685 VDPWR.n37 1.11531
R6277 VDPWR.n694 VDPWR.n610 1.1097
R6278 VDPWR.n1985 VDPWR.n1983 0.8197
R6279 VDPWR.n1984 VDPWR.n1906 0.8197
R6280 VDPWR.n1992 VDPWR.n1991 0.8197
R6281 VDPWR.n1908 VDPWR.n1907 0.8197
R6282 VDPWR.n2000 VDPWR.n1902 0.8197
R6283 VDPWR.n1999 VDPWR.n1900 0.8197
R6284 VDPWR.n1899 VDPWR.n1896 0.8197
R6285 VDPWR.n2008 VDPWR.n2007 0.8197
R6286 VDPWR.n1897 VDPWR.n1892 0.8197
R6287 VDPWR.n1582 VDPWR.n1580 0.8197
R6288 VDPWR.n1581 VDPWR.n1472 0.8197
R6289 VDPWR.n1471 VDPWR.n1468 0.8197
R6290 VDPWR.n1590 VDPWR.n1589 0.8197
R6291 VDPWR.n1503 VDPWR.n1469 0.8197
R6292 VDPWR.n1506 VDPWR.n1505 0.8197
R6293 VDPWR.n1511 VDPWR.n1502 0.8197
R6294 VDPWR.n1513 VDPWR.n1512 0.8197
R6295 VDPWR.n1524 VDPWR.n1490 0.8197
R6296 VDPWR.n1265 VDPWR.n1238 0.8197
R6297 VDPWR.n1264 VDPWR.n1241 0.8197
R6298 VDPWR.n1397 VDPWR.n1396 0.8197
R6299 VDPWR.n1324 VDPWR.n1242 0.8197
R6300 VDPWR.n1328 VDPWR.n1326 0.8197
R6301 VDPWR.n1330 VDPWR.n1329 0.8197
R6302 VDPWR.n1336 VDPWR.n1335 0.8197
R6303 VDPWR.n1332 VDPWR.n1331 0.8197
R6304 VDPWR.n1391 VDPWR.n1263 0.8197
R6305 VDPWR.n2554 VDPWR.n2553 0.8197
R6306 VDPWR.n2509 VDPWR.n709 0.8197
R6307 VDPWR.n2515 VDPWR.n2513 0.8197
R6308 VDPWR.n2519 VDPWR.n2516 0.8197
R6309 VDPWR.n2520 VDPWR.n2507 0.8197
R6310 VDPWR.n2525 VDPWR.n2524 0.8197
R6311 VDPWR.n2528 VDPWR.n2506 0.8197
R6312 VDPWR.n2530 VDPWR.n2529 0.8197
R6313 VDPWR.n2548 VDPWR.n730 0.8197
R6314 VDPWR.n2239 VDPWR.n2235 0.8197
R6315 VDPWR.n2238 VDPWR.n2137 0.8197
R6316 VDPWR.n2136 VDPWR.n2133 0.8197
R6317 VDPWR.n2247 VDPWR.n2246 0.8197
R6318 VDPWR.n2158 VDPWR.n2134 0.8197
R6319 VDPWR.n2160 VDPWR.n2159 0.8197
R6320 VDPWR.n2176 VDPWR.n2157 0.8197
R6321 VDPWR.n2175 VDPWR.n2154 0.8197
R6322 VDPWR.n2153 VDPWR.n2023 0.8197
R6323 VDPWR.n1052 VDPWR.n936 0.8197
R6324 VDPWR.n1048 VDPWR.n1047 0.8197
R6325 VDPWR.n967 VDPWR.n938 0.8197
R6326 VDPWR.n969 VDPWR.n968 0.8197
R6327 VDPWR.n976 VDPWR.n965 0.8197
R6328 VDPWR.n975 VDPWR.n962 0.8197
R6329 VDPWR.n961 VDPWR.n958 0.8197
R6330 VDPWR.n984 VDPWR.n983 0.8197
R6331 VDPWR.n956 VDPWR.n955 0.8197
R6332 VDPWR.n1188 VDPWR.n1129 0.8197
R6333 VDPWR.n1192 VDPWR.n1191 0.8197
R6334 VDPWR.n1127 VDPWR.n1126 0.8197
R6335 VDPWR.n1199 VDPWR.n1198 0.8197
R6336 VDPWR.n1202 VDPWR.n1125 0.8197
R6337 VDPWR.n1204 VDPWR.n1203 0.8197
R6338 VDPWR.n1211 VDPWR.n1122 0.8197
R6339 VDPWR.n1210 VDPWR.n1123 0.8197
R6340 VDPWR.n1216 VDPWR.n1102 0.8197
R6341 VDPWR.n1810 VDPWR.n878 0.8197
R6342 VDPWR.n1809 VDPWR.n876 0.8197
R6343 VDPWR.n875 VDPWR.n868 0.8197
R6344 VDPWR.n1818 VDPWR.n1817 0.8197
R6345 VDPWR.n873 VDPWR.n869 0.8197
R6346 VDPWR.n872 VDPWR.n871 0.8197
R6347 VDPWR.n1831 VDPWR.n860 0.8197
R6348 VDPWR.n1830 VDPWR.n858 0.8197
R6349 VDPWR.n857 VDPWR.n854 0.8197
R6350 VDPWR.n2270 VDPWR.n2121 0.8197
R6351 VDPWR.n2269 VDPWR.n2056 0.8197
R6352 VDPWR.n2055 VDPWR.n2047 0.8197
R6353 VDPWR.n2278 VDPWR.n2277 0.8197
R6354 VDPWR.n2053 VDPWR.n2048 0.8197
R6355 VDPWR.n2052 VDPWR.n2050 0.8197
R6356 VDPWR.n2292 VDPWR.n2037 0.8197
R6357 VDPWR.n2291 VDPWR.n2035 0.8197
R6358 VDPWR.n2034 VDPWR.n2031 0.8197
R6359 VDPWR.n357 VDPWR.n261 0.703977
R6360 VDPWR.n2610 VDPWR.n2593 0.65675
R6361 VDPWR.n307 VDPWR.n303 0.576295
R6362 VDPWR.n2570 VDPWR.n2569 0.542167
R6363 VDPWR.n124 VDPWR.n122 0.492597
R6364 VDPWR.n474 VDPWR.n473 0.206967
R6365 VDPWR.n2745 VDPWR.n3 0.206942
R6366 VDPWR.n385 VDPWR.n2 0.206942
R6367 VDPWR.n693 VDPWR.n611 0.199496
R6368 VDPWR.n502 VDPWR.n498 0.196005
R6369 VDPWR.n2565 VDPWR.n2564 0.188
R6370 VDPWR.n2568 VDPWR.n699 0.188
R6371 VDPWR.n2619 VDPWR.n2618 0.188
R6372 VDPWR.n609 VDPWR.n608 0.185879
R6373 VDPWR.n2678 VDPWR.n2653 0.15675
R6374 VDPWR.n2679 VDPWR.n2678 0.15675
R6375 VDPWR.n2682 VDPWR.n2679 0.15675
R6376 VDPWR.n2686 VDPWR.n2651 0.15675
R6377 VDPWR.n2687 VDPWR.n2686 0.15675
R6378 VDPWR.n2690 VDPWR.n2687 0.15675
R6379 VDPWR.n2694 VDPWR.n2649 0.15675
R6380 VDPWR.n2695 VDPWR.n2694 0.15675
R6381 VDPWR.n2698 VDPWR.n2695 0.15675
R6382 VDPWR.n2702 VDPWR.n2647 0.15675
R6383 VDPWR.n2703 VDPWR.n2702 0.15675
R6384 VDPWR.n2706 VDPWR.n2703 0.15675
R6385 VDPWR.n2710 VDPWR.n2645 0.15675
R6386 VDPWR.n633 VDPWR.n3 0.15675
R6387 VDPWR.n634 VDPWR.n633 0.15675
R6388 VDPWR.n635 VDPWR.n634 0.15675
R6389 VDPWR.n635 VDPWR.n630 0.15675
R6390 VDPWR.n639 VDPWR.n630 0.15675
R6391 VDPWR.n640 VDPWR.n639 0.15675
R6392 VDPWR.n641 VDPWR.n640 0.15675
R6393 VDPWR.n641 VDPWR.n627 0.15675
R6394 VDPWR.n627 VDPWR.n625 0.15675
R6395 VDPWR.n646 VDPWR.n625 0.15675
R6396 VDPWR.n647 VDPWR.n646 0.15675
R6397 VDPWR.n648 VDPWR.n647 0.15675
R6398 VDPWR.n648 VDPWR.n623 0.15675
R6399 VDPWR.n652 VDPWR.n623 0.15675
R6400 VDPWR.n653 VDPWR.n652 0.15675
R6401 VDPWR.n654 VDPWR.n653 0.15675
R6402 VDPWR.n654 VDPWR.n621 0.15675
R6403 VDPWR.n658 VDPWR.n621 0.15675
R6404 VDPWR.n659 VDPWR.n658 0.15675
R6405 VDPWR.n660 VDPWR.n659 0.15675
R6406 VDPWR.n660 VDPWR.n619 0.15675
R6407 VDPWR.n665 VDPWR.n619 0.15675
R6408 VDPWR.n666 VDPWR.n665 0.15675
R6409 VDPWR.n667 VDPWR.n666 0.15675
R6410 VDPWR.n667 VDPWR.n617 0.15675
R6411 VDPWR.n671 VDPWR.n617 0.15675
R6412 VDPWR.n672 VDPWR.n671 0.15675
R6413 VDPWR.n673 VDPWR.n672 0.15675
R6414 VDPWR.n673 VDPWR.n615 0.15675
R6415 VDPWR.n678 VDPWR.n615 0.15675
R6416 VDPWR.n679 VDPWR.n678 0.15675
R6417 VDPWR.n680 VDPWR.n679 0.15675
R6418 VDPWR.n680 VDPWR.n613 0.15675
R6419 VDPWR.n685 VDPWR.n613 0.15675
R6420 VDPWR.n686 VDPWR.n685 0.15675
R6421 VDPWR.n687 VDPWR.n686 0.15675
R6422 VDPWR.n687 VDPWR.n611 0.15675
R6423 VDPWR.n496 VDPWR.n245 0.15675
R6424 VDPWR.n492 VDPWR.n245 0.15675
R6425 VDPWR.n492 VDPWR.n491 0.15675
R6426 VDPWR.n491 VDPWR.n490 0.15675
R6427 VDPWR.n490 VDPWR.n248 0.15675
R6428 VDPWR.n486 VDPWR.n248 0.15675
R6429 VDPWR.n486 VDPWR.n485 0.15675
R6430 VDPWR.n485 VDPWR.n484 0.15675
R6431 VDPWR.n484 VDPWR.n250 0.15675
R6432 VDPWR.n480 VDPWR.n250 0.15675
R6433 VDPWR.n480 VDPWR.n479 0.15675
R6434 VDPWR.n479 VDPWR.n478 0.15675
R6435 VDPWR.n478 VDPWR.n253 0.15675
R6436 VDPWR.n474 VDPWR.n253 0.15675
R6437 VDPWR.n129 VDPWR.n122 0.15675
R6438 VDPWR.n130 VDPWR.n129 0.15675
R6439 VDPWR.n131 VDPWR.n130 0.15675
R6440 VDPWR.n131 VDPWR.n120 0.15675
R6441 VDPWR.n135 VDPWR.n120 0.15675
R6442 VDPWR.n136 VDPWR.n135 0.15675
R6443 VDPWR.n137 VDPWR.n136 0.15675
R6444 VDPWR.n137 VDPWR.n118 0.15675
R6445 VDPWR.n142 VDPWR.n118 0.15675
R6446 VDPWR.n143 VDPWR.n142 0.15675
R6447 VDPWR.n143 VDPWR.n115 0.15675
R6448 VDPWR.n147 VDPWR.n115 0.15675
R6449 VDPWR.n148 VDPWR.n147 0.15675
R6450 VDPWR.n149 VDPWR.n148 0.15675
R6451 VDPWR.n149 VDPWR.n112 0.15675
R6452 VDPWR.n153 VDPWR.n112 0.15675
R6453 VDPWR.n154 VDPWR.n153 0.15675
R6454 VDPWR.n155 VDPWR.n154 0.15675
R6455 VDPWR.n155 VDPWR.n110 0.15675
R6456 VDPWR.n159 VDPWR.n110 0.15675
R6457 VDPWR.n160 VDPWR.n159 0.15675
R6458 VDPWR.n160 VDPWR.n107 0.15675
R6459 VDPWR.n165 VDPWR.n107 0.15675
R6460 VDPWR.n166 VDPWR.n165 0.15675
R6461 VDPWR.n167 VDPWR.n166 0.15675
R6462 VDPWR.n167 VDPWR.n105 0.15675
R6463 VDPWR.n173 VDPWR.n105 0.15675
R6464 VDPWR.n174 VDPWR.n173 0.15675
R6465 VDPWR.n175 VDPWR.n174 0.15675
R6466 VDPWR.n175 VDPWR.n103 0.15675
R6467 VDPWR.n179 VDPWR.n103 0.15675
R6468 VDPWR.n180 VDPWR.n179 0.15675
R6469 VDPWR.n181 VDPWR.n180 0.15675
R6470 VDPWR.n181 VDPWR.n101 0.15675
R6471 VDPWR.n185 VDPWR.n101 0.15675
R6472 VDPWR.n186 VDPWR.n185 0.15675
R6473 VDPWR.n186 VDPWR.n99 0.15675
R6474 VDPWR.n191 VDPWR.n99 0.15675
R6475 VDPWR.n192 VDPWR.n191 0.15675
R6476 VDPWR.n193 VDPWR.n192 0.15675
R6477 VDPWR.n193 VDPWR.n97 0.15675
R6478 VDPWR.n199 VDPWR.n97 0.15675
R6479 VDPWR.n200 VDPWR.n199 0.15675
R6480 VDPWR.n578 VDPWR.n200 0.15675
R6481 VDPWR.n578 VDPWR.n577 0.15675
R6482 VDPWR.n577 VDPWR.n576 0.15675
R6483 VDPWR.n576 VDPWR.n201 0.15675
R6484 VDPWR.n572 VDPWR.n201 0.15675
R6485 VDPWR.n572 VDPWR.n571 0.15675
R6486 VDPWR.n571 VDPWR.n570 0.15675
R6487 VDPWR.n570 VDPWR.n203 0.15675
R6488 VDPWR.n566 VDPWR.n203 0.15675
R6489 VDPWR.n566 VDPWR.n565 0.15675
R6490 VDPWR.n565 VDPWR.n207 0.15675
R6491 VDPWR.n561 VDPWR.n207 0.15675
R6492 VDPWR.n561 VDPWR.n560 0.15675
R6493 VDPWR.n560 VDPWR.n559 0.15675
R6494 VDPWR.n559 VDPWR.n209 0.15675
R6495 VDPWR.n555 VDPWR.n209 0.15675
R6496 VDPWR.n555 VDPWR.n554 0.15675
R6497 VDPWR.n554 VDPWR.n553 0.15675
R6498 VDPWR.n553 VDPWR.n212 0.15675
R6499 VDPWR.n214 VDPWR.n212 0.15675
R6500 VDPWR.n548 VDPWR.n214 0.15675
R6501 VDPWR.n548 VDPWR.n547 0.15675
R6502 VDPWR.n547 VDPWR.n546 0.15675
R6503 VDPWR.n546 VDPWR.n217 0.15675
R6504 VDPWR.n542 VDPWR.n217 0.15675
R6505 VDPWR.n542 VDPWR.n541 0.15675
R6506 VDPWR.n541 VDPWR.n540 0.15675
R6507 VDPWR.n540 VDPWR.n221 0.15675
R6508 VDPWR.n536 VDPWR.n221 0.15675
R6509 VDPWR.n536 VDPWR.n535 0.15675
R6510 VDPWR.n535 VDPWR.n534 0.15675
R6511 VDPWR.n534 VDPWR.n224 0.15675
R6512 VDPWR.n226 VDPWR.n224 0.15675
R6513 VDPWR.n529 VDPWR.n226 0.15675
R6514 VDPWR.n529 VDPWR.n528 0.15675
R6515 VDPWR.n528 VDPWR.n527 0.15675
R6516 VDPWR.n527 VDPWR.n229 0.15675
R6517 VDPWR.n523 VDPWR.n229 0.15675
R6518 VDPWR.n523 VDPWR.n522 0.15675
R6519 VDPWR.n522 VDPWR.n521 0.15675
R6520 VDPWR.n521 VDPWR.n233 0.15675
R6521 VDPWR.n517 VDPWR.n233 0.15675
R6522 VDPWR.n517 VDPWR.n516 0.15675
R6523 VDPWR.n516 VDPWR.n515 0.15675
R6524 VDPWR.n515 VDPWR.n236 0.15675
R6525 VDPWR.n239 VDPWR.n236 0.15675
R6526 VDPWR.n510 VDPWR.n239 0.15675
R6527 VDPWR.n510 VDPWR.n509 0.15675
R6528 VDPWR.n509 VDPWR.n508 0.15675
R6529 VDPWR.n508 VDPWR.n241 0.15675
R6530 VDPWR.n504 VDPWR.n241 0.15675
R6531 VDPWR.n504 VDPWR.n503 0.15675
R6532 VDPWR.n503 VDPWR.n502 0.15675
R6533 VDPWR.n308 VDPWR.n307 0.15675
R6534 VDPWR.n309 VDPWR.n308 0.15675
R6535 VDPWR.n309 VDPWR.n287 0.15675
R6536 VDPWR.n287 VDPWR.n286 0.15675
R6537 VDPWR.n314 VDPWR.n286 0.15675
R6538 VDPWR.n315 VDPWR.n314 0.15675
R6539 VDPWR.n316 VDPWR.n315 0.15675
R6540 VDPWR.n316 VDPWR.n271 0.15675
R6541 VDPWR.n320 VDPWR.n271 0.15675
R6542 VDPWR.n321 VDPWR.n320 0.15675
R6543 VDPWR.n322 VDPWR.n321 0.15675
R6544 VDPWR.n322 VDPWR.n268 0.15675
R6545 VDPWR.n326 VDPWR.n268 0.15675
R6546 VDPWR.n327 VDPWR.n326 0.15675
R6547 VDPWR.n328 VDPWR.n327 0.15675
R6548 VDPWR.n328 VDPWR.n265 0.15675
R6549 VDPWR.n343 VDPWR.n265 0.15675
R6550 VDPWR.n344 VDPWR.n343 0.15675
R6551 VDPWR.n345 VDPWR.n344 0.15675
R6552 VDPWR.n345 VDPWR.n263 0.15675
R6553 VDPWR.n350 VDPWR.n263 0.15675
R6554 VDPWR.n351 VDPWR.n350 0.15675
R6555 VDPWR.n352 VDPWR.n351 0.15675
R6556 VDPWR.n352 VDPWR.n261 0.15675
R6557 VDPWR.n385 VDPWR.n383 0.15675
R6558 VDPWR.n389 VDPWR.n383 0.15675
R6559 VDPWR.n390 VDPWR.n389 0.15675
R6560 VDPWR.n391 VDPWR.n390 0.15675
R6561 VDPWR.n391 VDPWR.n381 0.15675
R6562 VDPWR.n395 VDPWR.n381 0.15675
R6563 VDPWR.n396 VDPWR.n395 0.15675
R6564 VDPWR.n396 VDPWR.n378 0.15675
R6565 VDPWR.n401 VDPWR.n378 0.15675
R6566 VDPWR.n402 VDPWR.n401 0.15675
R6567 VDPWR.n403 VDPWR.n402 0.15675
R6568 VDPWR.n403 VDPWR.n376 0.15675
R6569 VDPWR.n407 VDPWR.n376 0.15675
R6570 VDPWR.n408 VDPWR.n407 0.15675
R6571 VDPWR.n409 VDPWR.n408 0.15675
R6572 VDPWR.n409 VDPWR.n374 0.15675
R6573 VDPWR.n413 VDPWR.n374 0.15675
R6574 VDPWR.n414 VDPWR.n413 0.15675
R6575 VDPWR.n415 VDPWR.n414 0.15675
R6576 VDPWR.n438 VDPWR.n415 0.15675
R6577 VDPWR.n438 VDPWR.n437 0.15675
R6578 VDPWR.n437 VDPWR.n436 0.15675
R6579 VDPWR.n436 VDPWR.n417 0.15675
R6580 VDPWR.n431 VDPWR.n417 0.15675
R6581 VDPWR.n431 VDPWR.n430 0.15675
R6582 VDPWR.n430 VDPWR.n429 0.15675
R6583 VDPWR.n429 VDPWR.n420 0.15675
R6584 VDPWR.n425 VDPWR.n420 0.15675
R6585 VDPWR.n425 VDPWR.n424 0.15675
R6586 VDPWR.n424 VDPWR.n91 0.15675
R6587 VDPWR.n91 VDPWR.n89 0.15675
R6588 VDPWR.n589 VDPWR.n89 0.15675
R6589 VDPWR.n590 VDPWR.n589 0.15675
R6590 VDPWR.n592 VDPWR.n590 0.15675
R6591 VDPWR.n596 VDPWR.n87 0.15675
R6592 VDPWR.n597 VDPWR.n596 0.15675
R6593 VDPWR.n598 VDPWR.n597 0.15675
R6594 VDPWR.n598 VDPWR.n84 0.15675
R6595 VDPWR.n602 VDPWR.n84 0.15675
R6596 VDPWR.n603 VDPWR.n602 0.15675
R6597 VDPWR.n604 VDPWR.n603 0.15675
R6598 VDPWR.n604 VDPWR.n82 0.15675
R6599 VDPWR.n608 VDPWR.n82 0.15675
R6600 VDPWR.n497 VDPWR.n496 0.141125
R6601 VDPWR.n2711 VDPWR.n2642 0.131895
R6602 VDPWR.n2562 VDPWR.n701 0.1255
R6603 VDPWR.n2540 VDPWR.n2539 0.1255
R6604 VDPWR.n2625 VDPWR.n2624 0.1255
R6605 VDPWR.n591 VDPWR.n87 0.109875
R6606 VDPWR.n2675 VDPWR.n2655 0.0966335
R6607 VDPWR.n2655 VDPWR.n2653 0.09425
R6608 VDPWR.n2681 VDPWR.n2651 0.09425
R6609 VDPWR.n2689 VDPWR.n2649 0.09425
R6610 VDPWR.n2697 VDPWR.n2647 0.09425
R6611 VDPWR.n2705 VDPWR.n2645 0.09425
R6612 VDPWR.n2682 VDPWR.n2681 0.063
R6613 VDPWR.n2690 VDPWR.n2689 0.063
R6614 VDPWR.n2698 VDPWR.n2697 0.063
R6615 VDPWR.n2706 VDPWR.n2705 0.063
R6616 VDPWR.n2711 VDPWR.n2710 0.063
R6617 VDPWR.n2563 VDPWR.n2562 0.0626438
R6618 VDPWR.n2540 VDPWR.n2537 0.0626438
R6619 VDPWR.n2626 VDPWR.n2625 0.0626438
R6620 VDPWR.n592 VDPWR.n591 0.047375
R6621 VDPWR.n497 VDPWR.n80 0.0430057
R6622 VDPWR.n2569 VDPWR.n696 0.0421667
R6623 VDPWR.n2565 VDPWR.n697 0.0217373
R6624 VDPWR.n2568 VDPWR.n698 0.0217373
R6625 VDPWR.n700 VDPWR.n697 0.0217373
R6626 VDPWR.n700 VDPWR.n698 0.0217373
R6627 VDPWR.n2592 VDPWR.n2591 0.0217373
R6628 VDPWR.n2590 VDPWR.n695 0.0217373
R6629 VDPWR.n2593 VDPWR.n2592 0.0217373
R6630 VDPWR.n2567 VDPWR.n2566 0.0217373
R6631 VDPWR.n2590 VDPWR.n2589 0.0217373
R6632 VDPWR.n2566 VDPWR.n696 0.0217373
R6633 VDPWR.n2591 VDPWR.n2571 0.0217373
R6634 VDPWR.n2588 VDPWR.n2571 0.0217373
R6635 VDPWR.n2589 VDPWR.n2570 0.0217373
R6636 VDPWR.n2755 VDPWR.n2749 0.01225
R6637 VDPWR.n2753 VDPWR.n2749 0.01225
R6638 VDPWR.n2751 VDPWR.n1 0.0068649
R6639 VDPWR.n2754 VDPWR.n2750 0.0068649
R6640 VDPWR.n2752 VDPWR.n2747 0.0068649
R6641 VDPWR.n2756 VDPWR.n0 0.0068649
R6642 VDPWR.n2750 VDPWR.n2748 0.0068649
R6643 VDPWR.n2754 VDPWR.n2752 0.0068649
R6644 VDPWR.n2747 VDPWR.n0 0.0068649
R6645 VDPWR.n2753 VDPWR.n1 0.0068649
R6646 a_18180_33430.n0 a_18180_33430.n4 199.935
R6647 a_18180_33430.n0 a_18180_33430.n1 199.53
R6648 a_18180_33430.n0 a_18180_33430.n2 199.53
R6649 a_18180_33430.n0 a_18180_33430.n3 199.53
R6650 a_18180_33430.n5 a_18180_33430.n0 199.53
R6651 a_18180_33430.n0 a_18180_33430.t8 98.9938
R6652 a_18180_33430.n1 a_18180_33430.t7 48.0005
R6653 a_18180_33430.n1 a_18180_33430.t3 48.0005
R6654 a_18180_33430.n2 a_18180_33430.t10 48.0005
R6655 a_18180_33430.n2 a_18180_33430.t2 48.0005
R6656 a_18180_33430.n3 a_18180_33430.t5 48.0005
R6657 a_18180_33430.n3 a_18180_33430.t4 48.0005
R6658 a_18180_33430.n4 a_18180_33430.t6 48.0005
R6659 a_18180_33430.n4 a_18180_33430.t1 48.0005
R6660 a_18180_33430.t0 a_18180_33430.n5 48.0005
R6661 a_18180_33430.n5 a_18180_33430.t9 48.0005
R6662 a_25860_20180.n1 a_25860_20180.t3 600.206
R6663 a_25860_20180.t0 a_25860_20180.n5 576.192
R6664 a_25860_20180.n2 a_25860_20180.n1 568.072
R6665 a_25860_20180.n4 a_25860_20180.n2 392.486
R6666 a_25860_20180.n0 a_25860_20180.t2 289.791
R6667 a_25860_20180.n5 a_25860_20180.n4 168.067
R6668 a_25860_20180.n3 a_25860_20180.n0 97.9242
R6669 a_25860_20180.n4 a_25860_20180.n3 37.7572
R6670 a_25860_20180.n2 a_25860_20180.t4 32.1338
R6671 a_25860_20180.n1 a_25860_20180.t5 32.1338
R6672 a_25860_20180.n3 a_25860_20180.t1 32.1338
R6673 a_25860_20180.n5 a_25860_20180.n0 28.3357
R6674 a_26640_21760.t0 a_26640_21760.n0 421.027
R6675 a_26640_21760.n0 a_26640_21760.t2 348.81
R6676 a_26640_21760.n0 a_26640_21760.t1 316.159
R6677 a_24280_30060.t1 a_24280_30060.n2 500.086
R6678 a_24280_30060.n0 a_24280_30060.t2 490.034
R6679 a_24280_30060.t1 a_24280_30060.n2 461.389
R6680 a_24280_30060.n1 a_24280_30060.n0 449.233
R6681 a_24280_30060.n0 a_24280_30060.t3 345.433
R6682 a_24280_30060.n1 a_24280_30060.t0 177.577
R6683 a_24280_30060.n2 a_24280_30060.n1 48.3899
R6684 a_23100_30460.n1 a_23100_30460.t2 586.433
R6685 a_23100_30460.n2 a_23100_30460.n1 456.351
R6686 a_23100_30460.n0 a_23100_30460.t4 441.834
R6687 a_23100_30460.n0 a_23100_30460.t5 393.634
R6688 a_23100_30460.n3 a_23100_30460.n2 328.733
R6689 a_23100_30460.t0 a_23100_30460.n3 288.37
R6690 a_23100_30460.n1 a_23100_30460.t3 249.034
R6691 a_23100_30460.n3 a_23100_30460.t1 177.577
R6692 a_23100_30460.n2 a_23100_30460.n0 152.633
R6693 a_14730_30630.n4 a_14730_30630.n3 314.526
R6694 a_14730_30630.n5 a_14730_30630.t12 287.764
R6695 a_14730_30630.n6 a_14730_30630.t10 287.764
R6696 a_14730_30630.n5 a_14730_30630.t8 287.591
R6697 a_14730_30630.n7 a_14730_30630.t11 287.012
R6698 a_14730_30630.n8 a_14730_30630.t9 287.012
R6699 a_14730_30630.t0 a_14730_30630.n10 158.046
R6700 a_14730_30630.n2 a_14730_30630.n0 107.079
R6701 a_14730_30630.n2 a_14730_30630.n1 104.828
R6702 a_14730_30630.n10 a_14730_30630.t7 47.7913
R6703 a_14730_30630.n3 a_14730_30630.t1 39.4005
R6704 a_14730_30630.n3 a_14730_30630.t2 39.4005
R6705 a_14730_30630.n0 a_14730_30630.t6 13.1338
R6706 a_14730_30630.n0 a_14730_30630.t5 13.1338
R6707 a_14730_30630.n1 a_14730_30630.t3 13.1338
R6708 a_14730_30630.n1 a_14730_30630.t4 13.1338
R6709 a_14730_30630.n10 a_14730_30630.n9 13.0943
R6710 a_14730_30630.n9 a_14730_30630.n4 10.7505
R6711 a_14730_30630.n9 a_14730_30630.n8 6.78086
R6712 a_14730_30630.n4 a_14730_30630.n2 2.0005
R6713 a_14730_30630.n7 a_14730_30630.n6 0.579071
R6714 a_14730_30630.n8 a_14730_30630.n7 0.282643
R6715 a_14730_30630.n6 a_14730_30630.n5 0.2755
R6716 a_19910_25340.n4 a_19910_25340.n0 427.647
R6717 a_19910_25340.n1 a_19910_25340.t7 297.233
R6718 a_19910_25340.n5 a_19910_25340.n4 210.601
R6719 a_19910_25340.n3 a_19910_25340.t4 174.056
R6720 a_19910_25340.n2 a_19910_25340.n1 160.667
R6721 a_19910_25340.n4 a_19910_25340.n3 152
R6722 a_19910_25340.n1 a_19910_25340.t6 136.567
R6723 a_19910_25340.n2 a_19910_25340.t2 136.567
R6724 a_19910_25340.n5 a_19910_25340.t5 60.0005
R6725 a_19910_25340.t3 a_19910_25340.n5 60.0005
R6726 a_19910_25340.n0 a_19910_25340.t1 49.2505
R6727 a_19910_25340.n0 a_19910_25340.t0 49.2505
R6728 a_19910_25340.n3 a_19910_25340.n2 37.4894
R6729 a_19910_24200.n1 a_19910_24200.t6 377.567
R6730 a_19910_24200.n0 a_19910_24200.t8 297.233
R6731 a_19910_24200.n2 a_19910_24200.n1 233.476
R6732 a_19910_24200.n1 a_19910_24200.t7 216.9
R6733 a_19910_24200.n2 a_19910_24200.n0 213.998
R6734 a_19910_24200.n7 a_19910_24200.n6 205.862
R6735 a_19910_24200.n4 a_19910_24200.n3 178.903
R6736 a_19910_24200.n6 a_19910_24200.n5 178.901
R6737 a_19910_24200.n0 a_19910_24200.t9 136.567
R6738 a_19910_24200.n4 a_19910_24200.n2 66.8859
R6739 a_19910_24200.n6 a_19910_24200.n4 57.6005
R6740 a_19910_24200.n5 a_19910_24200.t3 24.6255
R6741 a_19910_24200.n5 a_19910_24200.t0 24.6255
R6742 a_19910_24200.n3 a_19910_24200.t5 24.6255
R6743 a_19910_24200.n3 a_19910_24200.t1 24.6255
R6744 a_19910_24200.t2 a_19910_24200.n7 15.0005
R6745 a_19910_24200.n7 a_19910_24200.t4 15.0005
R6746 a_19040_22530.t0 a_19040_22530.n6 1128.89
R6747 a_19040_22530.n3 a_19040_22530.n2 459.132
R6748 a_19040_22530.n2 a_19040_22530.n0 386.048
R6749 a_19040_22530.n2 a_19040_22530.n1 265
R6750 a_19040_22530.n3 a_19040_22530.t7 232.968
R6751 a_19040_22530.n4 a_19040_22530.t8 232.968
R6752 a_19040_22530.n5 a_19040_22530.t5 232.968
R6753 a_19040_22530.n6 a_19040_22530.t6 232.968
R6754 a_19040_22530.n4 a_19040_22530.n3 160.667
R6755 a_19040_22530.n5 a_19040_22530.n4 160.667
R6756 a_19040_22530.n6 a_19040_22530.n5 160.667
R6757 a_19040_22530.n1 a_19040_22530.t2 60.0005
R6758 a_19040_22530.n1 a_19040_22530.t1 60.0005
R6759 a_19040_22530.n0 a_19040_22530.t4 49.2505
R6760 a_19040_22530.n0 a_19040_22530.t3 49.2505
R6761 a_20480_25210.n5 a_20480_25210.n3 522.322
R6762 a_20480_25210.n11 a_20480_25210.t6 384.967
R6763 a_20480_25210.n0 a_20480_25210.t3 384.967
R6764 a_20480_25210.n0 a_20480_25210.t5 376.56
R6765 a_20480_25210.t7 a_20480_25210.n11 376.56
R6766 a_20480_25210.n8 a_20480_25210.n7 322.046
R6767 a_20480_25210.n10 a_20480_25210.n9 322.046
R6768 a_20480_25210.n2 a_20480_25210.n1 320.902
R6769 a_20480_25210.n5 a_20480_25210.n4 160.721
R6770 a_20480_25210.n10 a_20480_25210.n8 70.4005
R6771 a_20480_25210.n1 a_20480_25210.t9 49.2505
R6772 a_20480_25210.n1 a_20480_25210.t4 49.2505
R6773 a_20480_25210.n7 a_20480_25210.t0 49.2505
R6774 a_20480_25210.n7 a_20480_25210.t10 49.2505
R6775 a_20480_25210.n9 a_20480_25210.t8 49.2505
R6776 a_20480_25210.n9 a_20480_25210.t1 49.2505
R6777 a_20480_25210.n6 a_20480_25210.n5 37.763
R6778 a_20480_25210.n6 a_20480_25210.n2 36.2672
R6779 a_20480_25210.n4 a_20480_25210.t12 19.7005
R6780 a_20480_25210.n4 a_20480_25210.t2 19.7005
R6781 a_20480_25210.n3 a_20480_25210.t11 19.7005
R6782 a_20480_25210.n3 a_20480_25210.t13 19.7005
R6783 a_20480_25210.n8 a_20480_25210.n6 17.0672
R6784 a_20480_25210.n2 a_20480_25210.n0 9.6005
R6785 a_20480_25210.n11 a_20480_25210.n10 9.6005
R6786 w_20440_23530.n79 w_20440_23530.n78 585
R6787 w_20440_23530.n90 w_20440_23530.n89 585
R6788 w_20440_23530.n19 w_20440_23530.t50 384.967
R6789 w_20440_23530.n52 w_20440_23530.t54 384.967
R6790 w_20440_23530.n47 w_20440_23530.t46 384.967
R6791 w_20440_23530.n66 w_20440_23530.t38 384.967
R6792 w_20440_23530.n78 w_20440_23530.t58 374.878
R6793 w_20440_23530.n31 w_20440_23530.t42 352.834
R6794 w_20440_23530.n16 w_20440_23530.t48 341.752
R6795 w_20440_23530.n17 w_20440_23530.t57 341.752
R6796 w_20440_23530.n67 w_20440_23530.t41 341.752
R6797 w_20440_23530.n18 w_20440_23530.t52 341.752
R6798 w_20440_23530.n63 w_20440_23530.n62 322.046
R6799 w_20440_23530.n49 w_20440_23530.n48 322.046
R6800 w_20440_23530.n54 w_20440_23530.n50 322.046
R6801 w_20440_23530.n53 w_20440_23530.n51 322.046
R6802 w_20440_23530.n65 w_20440_23530.n64 322.046
R6803 w_20440_23530.n21 w_20440_23530.n20 322.046
R6804 w_20440_23530.t39 w_20440_23530.n67 304.659
R6805 w_20440_23530.n79 w_20440_23530.n73 290.733
R6806 w_20440_23530.n80 w_20440_23530.n79 290.733
R6807 w_20440_23530.n90 w_20440_23530.n9 290.733
R6808 w_20440_23530.n90 w_20440_23530.n10 290.733
R6809 w_20440_23530.n89 w_20440_23530.n11 230.308
R6810 w_20440_23530.n78 w_20440_23530.n69 230.308
R6811 w_20440_23530.n30 w_20440_23530.n15 230.308
R6812 w_20440_23530.n81 w_20440_23530.n80 188.536
R6813 w_20440_23530.n83 w_20440_23530.n17 185.001
R6814 w_20440_23530.n84 w_20440_23530.n16 185.001
R6815 w_20440_23530.n68 w_20440_23530.n18 185.001
R6816 w_20440_23530.n77 w_20440_23530.n76 185
R6817 w_20440_23530.n75 w_20440_23530.n74 185
R6818 w_20440_23530.n72 w_20440_23530.n71 185
R6819 w_20440_23530.n82 w_20440_23530.n81 185
R6820 w_20440_23530.n88 w_20440_23530.n87 185
R6821 w_20440_23530.n86 w_20440_23530.n14 185
R6822 w_20440_23530.n86 w_20440_23530.n85 185
R6823 w_20440_23530.n13 w_20440_23530.n12 185
R6824 w_20440_23530.t18 w_20440_23530.t14 145.038
R6825 w_20440_23530.n87 w_20440_23530.n86 120.001
R6826 w_20440_23530.n86 w_20440_23530.n12 120.001
R6827 w_20440_23530.n81 w_20440_23530.n71 120.001
R6828 w_20440_23530.n76 w_20440_23530.n75 120.001
R6829 w_20440_23530.n1 w_20440_23530.n32 119.737
R6830 w_20440_23530.n4 w_20440_23530.n29 119.737
R6831 w_20440_23530.n6 w_20440_23530.n27 119.737
R6832 w_20440_23530.n8 w_20440_23530.n25 119.737
R6833 w_20440_23530.n60 w_20440_23530.n23 119.737
R6834 w_20440_23530.n68 w_20440_23530.t51 119.656
R6835 w_20440_23530.n83 w_20440_23530.n82 108.779
R6836 w_20440_23530.t5 w_20440_23530.t4 94.2753
R6837 w_20440_23530.t28 w_20440_23530.t26 94.2753
R6838 w_20440_23530.n84 w_20440_23530.t16 94.2753
R6839 w_20440_23530.t47 w_20440_23530.t8 94.2753
R6840 w_20440_23530.t24 w_20440_23530.t0 94.2753
R6841 w_20440_23530.t51 w_20440_23530.t10 94.2753
R6842 w_20440_23530.t10 w_20440_23530.t6 94.2753
R6843 w_20440_23530.t6 w_20440_23530.t20 94.2753
R6844 w_20440_23530.t20 w_20440_23530.t22 94.2753
R6845 w_20440_23530.t22 w_20440_23530.t39 94.2753
R6846 w_20440_23530.t29 w_20440_23530.t12 83.3974
R6847 w_20440_23530.t55 w_20440_23530.t59 83.3974
R6848 w_20440_23530.t27 w_20440_23530.t43 76.1455
R6849 w_20440_23530.t30 w_20440_23530.t32 76.1455
R6850 w_20440_23530.n63 w_20440_23530.n61 75.7203
R6851 w_20440_23530.n54 w_20440_23530.n49 70.4005
R6852 w_20440_23530.n54 w_20440_23530.n53 70.4005
R6853 w_20440_23530.n63 w_20440_23530.n21 70.4005
R6854 w_20440_23530.n65 w_20440_23530.n63 70.4005
R6855 w_20440_23530.n82 w_20440_23530.n69 69.8479
R6856 w_20440_23530.n82 w_20440_23530.n70 69.8479
R6857 w_20440_23530.n85 w_20440_23530.n11 69.8479
R6858 w_20440_23530.n85 w_20440_23530.n15 69.8479
R6859 w_20440_23530.n85 w_20440_23530.t27 68.8936
R6860 w_20440_23530.t2 w_20440_23530.t30 68.8936
R6861 w_20440_23530.t34 w_20440_23530.t29 61.6417
R6862 w_20440_23530.t36 w_20440_23530.t55 61.6417
R6863 w_20440_23530.n55 w_20440_23530.n54 54.4005
R6864 w_20440_23530.t14 w_20440_23530.n84 50.7639
R6865 w_20440_23530.n62 w_20440_23530.t7 49.2505
R6866 w_20440_23530.n62 w_20440_23530.t21 49.2505
R6867 w_20440_23530.n48 w_20440_23530.t49 49.2505
R6868 w_20440_23530.n48 w_20440_23530.t9 49.2505
R6869 w_20440_23530.n50 w_20440_23530.t31 49.2505
R6870 w_20440_23530.n50 w_20440_23530.t25 49.2505
R6871 w_20440_23530.n51 w_20440_23530.t1 49.2505
R6872 w_20440_23530.n51 w_20440_23530.t56 49.2505
R6873 w_20440_23530.n64 w_20440_23530.t23 49.2505
R6874 w_20440_23530.n64 w_20440_23530.t40 49.2505
R6875 w_20440_23530.n20 w_20440_23530.t53 49.2505
R6876 w_20440_23530.n20 w_20440_23530.t11 49.2505
R6877 w_20440_23530.n15 w_20440_23530.n12 45.3071
R6878 w_20440_23530.n75 w_20440_23530.n70 45.3071
R6879 w_20440_23530.n76 w_20440_23530.n69 45.3071
R6880 w_20440_23530.n71 w_20440_23530.n70 45.3071
R6881 w_20440_23530.n87 w_20440_23530.n11 45.3071
R6882 w_20440_23530.t26 w_20440_23530.t18 39.886
R6883 w_20440_23530.n33 w_20440_23530.n2 39.4998
R6884 w_20440_23530.n61 w_20440_23530.n22 39.4988
R6885 w_20440_23530.t59 w_20440_23530.n83 36.26
R6886 w_20440_23530.t4 w_20440_23530.t34 32.6341
R6887 w_20440_23530.t0 w_20440_23530.t36 32.6341
R6888 w_20440_23530.n34 w_20440_23530.n33 32.0005
R6889 w_20440_23530.n34 w_20440_23530.n28 32.0005
R6890 w_20440_23530.n37 w_20440_23530.n28 32.0005
R6891 w_20440_23530.n38 w_20440_23530.n37 32.0005
R6892 w_20440_23530.n39 w_20440_23530.n38 32.0005
R6893 w_20440_23530.n39 w_20440_23530.n26 32.0005
R6894 w_20440_23530.n42 w_20440_23530.n26 32.0005
R6895 w_20440_23530.n43 w_20440_23530.n42 32.0005
R6896 w_20440_23530.n44 w_20440_23530.n43 32.0005
R6897 w_20440_23530.n44 w_20440_23530.n24 32.0005
R6898 w_20440_23530.n55 w_20440_23530.n24 32.0005
R6899 w_20440_23530.n57 w_20440_23530.n56 32.0005
R6900 w_20440_23530.n57 w_20440_23530.n22 32.0005
R6901 w_20440_23530.n47 w_20440_23530.n16 30.1875
R6902 w_20440_23530.n52 w_20440_23530.n17 30.1875
R6903 w_20440_23530.n67 w_20440_23530.n66 30.1875
R6904 w_20440_23530.n19 w_20440_23530.n18 30.1875
R6905 w_20440_23530.t16 w_20440_23530.t47 25.3822
R6906 w_20440_23530.t8 w_20440_23530.t2 25.3822
R6907 w_20440_23530.n31 w_20440_23530.n30 22.0449
R6908 w_20440_23530.n79 w_20440_23530.t61 19.7005
R6909 w_20440_23530.n32 w_20440_23530.t45 19.7005
R6910 w_20440_23530.n32 w_20440_23530.t35 19.7005
R6911 w_20440_23530.n29 w_20440_23530.t13 19.7005
R6912 w_20440_23530.n29 w_20440_23530.t19 19.7005
R6913 w_20440_23530.n27 w_20440_23530.t15 19.7005
R6914 w_20440_23530.n27 w_20440_23530.t17 19.7005
R6915 w_20440_23530.n25 w_20440_23530.t3 19.7005
R6916 w_20440_23530.n25 w_20440_23530.t33 19.7005
R6917 w_20440_23530.n23 w_20440_23530.t37 19.7005
R6918 w_20440_23530.n23 w_20440_23530.t60 19.7005
R6919 w_20440_23530.t44 w_20440_23530.n90 19.7005
R6920 w_20440_23530.n56 w_20440_23530.n55 19.2005
R6921 w_20440_23530.t43 w_20440_23530.t5 18.1303
R6922 w_20440_23530.t32 w_20440_23530.t24 18.1303
R6923 w_20440_23530.t12 w_20440_23530.t28 10.8784
R6924 w_20440_23530.n2 w_20440_23530.n31 9.95328
R6925 w_20440_23530.n49 w_20440_23530.n47 9.6005
R6926 w_20440_23530.n53 w_20440_23530.n52 9.6005
R6927 w_20440_23530.n66 w_20440_23530.n65 9.6005
R6928 w_20440_23530.n21 w_20440_23530.n19 9.6005
R6929 w_20440_23530.n59 w_20440_23530.n22 9.3005
R6930 w_20440_23530.n58 w_20440_23530.n57 9.3005
R6931 w_20440_23530.n56 w_20440_23530.n7 9.3005
R6932 w_20440_23530.n55 w_20440_23530.n8 9.3005
R6933 w_20440_23530.n46 w_20440_23530.n24 9.3005
R6934 w_20440_23530.n45 w_20440_23530.n44 9.3005
R6935 w_20440_23530.n43 w_20440_23530.n5 9.3005
R6936 w_20440_23530.n42 w_20440_23530.n6 9.3005
R6937 w_20440_23530.n41 w_20440_23530.n26 9.3005
R6938 w_20440_23530.n40 w_20440_23530.n39 9.3005
R6939 w_20440_23530.n38 w_20440_23530.n3 9.3005
R6940 w_20440_23530.n37 w_20440_23530.n4 9.3005
R6941 w_20440_23530.n36 w_20440_23530.n28 9.3005
R6942 w_20440_23530.n35 w_20440_23530.n34 9.3005
R6943 w_20440_23530.n33 w_20440_23530.n0 9.3005
R6944 w_20440_23530.n2 w_20440_23530.n1 0.0368314
R6945 w_20440_23530.n82 w_20440_23530.n68 7.25241
R6946 w_20440_23530.n74 w_20440_23530.n72 7.11161
R6947 w_20440_23530.n78 w_20440_23530.n77 7.11161
R6948 w_20440_23530.n89 w_20440_23530.n88 7.11161
R6949 w_20440_23530.n14 w_20440_23530.n13 7.11161
R6950 w_20440_23530.n74 w_20440_23530.n73 3.53508
R6951 w_20440_23530.n77 w_20440_23530.n73 3.53508
R6952 w_20440_23530.n80 w_20440_23530.n72 3.53508
R6953 w_20440_23530.n14 w_20440_23530.n10 3.53508
R6954 w_20440_23530.n30 w_20440_23530.n9 3.53508
R6955 w_20440_23530.n13 w_20440_23530.n9 3.53508
R6956 w_20440_23530.n88 w_20440_23530.n10 3.53508
R6957 w_20440_23530.n1 w_20440_23530.n0 0.15675
R6958 w_20440_23530.n35 w_20440_23530.n0 0.15675
R6959 w_20440_23530.n36 w_20440_23530.n35 0.15675
R6960 w_20440_23530.n4 w_20440_23530.n3 0.15675
R6961 w_20440_23530.n40 w_20440_23530.n3 0.15675
R6962 w_20440_23530.n41 w_20440_23530.n40 0.15675
R6963 w_20440_23530.n6 w_20440_23530.n5 0.15675
R6964 w_20440_23530.n45 w_20440_23530.n5 0.15675
R6965 w_20440_23530.n46 w_20440_23530.n45 0.15675
R6966 w_20440_23530.n8 w_20440_23530.n7 0.15675
R6967 w_20440_23530.n58 w_20440_23530.n7 0.15675
R6968 w_20440_23530.n59 w_20440_23530.n58 0.15675
R6969 w_20440_23530.n8 w_20440_23530.n46 0.15675
R6970 w_20440_23530.n6 w_20440_23530.n41 0.15675
R6971 w_20440_23530.n4 w_20440_23530.n36 0.15675
R6972 w_20440_23530.n61 w_20440_23530.n60 0.100307
R6973 w_20440_23530.n60 w_20440_23530.n59 0.09425
R6974 a_17884_25798.t8 a_17884_25798.n11 1456.66
R6975 a_17884_25798.n3 a_17884_25798.t10 377.567
R6976 a_17884_25798.n5 a_17884_25798.t11 377.567
R6977 a_17884_25798.n4 a_17884_25798.n3 257.067
R6978 a_17884_25798.n9 a_17884_25798.n8 257.067
R6979 a_17884_25798.n6 a_17884_25798.n5 257.067
R6980 a_17884_25798.n2 a_17884_25798.n1 159.12
R6981 a_17884_25798.n11 a_17884_25798.n0 154.321
R6982 a_17884_25798.n7 a_17884_25798.n2 153.601
R6983 a_17884_25798.n11 a_17884_25798.n10 152
R6984 a_17884_25798.n8 a_17884_25798.t0 120.501
R6985 a_17884_25798.n9 a_17884_25798.t6 120.501
R6986 a_17884_25798.n4 a_17884_25798.t2 120.501
R6987 a_17884_25798.n3 a_17884_25798.t12 120.501
R6988 a_17884_25798.n6 a_17884_25798.t4 120.501
R6989 a_17884_25798.n5 a_17884_25798.t9 120.501
R6990 a_17884_25798.n11 a_17884_25798.n2 108.8
R6991 a_17884_25798.n10 a_17884_25798.n4 85.6894
R6992 a_17884_25798.n10 a_17884_25798.n9 85.6894
R6993 a_17884_25798.n8 a_17884_25798.n7 85.6894
R6994 a_17884_25798.n7 a_17884_25798.n6 85.6894
R6995 a_17884_25798.n0 a_17884_25798.t3 19.7005
R6996 a_17884_25798.n0 a_17884_25798.t7 19.7005
R6997 a_17884_25798.n1 a_17884_25798.t1 19.7005
R6998 a_17884_25798.n1 a_17884_25798.t5 19.7005
R6999 a_26320_28790.n4 a_26320_28790.t0 782.52
R7000 a_26320_28790.t11 a_26320_28790.t2 514.134
R7001 a_26320_28790.t5 a_26320_28790.n5 377.567
R7002 a_26320_28790.n0 a_26320_28790.t3 377.567
R7003 a_26320_28790.n3 a_26320_28790.n2 321.334
R7004 a_26320_28790.n6 a_26320_28790.t5 318.702
R7005 a_26320_28790.n6 a_26320_28790.t11 307.909
R7006 a_26320_28790.n4 a_26320_28790.n3 275.341
R7007 a_26320_28790.n5 a_26320_28790.t7 265.101
R7008 a_26320_28790.t1 a_26320_28790.n7 233
R7009 a_26320_28790.n0 a_26320_28790.t8 168.701
R7010 a_26320_28790.n5 a_26320_28790.t6 136.567
R7011 a_26320_28790.n1 a_26320_28790.t4 136.567
R7012 a_26320_28790.n2 a_26320_28790.t9 136.567
R7013 a_26320_28790.n2 a_26320_28790.n1 128.534
R7014 a_26320_28790.n3 a_26320_28790.t10 126.927
R7015 a_26320_28790.n1 a_26320_28790.n0 48.2005
R7016 a_26320_28790.n7 a_26320_28790.n6 38.2642
R7017 a_26320_28790.n7 a_26320_28790.n4 26.4538
R7018 a_26420_30200.n0 a_26420_30200.t2 691.534
R7019 a_26420_30200.n1 a_26420_30200.t1 691.534
R7020 a_26420_30200.n0 a_26420_30200.t3 527.867
R7021 a_26420_30200.t0 a_26420_30200.n1 343.401
R7022 a_26420_30200.n1 a_26420_30200.n0 92.8005
R7023 a_13532_27710.t0 a_13532_27710.t16 170.145
R7024 a_13532_27710.t17 a_13532_27710.t10 0.1603
R7025 a_13532_27710.t11 a_13532_27710.t17 0.1603
R7026 a_13532_27710.t19 a_13532_27710.t11 0.1603
R7027 a_13532_27710.t3 a_13532_27710.t19 0.1603
R7028 a_13532_27710.t6 a_13532_27710.t3 0.1603
R7029 a_13532_27710.t4 a_13532_27710.t6 0.1603
R7030 a_13532_27710.t8 a_13532_27710.t4 0.1603
R7031 a_13532_27710.t14 a_13532_27710.t8 0.1603
R7032 a_13532_27710.t13 a_13532_27710.t20 0.1603
R7033 a_13532_27710.t7 a_13532_27710.t13 0.1603
R7034 a_13532_27710.t12 a_13532_27710.t7 0.1603
R7035 a_13532_27710.t5 a_13532_27710.t12 0.1603
R7036 a_13532_27710.t2 a_13532_27710.t5 0.1603
R7037 a_13532_27710.t18 a_13532_27710.t2 0.1603
R7038 a_13532_27710.t1 a_13532_27710.t18 0.1603
R7039 a_13532_27710.t16 a_13532_27710.t1 0.1603
R7040 a_13532_27710.t15 a_13532_27710.n0 0.159278
R7041 a_13532_27710.t20 a_13532_27710.t15 0.137822
R7042 a_13532_27710.n0 a_13532_27710.t14 0.1368
R7043 a_13532_27710.n0 a_13532_27710.t9 0.00152174
R7044 a_23100_27770.n0 a_23100_27770.t5 1180.9
R7045 a_23100_27770.n2 a_23100_27770.t3 522.168
R7046 a_23100_27770.t0 a_23100_27770.n4 458.818
R7047 a_23100_27770.t0 a_23100_27770.n4 429.281
R7048 a_23100_27770.n1 a_23100_27770.n0 417.733
R7049 a_23100_27770.n0 a_23100_27770.t2 232.968
R7050 a_23100_27770.n3 a_23100_27770.n2 228.8
R7051 a_23100_27770.n1 a_23100_27770.t4 217.905
R7052 a_23100_27770.n3 a_23100_27770.t1 164.775
R7053 a_23100_27770.n4 a_23100_27770.n3 60.248
R7054 a_23100_27770.n2 a_23100_27770.n1 15.063
R7055 a_23130_27670.t0 a_23130_27670.n8 458.818
R7056 a_23130_27670.t0 a_23130_27670.n8 429.281
R7057 a_23130_27670.n3 a_23130_27670.t6 326.658
R7058 a_23130_27670.t3 a_23130_27670.n5 297.233
R7059 a_23130_27670.n4 a_23130_27670.t7 297.233
R7060 a_23130_27670.n0 a_23130_27670.t2 294.829
R7061 a_23130_27670.n2 a_23130_27670.n1 257.067
R7062 a_23130_27670.n7 a_23130_27670.n6 242.494
R7063 a_23130_27670.n3 a_23130_27670.n2 226.942
R7064 a_23130_27670.n6 a_23130_27670.n1 226.942
R7065 a_23130_27670.n5 a_23130_27670.n4 216.9
R7066 a_23130_27670.n0 a_23130_27670.t1 151.976
R7067 a_23130_27670.n7 a_23130_27670.n0 137.601
R7068 a_23130_27670.n6 a_23130_27670.t3 92.3838
R7069 a_23130_27670.t7 a_23130_27670.n3 92.3838
R7070 a_23130_27670.n2 a_23130_27670.t5 80.3338
R7071 a_23130_27670.n4 a_23130_27670.t5 80.3338
R7072 a_23130_27670.t4 a_23130_27670.n1 80.3338
R7073 a_23130_27670.n5 a_23130_27670.t4 80.3338
R7074 a_23130_27670.n8 a_23130_27670.n7 34.648
R7075 a_19940_23090.n3 a_19940_23090.n1 418.048
R7076 a_19940_23090.n3 a_19940_23090.n2 360.447
R7077 a_19940_23090.n5 a_19940_23090.t3 328.175
R7078 a_19940_23090.n14 a_19940_23090.n0 306.601
R7079 a_19940_23090.t15 a_19940_23090.n9 297.233
R7080 a_19940_23090.n8 a_19940_23090.t14 297.233
R7081 a_19940_23090.t14 a_19940_23090.n7 297.233
R7082 a_19940_23090.n15 a_19940_23090.n14 249
R7083 a_19940_23090.n9 a_19940_23090.n8 216.9
R7084 a_19940_23090.n7 a_19940_23090.n6 216.9
R7085 a_19940_23090.n11 a_19940_23090.n10 210.351
R7086 a_19940_23090.n4 a_19940_23090.n3 208
R7087 a_19940_23090.n14 a_19940_23090.n13 208
R7088 a_19940_23090.n10 a_19940_23090.n6 180.75
R7089 a_19940_23090.n5 a_19940_23090.t1 118.627
R7090 a_19940_23090.n10 a_19940_23090.t15 92.3838
R7091 a_19940_23090.n7 a_19940_23090.t11 80.3338
R7092 a_19940_23090.n8 a_19940_23090.t11 80.3338
R7093 a_19940_23090.t10 a_19940_23090.n6 80.3338
R7094 a_19940_23090.n9 a_19940_23090.t10 80.3338
R7095 a_19940_23090.n13 a_19940_23090.t12 76.4829
R7096 a_19940_23090.n12 a_19940_23090.n11 73.0531
R7097 a_19940_23090.n4 a_19940_23090.t13 70.0829
R7098 a_19940_23090.n11 a_19940_23090.n5 62.8355
R7099 a_19940_23090.n0 a_19940_23090.t7 60.0005
R7100 a_19940_23090.n0 a_19940_23090.t6 60.0005
R7101 a_19940_23090.t9 a_19940_23090.n15 60.0005
R7102 a_19940_23090.n15 a_19940_23090.t8 60.0005
R7103 a_19940_23090.n13 a_19940_23090.n12 57.6005
R7104 a_19940_23090.n12 a_19940_23090.n4 54.4005
R7105 a_19940_23090.n1 a_19940_23090.t2 49.2505
R7106 a_19940_23090.n1 a_19940_23090.t0 49.2505
R7107 a_19940_23090.n2 a_19940_23090.t4 49.2505
R7108 a_19940_23090.n2 a_19940_23090.t5 49.2505
R7109 a_23100_30570.n4 a_23100_30570.n0 1295.28
R7110 a_23100_30570.n0 a_23100_30570.t3 586.433
R7111 a_23100_30570.n1 a_23100_30570.t5 388.813
R7112 a_23100_30570.n1 a_23100_30570.t6 356.68
R7113 a_23100_30570.n0 a_23100_30570.t4 249.034
R7114 a_23100_30570.n3 a_23100_30570.n1 225.601
R7115 a_23100_30570.t1 a_23100_30570.n4 221.411
R7116 a_23100_30570.n3 a_23100_30570.n2 163.677
R7117 a_23100_30570.n4 a_23100_30570.n3 84.24
R7118 a_23100_30570.n2 a_23100_30570.t2 24.0005
R7119 a_23100_30570.n2 a_23100_30570.t0 24.0005
R7120 a_23550_30490.t0 a_23550_30490.t1 39.4005
R7121 a_23100_30980.n0 a_23100_30980.t3 517.347
R7122 a_23100_30980.n2 a_23100_30980.n0 417.574
R7123 a_23100_30980.n2 a_23100_30980.n1 244.715
R7124 a_23100_30980.n0 a_23100_30980.t4 228.148
R7125 a_23100_30980.t1 a_23100_30980.n2 221.411
R7126 a_23100_30980.n1 a_23100_30980.t2 24.0005
R7127 a_23100_30980.n1 a_23100_30980.t0 24.0005
R7128 a_17884_25190.n2 a_17884_25190.t11 317.317
R7129 a_17884_25190.n9 a_17884_25190.t12 317.317
R7130 a_17884_25190.n3 a_17884_25190.n2 257.067
R7131 a_17884_25190.n10 a_17884_25190.n9 257.067
R7132 a_17884_25190.n8 a_17884_25190.n7 257.067
R7133 a_17884_25190.t8 a_17884_25190.n12 192.022
R7134 a_17884_25190.n6 a_17884_25190.n5 155.201
R7135 a_17884_25190.n12 a_17884_25190.n11 152
R7136 a_17884_25190.n1 a_17884_25190.n0 120.981
R7137 a_17884_25190.n5 a_17884_25190.n4 120.981
R7138 a_17884_25190.n5 a_17884_25190.n1 102.4
R7139 a_17884_25190.n6 a_17884_25190.n3 85.6894
R7140 a_17884_25190.n11 a_17884_25190.n10 85.6894
R7141 a_17884_25190.n11 a_17884_25190.n8 85.6894
R7142 a_17884_25190.n7 a_17884_25190.n6 85.6894
R7143 a_17884_25190.n3 a_17884_25190.t2 60.2505
R7144 a_17884_25190.n2 a_17884_25190.t9 60.2505
R7145 a_17884_25190.n7 a_17884_25190.t6 60.2505
R7146 a_17884_25190.n8 a_17884_25190.t0 60.2505
R7147 a_17884_25190.n10 a_17884_25190.t4 60.2505
R7148 a_17884_25190.n9 a_17884_25190.t10 60.2505
R7149 a_17884_25190.n0 a_17884_25190.t1 24.0005
R7150 a_17884_25190.n0 a_17884_25190.t5 24.0005
R7151 a_17884_25190.n4 a_17884_25190.t3 24.0005
R7152 a_17884_25190.n4 a_17884_25190.t7 24.0005
R7153 a_17884_25190.n12 a_17884_25190.n1 3.2005
R7154 a_19250_24340.n6 a_19250_24340.n4 482.582
R7155 a_19250_24340.n10 a_19250_24340.t5 304.634
R7156 a_19250_24340.n0 a_19250_24340.t2 304.634
R7157 a_19250_24340.n0 a_19250_24340.t4 276.289
R7158 a_19250_24340.t6 a_19250_24340.n10 276.289
R7159 a_19250_24340.n2 a_19250_24340.n1 210.601
R7160 a_19250_24340.n9 a_19250_24340.n8 210.601
R7161 a_19250_24340.n7 a_19250_24340.n3 207.4
R7162 a_19250_24340.n6 a_19250_24340.n5 120.981
R7163 a_19250_24340.n7 a_19250_24340.n2 64.0005
R7164 a_19250_24340.n9 a_19250_24340.n7 64.0005
R7165 a_19250_24340.n1 a_19250_24340.t8 60.0005
R7166 a_19250_24340.n1 a_19250_24340.t3 60.0005
R7167 a_19250_24340.n3 a_19250_24340.t0 60.0005
R7168 a_19250_24340.n3 a_19250_24340.t9 60.0005
R7169 a_19250_24340.n8 a_19250_24340.t7 60.0005
R7170 a_19250_24340.n8 a_19250_24340.t1 60.0005
R7171 a_19250_24340.n7 a_19250_24340.n6 47.363
R7172 a_19250_24340.n5 a_19250_24340.t12 24.0005
R7173 a_19250_24340.n5 a_19250_24340.t10 24.0005
R7174 a_19250_24340.n4 a_19250_24340.t11 24.0005
R7175 a_19250_24340.n4 a_19250_24340.t13 24.0005
R7176 a_19250_24340.n2 a_19250_24340.n0 9.6005
R7177 a_19250_24340.n10 a_19250_24340.n9 9.6005
R7178 a_19190_29290.n15 a_19190_29290.t18 310.488
R7179 a_19190_29290.n1 a_19190_29290.t21 310.488
R7180 a_19190_29290.n6 a_19190_29290.t17 310.488
R7181 a_19190_29290.n4 a_19190_29290.n0 297.433
R7182 a_19190_29290.n9 a_19190_29290.n5 297.433
R7183 a_19190_29290.n19 a_19190_29290.n18 297.433
R7184 a_19190_29290.n13 a_19190_29290.t15 248.133
R7185 a_19190_29290.n13 a_19190_29290.n12 199.383
R7186 a_19190_29290.n14 a_19190_29290.n11 194.883
R7187 a_19190_29290.n17 a_19190_29290.t10 184.097
R7188 a_19190_29290.n3 a_19190_29290.t6 184.097
R7189 a_19190_29290.n8 a_19190_29290.t4 184.097
R7190 a_19190_29290.n16 a_19190_29290.n15 167.094
R7191 a_19190_29290.n2 a_19190_29290.n1 167.094
R7192 a_19190_29290.n7 a_19190_29290.n6 167.094
R7193 a_19190_29290.n18 a_19190_29290.n17 161.3
R7194 a_19190_29290.n4 a_19190_29290.n3 161.3
R7195 a_19190_29290.n9 a_19190_29290.n8 161.3
R7196 a_19190_29290.n16 a_19190_29290.t8 120.501
R7197 a_19190_29290.n15 a_19190_29290.t19 120.501
R7198 a_19190_29290.n2 a_19190_29290.t0 120.501
R7199 a_19190_29290.n1 a_19190_29290.t20 120.501
R7200 a_19190_29290.n7 a_19190_29290.t2 120.501
R7201 a_19190_29290.n6 a_19190_29290.t22 120.501
R7202 a_19190_29290.n12 a_19190_29290.t12 48.0005
R7203 a_19190_29290.n12 a_19190_29290.t13 48.0005
R7204 a_19190_29290.n11 a_19190_29290.t14 48.0005
R7205 a_19190_29290.n11 a_19190_29290.t16 48.0005
R7206 a_19190_29290.n17 a_19190_29290.n16 40.7027
R7207 a_19190_29290.n3 a_19190_29290.n2 40.7027
R7208 a_19190_29290.n8 a_19190_29290.n7 40.7027
R7209 a_19190_29290.n0 a_19190_29290.t1 39.4005
R7210 a_19190_29290.n0 a_19190_29290.t7 39.4005
R7211 a_19190_29290.n5 a_19190_29290.t3 39.4005
R7212 a_19190_29290.n5 a_19190_29290.t5 39.4005
R7213 a_19190_29290.n19 a_19190_29290.t9 39.4005
R7214 a_19190_29290.t11 a_19190_29290.n19 39.4005
R7215 a_19190_29290.n10 a_19190_29290.n4 6.6255
R7216 a_19190_29290.n10 a_19190_29290.n9 6.6255
R7217 a_19190_29290.n14 a_19190_29290.n13 5.2505
R7218 a_19190_29290.n18 a_19190_29290.n10 4.5005
R7219 a_19190_29290.n18 a_19190_29290.n14 0.78175
R7220 a_17540_31010.n1 a_17540_31010.t7 238.322
R7221 a_17540_31010.n1 a_17540_31010.t6 238.322
R7222 a_17540_31010.n3 a_17540_31010.n1 168.8
R7223 a_17540_31010.n0 a_17540_31010.t1 130
R7224 a_17540_31010.n5 a_17540_31010.n4 105.171
R7225 a_17540_31010.n3 a_17540_31010.n2 105.171
R7226 a_17540_31010.n0 a_17540_31010.t0 83.3658
R7227 a_17540_31010.n4 a_17540_31010.n0 35.4806
R7228 a_17540_31010.n2 a_17540_31010.t3 13.1338
R7229 a_17540_31010.n2 a_17540_31010.t2 13.1338
R7230 a_17540_31010.n5 a_17540_31010.t4 13.1338
R7231 a_17540_31010.t5 a_17540_31010.n5 13.1338
R7232 a_17540_31010.n4 a_17540_31010.n3 3.3755
R7233 a_26390_26310.n9 a_26390_26310.t2 729.933
R7234 a_26390_26310.n8 a_26390_26310.t1 729.933
R7235 a_26390_26310.n3 a_26390_26310.n2 718.41
R7236 a_26390_26310.n2 a_26390_26310.n1 660.706
R7237 a_26390_26310.n0 a_26390_26310.t11 361.5
R7238 a_26390_26310.n7 a_26390_26310.n6 342.757
R7239 a_26390_26310.n0 a_26390_26310.t4 281.168
R7240 a_26390_26310.t0 a_26390_26310.n9 260.733
R7241 a_26390_26310.n4 a_26390_26310.n3 224.934
R7242 a_26390_26310.n7 a_26390_26310.t3 190.123
R7243 a_26390_26310.n8 a_26390_26310.n7 180.8
R7244 a_26390_26310.n3 a_26390_26310.t8 168.701
R7245 a_26390_26310.n0 a_26390_26310.t10 152.633
R7246 a_26390_26310.n1 a_26390_26310.t6 152.633
R7247 a_26390_26310.n4 a_26390_26310.t12 136.567
R7248 a_26390_26310.n5 a_26390_26310.t9 136.567
R7249 a_26390_26310.n6 a_26390_26310.t5 136.567
R7250 a_26390_26310.n2 a_26390_26310.t7 131.976
R7251 a_26390_26310.n1 a_26390_26310.n0 128.534
R7252 a_26390_26310.n5 a_26390_26310.n4 128.534
R7253 a_26390_26310.n6 a_26390_26310.n5 128.534
R7254 a_26390_26310.n9 a_26390_26310.n8 57.6005
R7255 a_26420_26230.t0 a_26420_26230.t1 96.0005
R7256 a_26420_26340.n0 a_26420_26340.t1 713.933
R7257 a_26420_26340.n0 a_26420_26340.t2 314.233
R7258 a_26420_26340.t0 a_26420_26340.n0 308.2
R7259 a_18180_28430.n0 a_18180_28430.n2 199.935
R7260 a_18180_28430.n0 a_18180_28430.n3 199.53
R7261 a_18180_28430.n0 a_18180_28430.n4 199.53
R7262 a_18180_28430.n1 a_18180_28430.n5 199.53
R7263 a_18180_28430.n6 a_18180_28430.n1 199.53
R7264 a_18180_28430.n1 a_18180_28430.t5 55.175
R7265 a_18180_28430.n2 a_18180_28430.t10 48.0005
R7266 a_18180_28430.n2 a_18180_28430.t1 48.0005
R7267 a_18180_28430.n3 a_18180_28430.t2 48.0005
R7268 a_18180_28430.n3 a_18180_28430.t6 48.0005
R7269 a_18180_28430.n4 a_18180_28430.t8 48.0005
R7270 a_18180_28430.n4 a_18180_28430.t0 48.0005
R7271 a_18180_28430.n5 a_18180_28430.t4 48.0005
R7272 a_18180_28430.n5 a_18180_28430.t7 48.0005
R7273 a_18180_28430.t9 a_18180_28430.n6 48.0005
R7274 a_18180_28430.n6 a_18180_28430.t3 48.0005
R7275 a_18180_28430.n1 a_18180_28430.n0 1.09425
R7276 a_14990_33500.n3 a_14990_33500.t6 291.503
R7277 a_14990_33500.n3 a_14990_33500.t10 291.288
R7278 a_14990_33500.n4 a_14990_33500.t8 291.288
R7279 a_14990_33500.n5 a_14990_33500.t9 291.288
R7280 a_14990_33500.n6 a_14990_33500.t7 291.288
R7281 a_14990_33500.t0 a_14990_33500.n8 165.601
R7282 a_14990_33500.n8 a_14990_33500.t1 108.424
R7283 a_14990_33500.n2 a_14990_33500.n0 105.609
R7284 a_14990_33500.n2 a_14990_33500.n1 104.484
R7285 a_14990_33500.n8 a_14990_33500.n7 21.4246
R7286 a_14990_33500.n7 a_14990_33500.n2 14.2349
R7287 a_14990_33500.n0 a_14990_33500.t5 13.1338
R7288 a_14990_33500.n0 a_14990_33500.t4 13.1338
R7289 a_14990_33500.n1 a_14990_33500.t3 13.1338
R7290 a_14990_33500.n1 a_14990_33500.t2 13.1338
R7291 a_14990_33500.n7 a_14990_33500.n6 6.43621
R7292 a_14990_33500.n4 a_14990_33500.n3 0.643357
R7293 a_14990_33500.n6 a_14990_33500.n5 0.643357
R7294 a_14990_33500.n5 a_14990_33500.n4 0.214786
R7295 a_26390_27520.n0 a_26390_27520.t0 663.801
R7296 a_26390_27520.t5 a_26390_27520.t3 514.134
R7297 a_26390_27520.n0 a_26390_27520.t5 479.284
R7298 a_26390_27520.n3 a_26390_27520.n2 320.7
R7299 a_26390_27520.t1 a_26390_27520.n3 275.454
R7300 a_26390_27520.n2 a_26390_27520.t2 265.101
R7301 a_26390_27520.n1 a_26390_27520.t6 265.101
R7302 a_26390_27520.n1 a_26390_27520.t4 136.567
R7303 a_26390_27520.n2 a_26390_27520.n1 112.468
R7304 a_26390_27520.n3 a_26390_27520.n0 97.9205
R7305 a_26310_26200.n8 a_26310_26200.n7 949.764
R7306 a_26310_26200.n3 a_26310_26200.n2 895.144
R7307 a_26310_26200.t10 a_26310_26200.t8 819.4
R7308 a_26310_26200.n10 a_26310_26200.n9 628.734
R7309 a_26310_26200.n2 a_26310_26200.n1 496.262
R7310 a_26310_26200.n0 a_26310_26200.t5 361.5
R7311 a_26310_26200.n8 a_26310_26200.t10 336.25
R7312 a_26310_26200.n7 a_26310_26200.n6 321.334
R7313 a_26310_26200.n0 a_26310_26200.t7 281.168
R7314 a_26310_26200.n9 a_26310_26200.t2 257.534
R7315 a_26310_26200.n4 a_26310_26200.n3 208.868
R7316 a_26310_26200.n4 a_26310_26200.t3 168.701
R7317 a_26310_26200.n3 a_26310_26200.t14 168.701
R7318 a_26310_26200.n0 a_26310_26200.t4 152.633
R7319 a_26310_26200.n1 a_26310_26200.t11 152.633
R7320 a_26310_26200.n5 a_26310_26200.t12 136.567
R7321 a_26310_26200.n6 a_26310_26200.t6 136.567
R7322 a_26310_26200.n2 a_26310_26200.t9 131.976
R7323 a_26310_26200.n1 a_26310_26200.n0 128.534
R7324 a_26310_26200.n6 a_26310_26200.n5 128.534
R7325 a_26310_26200.n7 a_26310_26200.t13 126.927
R7326 a_26310_26200.n10 a_26310_26200.t0 78.8005
R7327 a_26310_26200.t1 a_26310_26200.n10 78.8005
R7328 a_26310_26200.n5 a_26310_26200.n4 48.2005
R7329 a_26310_26200.n9 a_26310_26200.n8 11.2005
R7330 a_24280_30570.n4 a_24280_30570.n3 1295.28
R7331 a_24280_30570.n3 a_24280_30570.t4 586.433
R7332 a_24280_30570.n0 a_24280_30570.t3 388.813
R7333 a_24280_30570.n0 a_24280_30570.t5 356.68
R7334 a_24280_30570.n3 a_24280_30570.t6 249.034
R7335 a_24280_30570.n2 a_24280_30570.n0 225.601
R7336 a_24280_30570.t2 a_24280_30570.n4 221.411
R7337 a_24280_30570.n2 a_24280_30570.n1 163.678
R7338 a_24280_30570.n4 a_24280_30570.n2 84.24
R7339 a_24280_30570.n1 a_24280_30570.t0 24.0005
R7340 a_24280_30570.n1 a_24280_30570.t1 24.0005
R7341 a_24310_31390.t0 a_24310_31390.t1 39.4005
R7342 a_23100_30050.t4 a_23100_30050.t5 835.467
R7343 a_23100_30050.n3 a_23100_30050.t4 564.496
R7344 a_23100_30050.n2 a_23100_30050.t6 538.234
R7345 a_23100_30050.n1 a_23100_30050.t8 517.347
R7346 a_23100_30050.n3 a_23100_30050.n2 431.12
R7347 a_23100_30050.n4 a_23100_30050.n1 369.601
R7348 a_23100_30050.n2 a_23100_30050.t7 297.233
R7349 a_23100_30050.n5 a_23100_30050.n0 244.716
R7350 a_23100_30050.n1 a_23100_30050.t3 228.148
R7351 a_23100_30050.t1 a_23100_30050.n5 221.411
R7352 a_23100_30050.n5 a_23100_30050.n4 47.9734
R7353 a_23100_30050.n4 a_23100_30050.n3 39.5568
R7354 a_23100_30050.n0 a_23100_30050.t2 24.0005
R7355 a_23100_30050.n0 a_23100_30050.t0 24.0005
R7356 a_24280_31090.n2 a_24280_31090.n1 1295.28
R7357 a_24280_31090.t6 a_24280_31090.t4 1188.93
R7358 a_24280_31090.t4 a_24280_31090.t3 835.467
R7359 a_24280_31090.n1 a_24280_31090.t5 586.433
R7360 a_24280_31090.n1 a_24280_31090.t6 249.034
R7361 a_24280_31090.n2 a_24280_31090.n0 247.916
R7362 a_24280_31090.t0 a_24280_31090.n2 221.411
R7363 a_24280_31090.n0 a_24280_31090.t2 24.0005
R7364 a_24280_31090.n0 a_24280_31090.t1 24.0005
R7365 a_24310_31010.t0 a_24310_31010.t1 39.4005
R7366 a_26390_28180.n0 a_26390_28180.t3 729.933
R7367 a_26390_28180.n1 a_26390_28180.t4 547.134
R7368 a_26390_28180.n0 a_26390_28180.t1 260.733
R7369 a_26390_28180.n2 a_26390_28180.n1 212.733
R7370 a_26390_28180.n1 a_26390_28180.n0 57.6005
R7371 a_26390_28180.t2 a_26390_28180.n2 48.0005
R7372 a_26390_28180.n2 a_26390_28180.t0 48.0005
R7373 a_19910_24460.n0 a_19910_24460.t8 1132.7
R7374 a_19910_24460.n1 a_19910_24460.n0 915.801
R7375 a_19910_24460.n12 a_19910_24460.n2 706.639
R7376 a_19910_24460.n2 a_19910_24460.n1 385.601
R7377 a_19910_24460.n4 a_19910_24460.t11 377.567
R7378 a_19910_24460.n3 a_19910_24460.t9 297.233
R7379 a_19910_24460.n5 a_19910_24460.n3 237.851
R7380 a_19910_24460.n9 a_19910_24460.n7 236.501
R7381 a_19910_24460.n5 a_19910_24460.n4 232.809
R7382 a_19910_24460.n0 a_19910_24460.t15 216.9
R7383 a_19910_24460.n1 a_19910_24460.t12 216.9
R7384 a_19910_24460.n2 a_19910_24460.t13 216.9
R7385 a_19910_24460.n4 a_19910_24460.t10 216.9
R7386 a_19910_24460.n9 a_19910_24460.n8 178.901
R7387 a_19910_24460.n3 a_19910_24460.t14 136.567
R7388 a_19910_24460.t0 a_19910_24460.n13 126.139
R7389 a_19910_24460.n11 a_19910_24460.n10 117.546
R7390 a_19910_24460.n10 a_19910_24460.n6 113.061
R7391 a_19910_24460.n11 a_19910_24460.n5 51.2088
R7392 a_19910_24460.n10 a_19910_24460.n9 35.2005
R7393 a_19910_24460.n8 a_19910_24460.t4 24.6255
R7394 a_19910_24460.n8 a_19910_24460.t3 24.6255
R7395 a_19910_24460.n7 a_19910_24460.t6 24.6255
R7396 a_19910_24460.n7 a_19910_24460.t5 24.6255
R7397 a_19910_24460.n6 a_19910_24460.t1 15.0005
R7398 a_19910_24460.n6 a_19910_24460.t2 15.0005
R7399 a_19910_24460.n12 a_19910_24460.n11 11.5239
R7400 a_19910_24460.n13 a_19910_24460.t7 3.82928
R7401 a_19910_24460.n13 a_19910_24460.n12 0.09475
R7402 a_25860_21760.n0 a_25860_21760.t1 284.2
R7403 a_25860_21760.n0 a_25860_21760.t2 233
R7404 a_25860_21760.t0 a_25860_21760.n0 184.191
R7405 a_19940_24490.n1 a_19940_24490.t7 335.793
R7406 a_19940_24490.n5 a_19940_24490.n4 325.248
R7407 a_19940_24490.n4 a_19940_24490.n0 313
R7408 a_19940_24490.n3 a_19940_24490.t4 252.248
R7409 a_19940_24490.n1 a_19940_24490.t6 216.9
R7410 a_19940_24490.n2 a_19940_24490.t2 216.9
R7411 a_19940_24490.n2 a_19940_24490.n1 160.667
R7412 a_19940_24490.n4 a_19940_24490.n3 152
R7413 a_19940_24490.n0 a_19940_24490.t0 60.0005
R7414 a_19940_24490.n0 a_19940_24490.t1 60.0005
R7415 a_19940_24490.n5 a_19940_24490.t5 49.2505
R7416 a_19940_24490.t3 a_19940_24490.n5 49.2505
R7417 a_19940_24490.n3 a_19940_24490.n2 35.3472
R7418 a_23100_29610.n0 a_23100_29610.t3 490.034
R7419 a_23100_29610.n1 a_23100_29610.n0 457.233
R7420 a_23100_29610.n0 a_23100_29610.t4 345.433
R7421 a_23100_29610.n2 a_23100_29610.n1 226.887
R7422 a_23100_29610.n1 a_23100_29610.t2 172.458
R7423 a_23100_29610.t0 a_23100_29610.n2 19.7005
R7424 a_23100_29610.n2 a_23100_29610.t1 19.7005
R7425 a_23100_29280.t0 a_23100_29280.n2 500.086
R7426 a_23100_29280.n0 a_23100_29280.t2 490.034
R7427 a_23100_29280.t0 a_23100_29280.n2 461.389
R7428 a_23100_29280.n1 a_23100_29280.n0 449.233
R7429 a_23100_29280.n0 a_23100_29280.t3 345.433
R7430 a_23100_29280.n1 a_23100_29280.t1 177.577
R7431 a_23100_29280.n2 a_23100_29280.n1 48.3899
R7432 a_14558_34050.n0 a_14558_34050.t25 403.952
R7433 a_14558_34050.n18 a_14558_34050.t26 403.755
R7434 a_14558_34050.n17 a_14558_34050.t23 403.755
R7435 a_14558_34050.n16 a_14558_34050.t14 403.755
R7436 a_14558_34050.n15 a_14558_34050.t27 403.755
R7437 a_14558_34050.n14 a_14558_34050.t18 403.755
R7438 a_14558_34050.n13 a_14558_34050.t11 403.755
R7439 a_14558_34050.n12 a_14558_34050.t24 403.755
R7440 a_14558_34050.n11 a_14558_34050.t16 403.755
R7441 a_14558_34050.n10 a_14558_34050.t29 403.755
R7442 a_14558_34050.n9 a_14558_34050.t20 403.755
R7443 a_14558_34050.n8 a_14558_34050.t21 403.755
R7444 a_14558_34050.n7 a_14558_34050.t17 403.755
R7445 a_14558_34050.n6 a_14558_34050.t10 403.755
R7446 a_14558_34050.n5 a_14558_34050.t22 403.755
R7447 a_14558_34050.n4 a_14558_34050.t13 403.755
R7448 a_14558_34050.n3 a_14558_34050.t15 403.755
R7449 a_14558_34050.n2 a_14558_34050.t28 403.755
R7450 a_14558_34050.n1 a_14558_34050.t19 403.755
R7451 a_14558_34050.n0 a_14558_34050.t12 403.755
R7452 a_14558_34050.n26 a_14558_34050.n25 301.933
R7453 a_14558_34050.n24 a_14558_34050.n23 301.933
R7454 a_14558_34050.n22 a_14558_34050.n21 301.933
R7455 a_14558_34050.n20 a_14558_34050.n19 301.933
R7456 a_14558_34050.t9 a_14558_34050.n27 157.238
R7457 a_14558_34050.n20 a_14558_34050.t2 103.826
R7458 a_14558_34050.n25 a_14558_34050.t1 39.4005
R7459 a_14558_34050.n25 a_14558_34050.t4 39.4005
R7460 a_14558_34050.n23 a_14558_34050.t5 39.4005
R7461 a_14558_34050.n23 a_14558_34050.t6 39.4005
R7462 a_14558_34050.n21 a_14558_34050.t7 39.4005
R7463 a_14558_34050.n21 a_14558_34050.t8 39.4005
R7464 a_14558_34050.n19 a_14558_34050.t3 39.4005
R7465 a_14558_34050.n19 a_14558_34050.t0 39.4005
R7466 a_14558_34050.n27 a_14558_34050.n18 10.3335
R7467 a_14558_34050.n27 a_14558_34050.n26 5.313
R7468 a_14558_34050.n9 a_14558_34050.n8 1.6255
R7469 a_14558_34050.n26 a_14558_34050.n24 1.1255
R7470 a_14558_34050.n24 a_14558_34050.n22 1.1255
R7471 a_14558_34050.n22 a_14558_34050.n20 1.1255
R7472 a_14558_34050.n18 a_14558_34050.n17 0.196929
R7473 a_14558_34050.n17 a_14558_34050.n16 0.196929
R7474 a_14558_34050.n16 a_14558_34050.n15 0.196929
R7475 a_14558_34050.n15 a_14558_34050.n14 0.196929
R7476 a_14558_34050.n14 a_14558_34050.n13 0.196929
R7477 a_14558_34050.n13 a_14558_34050.n12 0.196929
R7478 a_14558_34050.n12 a_14558_34050.n11 0.196929
R7479 a_14558_34050.n11 a_14558_34050.n10 0.196929
R7480 a_14558_34050.n10 a_14558_34050.n9 0.196929
R7481 a_14558_34050.n8 a_14558_34050.n7 0.196929
R7482 a_14558_34050.n7 a_14558_34050.n6 0.196929
R7483 a_14558_34050.n6 a_14558_34050.n5 0.196929
R7484 a_14558_34050.n5 a_14558_34050.n4 0.196929
R7485 a_14558_34050.n4 a_14558_34050.n3 0.196929
R7486 a_14558_34050.n3 a_14558_34050.n2 0.196929
R7487 a_14558_34050.n2 a_14558_34050.n1 0.196929
R7488 a_14558_34050.n1 a_14558_34050.n0 0.196929
R7489 a_22190_29430.n5 a_22190_29430.n4 1269.42
R7490 a_22190_29430.n11 a_22190_29430.n10 297.663
R7491 a_22190_29430.n21 a_22190_29430.n20 297.663
R7492 a_22190_29430.n19 a_22190_29430.n18 297.663
R7493 a_22190_29430.n17 a_22190_29430.n15 297.663
R7494 a_22190_29430.n14 a_22190_29430.n13 297.663
R7495 a_22190_29430.n25 a_22190_29430.n24 297.663
R7496 a_22190_29430.n5 a_22190_29430.t2 275.325
R7497 a_22190_29430.n7 a_22190_29430.n6 248.4
R7498 a_22190_29430.n2 a_22190_29430.t5 239.3
R7499 a_22190_29430.n2 a_22190_29430.t4 207.504
R7500 a_22190_29430.n8 a_22190_29430.n2 166.232
R7501 a_22190_29430.n4 a_22190_29430.t19 151.792
R7502 a_22190_29430.n6 a_22190_29430.t0 140.583
R7503 a_22190_29430.n6 a_22190_29430.t2 140.583
R7504 a_22190_29430.n7 a_22190_29430.n3 98.6614
R7505 a_22190_29430.t0 a_22190_29430.n5 80.3338
R7506 a_22190_29430.n4 a_22190_29430.t18 44.2902
R7507 a_22190_29430.n10 a_22190_29430.t6 39.4005
R7508 a_22190_29430.n10 a_22190_29430.t11 39.4005
R7509 a_22190_29430.n20 a_22190_29430.t10 39.4005
R7510 a_22190_29430.n20 a_22190_29430.t15 39.4005
R7511 a_22190_29430.n18 a_22190_29430.t14 39.4005
R7512 a_22190_29430.n18 a_22190_29430.t8 39.4005
R7513 a_22190_29430.n15 a_22190_29430.t12 39.4005
R7514 a_22190_29430.n15 a_22190_29430.t16 39.4005
R7515 a_22190_29430.n13 a_22190_29430.t9 39.4005
R7516 a_22190_29430.n13 a_22190_29430.t7 39.4005
R7517 a_22190_29430.n25 a_22190_29430.t13 39.4005
R7518 a_22190_29430.t17 a_22190_29430.n25 39.4005
R7519 a_22190_29430.n8 a_22190_29430.n7 17.0229
R7520 a_22190_29430.n3 a_22190_29430.t3 15.0005
R7521 a_22190_29430.n3 a_22190_29430.t1 15.0005
R7522 a_22190_29430.n23 a_22190_29430.n11 4.84425
R7523 a_22190_29430.n16 a_22190_29430.n14 4.84425
R7524 a_22190_29430.n17 a_22190_29430.n16 4.5005
R7525 a_22190_29430.n19 a_22190_29430.n12 4.5005
R7526 a_22190_29430.n22 a_22190_29430.n21 4.5005
R7527 a_22190_29430.n24 a_22190_29430.n23 4.5005
R7528 a_22190_29430.n9 a_22190_29430.n8 9.35425
R7529 a_22190_29430.n0 a_22190_29430.n14 1.85607
R7530 a_22190_29430.n11 a_22190_29430.n9 1.74185
R7531 a_22190_29430.n21 a_22190_29430.n1 1.74185
R7532 a_22190_29430.n0 a_22190_29430.n19 1.74185
R7533 a_22190_29430.n0 a_22190_29430.n17 1.74185
R7534 a_22190_29430.n24 a_22190_29430.n1 1.74185
R7535 a_22190_29430.n23 a_22190_29430.n22 0.34425
R7536 a_22190_29430.n22 a_22190_29430.n12 0.34425
R7537 a_22190_29430.n16 a_22190_29430.n12 0.34425
R7538 a_22190_29430.n1 a_22190_29430.n0 0.229667
R7539 a_22190_29430.n9 a_22190_29430.n1 0.229667
R7540 a_26300_23070.n2 a_26300_23070.t0 755.889
R7541 a_26300_23070.n1 a_26300_23070.t4 343.034
R7542 a_26300_23070.t1 a_26300_23070.n2 270.334
R7543 a_26300_23070.n1 a_26300_23070.n0 212.733
R7544 a_26300_23070.n0 a_26300_23070.t3 48.0005
R7545 a_26300_23070.n0 a_26300_23070.t2 48.0005
R7546 a_26300_23070.n2 a_26300_23070.n1 35.2005
R7547 a_26300_22300.t4 a_26300_22300.t3 1012.2
R7548 a_26300_22300.n1 a_26300_22300.t0 663.801
R7549 a_26300_22300.t5 a_26300_22300.t6 401.668
R7550 a_26300_22300.n2 a_26300_22300.n0 400.901
R7551 a_26300_22300.n0 a_26300_22300.t2 377.567
R7552 a_26300_22300.n1 a_26300_22300.t4 361.661
R7553 a_26300_22300.t1 a_26300_22300.n2 314.601
R7554 a_26300_22300.n0 a_26300_22300.t5 281.168
R7555 a_26300_22300.n2 a_26300_22300.n1 73.6005
R7556 a_26420_27440.t0 a_26420_27440.t1 96.0005
R7557 a_26390_29930.n0 a_26390_29930.t3 767.801
R7558 a_26390_29930.n1 a_26390_29930.t4 343.949
R7559 a_26390_29930.n0 a_26390_29930.t1 260.733
R7560 a_26390_29930.n2 a_26390_29930.n1 212.733
R7561 a_26390_29930.n1 a_26390_29930.n0 57.6005
R7562 a_26390_29930.t2 a_26390_29930.n2 48.0005
R7563 a_26390_29930.n2 a_26390_29930.t0 48.0005
R7564 a_14140_28370.n2 a_14140_28370.n0 302.507
R7565 a_14140_28370.n10 a_14140_28370.n9 302.163
R7566 a_14140_28370.n8 a_14140_28370.n7 302.163
R7567 a_14140_28370.n6 a_14140_28370.n5 302.163
R7568 a_14140_28370.n4 a_14140_28370.n3 302.163
R7569 a_14140_28370.n2 a_14140_28370.n1 302.163
R7570 a_14140_28370.n11 a_14140_28370.t13 291.503
R7571 a_14140_28370.n14 a_14140_28370.t17 291.288
R7572 a_14140_28370.n13 a_14140_28370.t15 291.288
R7573 a_14140_28370.n12 a_14140_28370.t16 291.288
R7574 a_14140_28370.n11 a_14140_28370.t14 291.288
R7575 a_14140_28370.t0 a_14140_28370.n15 173.233
R7576 a_14140_28370.n9 a_14140_28370.t1 39.4005
R7577 a_14140_28370.n9 a_14140_28370.t5 39.4005
R7578 a_14140_28370.n7 a_14140_28370.t7 39.4005
R7579 a_14140_28370.n7 a_14140_28370.t11 39.4005
R7580 a_14140_28370.n5 a_14140_28370.t4 39.4005
R7581 a_14140_28370.n5 a_14140_28370.t9 39.4005
R7582 a_14140_28370.n3 a_14140_28370.t12 39.4005
R7583 a_14140_28370.n3 a_14140_28370.t6 39.4005
R7584 a_14140_28370.n1 a_14140_28370.t10 39.4005
R7585 a_14140_28370.n1 a_14140_28370.t3 39.4005
R7586 a_14140_28370.n0 a_14140_28370.t8 39.4005
R7587 a_14140_28370.n0 a_14140_28370.t2 39.4005
R7588 a_14140_28370.n15 a_14140_28370.n10 12.0474
R7589 a_14140_28370.n15 a_14140_28370.n14 6.4005
R7590 a_14140_28370.n14 a_14140_28370.n13 0.643357
R7591 a_14140_28370.n12 a_14140_28370.n11 0.643357
R7592 a_14140_28370.n10 a_14140_28370.n8 0.34425
R7593 a_14140_28370.n8 a_14140_28370.n6 0.34425
R7594 a_14140_28370.n6 a_14140_28370.n4 0.34425
R7595 a_14140_28370.n4 a_14140_28370.n2 0.34425
R7596 a_14140_28370.n13 a_14140_28370.n12 0.214786
R7597 a_26390_31270.n0 a_26390_31270.t3 729.933
R7598 a_26390_31270.n1 a_26390_31270.t4 547.134
R7599 a_26390_31270.n0 a_26390_31270.t0 260.733
R7600 a_26390_31270.n2 a_26390_31270.n1 212.733
R7601 a_26390_31270.n1 a_26390_31270.n0 57.6005
R7602 a_26390_31270.n2 a_26390_31270.t1 48.0005
R7603 a_26390_31270.t2 a_26390_31270.n2 48.0005
R7604 a_13370_29270.t0 a_13370_29270.n130 132.74
R7605 a_13370_29270.n120 a_13370_29270.n5 83.5719
R7606 a_13370_29270.n115 a_13370_29270.n6 83.5719
R7607 a_13370_29270.n127 a_13370_29270.n126 83.5719
R7608 a_13370_29270.n40 a_13370_29270.n2 83.5719
R7609 a_13370_29270.n43 a_13370_29270.n41 83.5719
R7610 a_13370_29270.n50 a_13370_29270.n49 83.5719
R7611 a_13370_29270.n60 a_13370_29270.n59 83.5719
R7612 a_13370_29270.n58 a_13370_29270.n57 83.5719
R7613 a_13370_29270.n56 a_13370_29270.n55 83.5719
R7614 a_13370_29270.n93 a_13370_29270.n14 83.5719
R7615 a_13370_29270.n92 a_13370_29270.n91 83.5719
R7616 a_13370_29270.n83 a_13370_29270.n17 83.5719
R7617 a_13370_29270.n76 a_13370_29270.n18 83.5719
R7618 a_13370_29270.n78 a_13370_29270.n77 83.5719
R7619 a_13370_29270.n70 a_13370_29270.n22 83.5719
R7620 a_13370_29270.n108 a_13370_29270.n107 83.5719
R7621 a_13370_29270.n106 a_13370_29270.n105 83.5719
R7622 a_13370_29270.n104 a_13370_29270.n103 83.5719
R7623 a_13370_29270.n122 a_13370_29270.n5 73.3165
R7624 a_13370_29270.n45 a_13370_29270.n41 73.3165
R7625 a_13370_29270.n56 a_13370_29270.n29 73.3165
R7626 a_13370_29270.n92 a_13370_29270.n15 73.3165
R7627 a_13370_29270.n77 a_13370_29270.n75 73.3165
R7628 a_13370_29270.n104 a_13370_29270.n12 73.3165
R7629 a_13370_29270.n126 a_13370_29270.n125 73.19
R7630 a_13370_29270.n49 a_13370_29270.n48 73.19
R7631 a_13370_29270.n61 a_13370_29270.n60 73.19
R7632 a_13370_29270.n85 a_13370_29270.n17 73.19
R7633 a_13370_29270.n72 a_13370_29270.n22 73.19
R7634 a_13370_29270.n109 a_13370_29270.n108 73.19
R7635 a_13370_29270.n116 a_13370_29270.t7 65.0331
R7636 a_13370_29270.n94 a_13370_29270.t2 65.0331
R7637 a_13370_29270.t4 a_13370_29270.n36 36.6632
R7638 a_13370_29270.n23 a_13370_29270.t8 36.6632
R7639 a_13370_29270.n115 a_13370_29270.n5 26.074
R7640 a_13370_29270.n41 a_13370_29270.n40 26.074
R7641 a_13370_29270.n58 a_13370_29270.n56 26.074
R7642 a_13370_29270.n93 a_13370_29270.n92 26.074
R7643 a_13370_29270.n77 a_13370_29270.n76 26.074
R7644 a_13370_29270.n106 a_13370_29270.n104 26.074
R7645 a_13370_29270.n126 a_13370_29270.t1 25.7843
R7646 a_13370_29270.n49 a_13370_29270.t4 25.7843
R7647 a_13370_29270.n60 a_13370_29270.t3 25.7843
R7648 a_13370_29270.t5 a_13370_29270.n17 25.7843
R7649 a_13370_29270.t8 a_13370_29270.n22 25.7843
R7650 a_13370_29270.n108 a_13370_29270.t6 25.7843
R7651 a_13370_29270.n98 a_13370_29270.n10 9.3005
R7652 a_13370_29270.n98 a_13370_29270.n8 9.3005
R7653 a_13370_29270.n98 a_13370_29270.n11 9.3005
R7654 a_13370_29270.n113 a_13370_29270.n98 9.3005
R7655 a_13370_29270.n100 a_13370_29270.n10 9.3005
R7656 a_13370_29270.n100 a_13370_29270.n8 9.3005
R7657 a_13370_29270.n100 a_13370_29270.n11 9.3005
R7658 a_13370_29270.n113 a_13370_29270.n100 9.3005
R7659 a_13370_29270.n97 a_13370_29270.n10 9.3005
R7660 a_13370_29270.n97 a_13370_29270.n8 9.3005
R7661 a_13370_29270.n97 a_13370_29270.n11 9.3005
R7662 a_13370_29270.n113 a_13370_29270.n97 9.3005
R7663 a_13370_29270.n112 a_13370_29270.n10 9.3005
R7664 a_13370_29270.n112 a_13370_29270.n8 9.3005
R7665 a_13370_29270.n112 a_13370_29270.n11 9.3005
R7666 a_13370_29270.n113 a_13370_29270.n112 9.3005
R7667 a_13370_29270.n96 a_13370_29270.n10 9.3005
R7668 a_13370_29270.n96 a_13370_29270.n8 9.3005
R7669 a_13370_29270.n96 a_13370_29270.n11 9.3005
R7670 a_13370_29270.n96 a_13370_29270.n7 9.3005
R7671 a_13370_29270.n113 a_13370_29270.n96 9.3005
R7672 a_13370_29270.n114 a_13370_29270.n10 9.3005
R7673 a_13370_29270.n114 a_13370_29270.n8 9.3005
R7674 a_13370_29270.n114 a_13370_29270.n11 9.3005
R7675 a_13370_29270.n114 a_13370_29270.n7 9.3005
R7676 a_13370_29270.n114 a_13370_29270.n113 9.3005
R7677 a_13370_29270.n31 a_13370_29270.n27 9.3005
R7678 a_13370_29270.n31 a_13370_29270.n26 9.3005
R7679 a_13370_29270.n31 a_13370_29270.n28 9.3005
R7680 a_13370_29270.n65 a_13370_29270.n31 9.3005
R7681 a_13370_29270.n33 a_13370_29270.n27 9.3005
R7682 a_13370_29270.n33 a_13370_29270.n26 9.3005
R7683 a_13370_29270.n33 a_13370_29270.n28 9.3005
R7684 a_13370_29270.n65 a_13370_29270.n33 9.3005
R7685 a_13370_29270.n30 a_13370_29270.n27 9.3005
R7686 a_13370_29270.n30 a_13370_29270.n26 9.3005
R7687 a_13370_29270.n30 a_13370_29270.n28 9.3005
R7688 a_13370_29270.n65 a_13370_29270.n30 9.3005
R7689 a_13370_29270.n35 a_13370_29270.n27 9.3005
R7690 a_13370_29270.n35 a_13370_29270.n26 9.3005
R7691 a_13370_29270.n35 a_13370_29270.n28 9.3005
R7692 a_13370_29270.n65 a_13370_29270.n35 9.3005
R7693 a_13370_29270.n66 a_13370_29270.n27 9.3005
R7694 a_13370_29270.n66 a_13370_29270.n26 9.3005
R7695 a_13370_29270.n66 a_13370_29270.n28 9.3005
R7696 a_13370_29270.n66 a_13370_29270.n25 9.3005
R7697 a_13370_29270.n66 a_13370_29270.n65 9.3005
R7698 a_13370_29270.n64 a_13370_29270.n27 9.3005
R7699 a_13370_29270.n64 a_13370_29270.n26 9.3005
R7700 a_13370_29270.n64 a_13370_29270.n28 9.3005
R7701 a_13370_29270.n64 a_13370_29270.n25 9.3005
R7702 a_13370_29270.n65 a_13370_29270.n64 9.3005
R7703 a_13370_29270.n99 a_13370_29270.n7 4.64654
R7704 a_13370_29270.n110 a_13370_29270.n102 4.64654
R7705 a_13370_29270.n101 a_13370_29270.n7 4.64654
R7706 a_13370_29270.n111 a_13370_29270.n110 4.64654
R7707 a_13370_29270.n110 a_13370_29270.n9 4.64654
R7708 a_13370_29270.n32 a_13370_29270.n25 4.64654
R7709 a_13370_29270.n62 a_13370_29270.n54 4.64654
R7710 a_13370_29270.n34 a_13370_29270.n25 4.64654
R7711 a_13370_29270.n62 a_13370_29270.n24 4.64654
R7712 a_13370_29270.n63 a_13370_29270.n62 4.64654
R7713 a_13370_29270.n125 a_13370_29270.n124 2.36206
R7714 a_13370_29270.n48 a_13370_29270.n47 2.36206
R7715 a_13370_29270.n86 a_13370_29270.n85 2.36206
R7716 a_13370_29270.n73 a_13370_29270.n72 2.36206
R7717 a_13370_29270.n123 a_13370_29270.n122 2.19742
R7718 a_13370_29270.n46 a_13370_29270.n45 2.19742
R7719 a_13370_29270.n87 a_13370_29270.n15 2.19742
R7720 a_13370_29270.n75 a_13370_29270.n74 2.19742
R7721 a_13370_29270.n51 a_13370_29270.n36 1.80777
R7722 a_13370_29270.n69 a_13370_29270.n23 1.80777
R7723 a_13370_29270.n116 a_13370_29270.n6 1.56484
R7724 a_13370_29270.n94 a_13370_29270.n14 1.56484
R7725 a_13370_29270.n71 a_13370_29270.n21 1.5505
R7726 a_13370_29270.n69 a_13370_29270.n68 1.5505
R7727 a_13370_29270.n84 a_13370_29270.n16 1.5505
R7728 a_13370_29270.n82 a_13370_29270.n81 1.5505
R7729 a_13370_29270.n80 a_13370_29270.n79 1.5505
R7730 a_13370_29270.n20 a_13370_29270.n19 1.5505
R7731 a_13370_29270.n90 a_13370_29270.n13 1.5505
R7732 a_13370_29270.n89 a_13370_29270.n88 1.5505
R7733 a_13370_29270.n38 a_13370_29270.n37 1.5505
R7734 a_13370_29270.n52 a_13370_29270.n51 1.5505
R7735 a_13370_29270.n3 a_13370_29270.n1 1.5505
R7736 a_13370_29270.n129 a_13370_29270.n128 1.5505
R7737 a_13370_29270.n42 a_13370_29270.n0 1.5505
R7738 a_13370_29270.n44 a_13370_29270.n39 1.5505
R7739 a_13370_29270.n119 a_13370_29270.n118 1.5505
R7740 a_13370_29270.n121 a_13370_29270.n4 1.5505
R7741 a_13370_29270.n127 a_13370_29270.n3 1.25468
R7742 a_13370_29270.n50 a_13370_29270.n38 1.25468
R7743 a_13370_29270.n59 a_13370_29270.n27 1.25468
R7744 a_13370_29270.n84 a_13370_29270.n83 1.25468
R7745 a_13370_29270.n71 a_13370_29270.n70 1.25468
R7746 a_13370_29270.n107 a_13370_29270.n10 1.25468
R7747 a_13370_29270.n122 a_13370_29270.n121 1.19225
R7748 a_13370_29270.n45 a_13370_29270.n44 1.19225
R7749 a_13370_29270.n29 a_13370_29270.n25 1.19225
R7750 a_13370_29270.n89 a_13370_29270.n15 1.19225
R7751 a_13370_29270.n75 a_13370_29270.n20 1.19225
R7752 a_13370_29270.n12 a_13370_29270.n7 1.19225
R7753 a_13370_29270.n128 a_13370_29270.n2 1.07024
R7754 a_13370_29270.n57 a_13370_29270.n26 1.07024
R7755 a_13370_29270.n82 a_13370_29270.n18 1.07024
R7756 a_13370_29270.n105 a_13370_29270.n8 1.07024
R7757 a_13370_29270.n67 a_13370_29270.n23 1.04793
R7758 a_13370_29270.n53 a_13370_29270.n36 1.04793
R7759 a_13370_29270.n125 a_13370_29270.n3 1.0237
R7760 a_13370_29270.n48 a_13370_29270.n38 1.0237
R7761 a_13370_29270.n61 a_13370_29270.n27 1.0237
R7762 a_13370_29270.n85 a_13370_29270.n84 1.0237
R7763 a_13370_29270.n72 a_13370_29270.n71 1.0237
R7764 a_13370_29270.n109 a_13370_29270.n10 1.0237
R7765 a_13370_29270.n121 a_13370_29270.n120 0.959578
R7766 a_13370_29270.n44 a_13370_29270.n43 0.959578
R7767 a_13370_29270.n55 a_13370_29270.n25 0.959578
R7768 a_13370_29270.n91 a_13370_29270.n89 0.959578
R7769 a_13370_29270.n78 a_13370_29270.n20 0.959578
R7770 a_13370_29270.n103 a_13370_29270.n7 0.959578
R7771 a_13370_29270.n120 a_13370_29270.n119 0.885803
R7772 a_13370_29270.n43 a_13370_29270.n42 0.885803
R7773 a_13370_29270.n55 a_13370_29270.n28 0.885803
R7774 a_13370_29270.n91 a_13370_29270.n90 0.885803
R7775 a_13370_29270.n79 a_13370_29270.n78 0.885803
R7776 a_13370_29270.n103 a_13370_29270.n11 0.885803
R7777 a_13370_29270.n62 a_13370_29270.n61 0.812055
R7778 a_13370_29270.n110 a_13370_29270.n109 0.812055
R7779 a_13370_29270.n119 a_13370_29270.n6 0.77514
R7780 a_13370_29270.n42 a_13370_29270.n2 0.77514
R7781 a_13370_29270.n57 a_13370_29270.n28 0.77514
R7782 a_13370_29270.n90 a_13370_29270.n14 0.77514
R7783 a_13370_29270.n79 a_13370_29270.n18 0.77514
R7784 a_13370_29270.n105 a_13370_29270.n11 0.77514
R7785 a_13370_29270.n65 a_13370_29270.n29 0.647417
R7786 a_13370_29270.n113 a_13370_29270.n12 0.647417
R7787 a_13370_29270.n128 a_13370_29270.n127 0.590702
R7788 a_13370_29270.n51 a_13370_29270.n50 0.590702
R7789 a_13370_29270.n59 a_13370_29270.n26 0.590702
R7790 a_13370_29270.n83 a_13370_29270.n82 0.590702
R7791 a_13370_29270.n70 a_13370_29270.n69 0.590702
R7792 a_13370_29270.n107 a_13370_29270.n8 0.590702
R7793 a_13370_29270.n95 a_13370_29270.n94 0.531214
R7794 a_13370_29270.n117 a_13370_29270.n116 0.531214
R7795 a_13370_29270.t7 a_13370_29270.n115 0.290206
R7796 a_13370_29270.n40 a_13370_29270.t1 0.290206
R7797 a_13370_29270.t3 a_13370_29270.n58 0.290206
R7798 a_13370_29270.t2 a_13370_29270.n93 0.290206
R7799 a_13370_29270.n76 a_13370_29270.t5 0.290206
R7800 a_13370_29270.t6 a_13370_29270.n106 0.290206
R7801 a_13370_29270.n74 a_13370_29270.n73 0.154071
R7802 a_13370_29270.n87 a_13370_29270.n86 0.154071
R7803 a_13370_29270.n47 a_13370_29270.n46 0.154071
R7804 a_13370_29270.n124 a_13370_29270.n123 0.154071
R7805 a_13370_29270.n117 a_13370_29270.n114 0.137464
R7806 a_13370_29270.n64 a_13370_29270.n53 0.137464
R7807 a_13370_29270.n96 a_13370_29270.n95 0.134964
R7808 a_13370_29270.n67 a_13370_29270.n66 0.134964
R7809 a_13370_29270.n68 a_13370_29270.n21 0.0183571
R7810 a_13370_29270.n73 a_13370_29270.n21 0.0183571
R7811 a_13370_29270.n74 a_13370_29270.n19 0.0183571
R7812 a_13370_29270.n80 a_13370_29270.n19 0.0183571
R7813 a_13370_29270.n81 a_13370_29270.n80 0.0183571
R7814 a_13370_29270.n81 a_13370_29270.n16 0.0183571
R7815 a_13370_29270.n86 a_13370_29270.n16 0.0183571
R7816 a_13370_29270.n88 a_13370_29270.n87 0.0183571
R7817 a_13370_29270.n88 a_13370_29270.n13 0.0183571
R7818 a_13370_29270.n52 a_13370_29270.n37 0.0183571
R7819 a_13370_29270.n47 a_13370_29270.n37 0.0183571
R7820 a_13370_29270.n46 a_13370_29270.n39 0.0183571
R7821 a_13370_29270.n39 a_13370_29270.n0 0.0183571
R7822 a_13370_29270.n129 a_13370_29270.n1 0.0183571
R7823 a_13370_29270.n124 a_13370_29270.n1 0.0183571
R7824 a_13370_29270.n123 a_13370_29270.n4 0.0183571
R7825 a_13370_29270.n118 a_13370_29270.n4 0.0183571
R7826 a_13370_29270.n68 a_13370_29270.n67 0.0106786
R7827 a_13370_29270.n53 a_13370_29270.n52 0.0106786
R7828 a_13370_29270.n130 a_13370_29270.n129 0.0106786
R7829 a_13370_29270.n114 a_13370_29270.n9 0.00992001
R7830 a_13370_29270.n100 a_13370_29270.n99 0.00992001
R7831 a_13370_29270.n102 a_13370_29270.n97 0.00992001
R7832 a_13370_29270.n112 a_13370_29270.n101 0.00992001
R7833 a_13370_29270.n111 a_13370_29270.n96 0.00992001
R7834 a_13370_29270.n98 a_13370_29270.n9 0.00992001
R7835 a_13370_29270.n99 a_13370_29270.n98 0.00992001
R7836 a_13370_29270.n102 a_13370_29270.n100 0.00992001
R7837 a_13370_29270.n101 a_13370_29270.n97 0.00992001
R7838 a_13370_29270.n112 a_13370_29270.n111 0.00992001
R7839 a_13370_29270.n64 a_13370_29270.n63 0.00992001
R7840 a_13370_29270.n33 a_13370_29270.n32 0.00992001
R7841 a_13370_29270.n54 a_13370_29270.n30 0.00992001
R7842 a_13370_29270.n35 a_13370_29270.n34 0.00992001
R7843 a_13370_29270.n66 a_13370_29270.n24 0.00992001
R7844 a_13370_29270.n63 a_13370_29270.n31 0.00992001
R7845 a_13370_29270.n32 a_13370_29270.n31 0.00992001
R7846 a_13370_29270.n54 a_13370_29270.n33 0.00992001
R7847 a_13370_29270.n34 a_13370_29270.n30 0.00992001
R7848 a_13370_29270.n35 a_13370_29270.n24 0.00992001
R7849 a_13370_29270.n95 a_13370_29270.n13 0.00817857
R7850 a_13370_29270.n130 a_13370_29270.n0 0.00817857
R7851 a_13370_29270.n118 a_13370_29270.n117 0.00817857
R7852 a_24280_31990.n3 a_24280_31990.t7 796.295
R7853 a_24280_31990.n1 a_24280_31990.t1 761.4
R7854 a_24280_31990.n4 a_24280_31990.n3 631.564
R7855 a_24280_31990.n0 a_24280_31990.t2 538.234
R7856 a_24280_31990.t7 a_24280_31990.t5 514.134
R7857 a_24280_31990.n1 a_24280_31990.n0 435.952
R7858 a_24280_31990.n2 a_24280_31990.t4 313.3
R7859 a_24280_31990.n0 a_24280_31990.t3 297.233
R7860 a_24280_31990.t0 a_24280_31990.n4 233
R7861 a_24280_31990.n2 a_24280_31990.t6 200.833
R7862 a_24280_31990.n3 a_24280_31990.n2 160.667
R7863 a_24280_31990.n4 a_24280_31990.n1 46.7205
R7864 a_26640_21160.t0 a_26640_21160.n0 421.027
R7865 a_26640_21160.n0 a_26640_21160.t2 348.81
R7866 a_26640_21160.n0 a_26640_21160.t1 316.159
R7867 a_24280_27770.n0 a_24280_27770.t3 1004.17
R7868 a_24280_27770.n2 a_24280_27770.n1 545.634
R7869 a_24280_27770.t1 a_24280_27770.n3 458.818
R7870 a_24280_27770.t1 a_24280_27770.n3 429.281
R7871 a_24280_27770.n1 a_24280_27770.t5 425.767
R7872 a_24280_27770.n1 a_24280_27770.n0 417.733
R7873 a_24280_27770.n0 a_24280_27770.t2 409.7
R7874 a_24280_27770.n1 a_24280_27770.t4 409.7
R7875 a_24280_27770.n2 a_24280_27770.t0 173.095
R7876 a_24280_27770.n3 a_24280_27770.n2 36.568
R7877 a_24310_27670.t1 a_24310_27670.n4 458.818
R7878 a_24310_27670.t1 a_24310_27670.n4 429.281
R7879 a_24310_27670.t5 a_24310_27670.t3 377.567
R7880 a_24310_27670.n0 a_24310_27670.t4 326.658
R7881 a_24310_27670.n2 a_24310_27670.n1 252.345
R7882 a_24310_27670.n1 a_24310_27670.n0 196.817
R7883 a_24310_27670.n3 a_24310_27670.t0 164.775
R7884 a_24310_27670.n2 a_24310_27670.t2 164.775
R7885 a_24310_27670.n3 a_24310_27670.n2 112.001
R7886 a_24310_27670.n1 a_24310_27670.t5 92.3838
R7887 a_24310_27670.t3 a_24310_27670.n0 92.3838
R7888 a_24310_27670.n4 a_24310_27670.n3 60.248
R7889 a_23130_29200.t0 a_23130_29200.n2 500.086
R7890 a_23130_29200.n0 a_23130_29200.t2 490.034
R7891 a_23130_29200.t0 a_23130_29200.n2 461.389
R7892 a_23130_29200.n1 a_23130_29200.n0 368.524
R7893 a_23130_29200.n0 a_23130_29200.t3 345.433
R7894 a_23130_29200.n1 a_23130_29200.t1 177.577
R7895 a_23130_29200.n2 a_23130_29200.n1 48.3899
R7896 a_24280_29730.t0 a_24280_29730.n2 500.086
R7897 a_24280_29730.n0 a_24280_29730.t2 490.034
R7898 a_24280_29730.t0 a_24280_29730.n2 461.389
R7899 a_24280_29730.n1 a_24280_29730.n0 449.233
R7900 a_24280_29730.n0 a_24280_29730.t3 345.433
R7901 a_24280_29730.n1 a_24280_29730.t1 177.577
R7902 a_24280_29730.n2 a_24280_29730.n1 48.3899
R7903 a_26300_24370.n0 a_26300_24370.t1 755.889
R7904 a_26300_24370.n1 a_26300_24370.t4 343.034
R7905 a_26300_24370.n0 a_26300_24370.t3 270.334
R7906 a_26300_24370.n2 a_26300_24370.n1 212.733
R7907 a_26300_24370.t0 a_26300_24370.n2 48.0005
R7908 a_26300_24370.n2 a_26300_24370.t2 48.0005
R7909 a_26300_24370.n1 a_26300_24370.n0 35.2005
R7910 a_26300_23600.t4 a_26300_23600.t3 1012.2
R7911 a_26300_23600.n1 a_26300_23600.t0 663.801
R7912 a_26300_23600.t5 a_26300_23600.t6 401.668
R7913 a_26300_23600.n2 a_26300_23600.n0 400.901
R7914 a_26300_23600.n0 a_26300_23600.t2 377.567
R7915 a_26300_23600.n1 a_26300_23600.t4 361.661
R7916 a_26300_23600.t1 a_26300_23600.n2 314.601
R7917 a_26300_23600.n0 a_26300_23600.t5 281.168
R7918 a_26300_23600.n2 a_26300_23600.n1 73.6005
R7919 a_26390_30500.n0 a_26390_30500.t0 719.801
R7920 a_26390_30500.t3 a_26390_30500.t2 514.134
R7921 a_26390_30500.n0 a_26390_30500.t3 332.783
R7922 a_26390_30500.t1 a_26390_30500.n0 330.601
R7923 a_26420_30420.n0 a_26420_30420.t2 531.067
R7924 a_26420_30420.n0 a_26420_30420.t1 48.0005
R7925 a_26420_30420.t0 a_26420_30420.n0 48.0005
R7926 ua[1].n3 ua[1].n1 409.7
R7927 ua[1].t4 ua[1].t6 401.668
R7928 ua[1].n1 ua[1].t3 377.567
R7929 ua[1].n0 ua[1].t0 372.118
R7930 ua[1].n1 ua[1].t4 281.168
R7931 ua[1].n2 ua[1].t5 249.034
R7932 ua[1].n0 ua[1].t1 247.934
R7933 ua[1].n3 ua[1].n2 200.833
R7934 ua[1].n4 ua[1].n3 171.457
R7935 ua[1].n2 ua[1].t2 168.701
R7936 ua[1].n4 ua[1].n0 65.3005
R7937 ua[1] ua[1].n4 18.0284
R7938 a_26400_21130.n1 a_26400_21130.n0 413.634
R7939 a_26400_21130.t1 a_26400_21130.n1 372.118
R7940 a_26400_21130.n0 a_26400_21130.t2 249.034
R7941 a_26400_21130.n1 a_26400_21130.t0 247.934
R7942 a_26400_21130.n0 a_26400_21130.t3 168.701
R7943 a_26420_27220.n0 a_26420_27220.t1 691.534
R7944 a_26420_27220.n1 a_26420_27220.t2 663.801
R7945 a_26420_27220.n0 a_26420_27220.t3 527.867
R7946 a_26420_27220.t0 a_26420_27220.n1 372.2
R7947 a_26420_27220.n1 a_26420_27220.n0 85.3338
R7948 a_26390_32300.n0 a_26390_32300.t0 767.801
R7949 a_26390_32300.n1 a_26390_32300.t4 343.034
R7950 a_26390_32300.n0 a_26390_32300.t1 260.733
R7951 a_26390_32300.n2 a_26390_32300.n1 212.733
R7952 a_26390_32300.n1 a_26390_32300.n0 57.6005
R7953 a_26390_32300.n2 a_26390_32300.t2 48.0005
R7954 a_26390_32300.t3 a_26390_32300.n2 48.0005
R7955 ua[0] ua[0].n0 546.412
R7956 ua[0].n0 ua[0].t0 538.234
R7957 ua[0].n0 ua[0].t1 297.233
R7958 a_23550_31910.t0 a_23550_31910.t1 39.4005
R7959 a_26300_24900.t4 a_26300_24900.t2 1012.2
R7960 a_26300_24900.n1 a_26300_24900.t0 663.801
R7961 a_26300_24900.t5 a_26300_24900.t6 401.668
R7962 a_26300_24900.n2 a_26300_24900.n0 400.901
R7963 a_26300_24900.n1 a_26300_24900.t4 361.661
R7964 a_26300_24900.t1 a_26300_24900.n2 314.601
R7965 a_26300_24900.n0 a_26300_24900.t5 281.168
R7966 a_26300_24900.n0 a_26300_24900.t3 232.968
R7967 a_26300_24900.n2 a_26300_24900.n1 73.6005
R7968 a_24310_30490.t0 a_24310_30490.t1 39.4005
R7969 a_24280_30980.n1 a_24280_30980.t3 517.347
R7970 a_24280_30980.n2 a_24280_30980.n1 417.574
R7971 a_24280_30980.n2 a_24280_30980.n0 244.716
R7972 a_24280_30980.n1 a_24280_30980.t4 228.148
R7973 a_24280_30980.t0 a_24280_30980.n2 221.411
R7974 a_24280_30980.n0 a_24280_30980.t1 24.0005
R7975 a_24280_30980.n0 a_24280_30980.t2 24.0005
R7976 a_26400_20530.n1 a_26400_20530.n0 413.634
R7977 a_26400_20530.t0 a_26400_20530.n1 372.118
R7978 a_26400_20530.n0 a_26400_20530.t2 249.034
R7979 a_26400_20530.n1 a_26400_20530.t1 247.934
R7980 a_26400_20530.n0 a_26400_20530.t3 168.701
R7981 a_26640_20560.t0 a_26640_20560.n0 421.027
R7982 a_26640_20560.n0 a_26640_20560.t2 348.81
R7983 a_26640_20560.n0 a_26640_20560.t1 316.159
R7984 a_26740_30530.t0 a_26740_30530.t1 157.601
R7985 a_23020_31090.n2 a_23020_31090.n0 1295.28
R7986 a_23020_31090.t4 a_23020_31090.t6 1188.93
R7987 a_23020_31090.t6 a_23020_31090.t5 835.467
R7988 a_23020_31090.n0 a_23020_31090.t3 586.433
R7989 a_23020_31090.n0 a_23020_31090.t4 249.034
R7990 a_23020_31090.n2 a_23020_31090.n1 247.917
R7991 a_23020_31090.t2 a_23020_31090.n2 221.411
R7992 a_23020_31090.n1 a_23020_31090.t0 24.0005
R7993 a_23020_31090.n1 a_23020_31090.t1 24.0005
R7994 a_26300_22410.n4 a_26300_22410.t0 758.734
R7995 a_26300_22410.t1 a_26300_22410.n5 758.734
R7996 a_26300_22410.n0 a_26300_22410.t4 538.234
R7997 a_26300_22410.n3 a_26300_22410.n2 342.757
R7998 a_26300_22410.n5 a_26300_22410.t2 260.733
R7999 a_26300_22410.n3 a_26300_22410.t6 190.123
R8000 a_26300_22410.n4 a_26300_22410.n3 180.8
R8001 a_26300_22410.n0 a_26300_22410.t5 136.567
R8002 a_26300_22410.n1 a_26300_22410.t3 136.567
R8003 a_26300_22410.n2 a_26300_22410.t7 136.567
R8004 a_26300_22410.n1 a_26300_22410.n0 128.534
R8005 a_26300_22410.n2 a_26300_22410.n1 128.534
R8006 a_26300_22410.n5 a_26300_22410.n4 57.6005
R8007 a_26390_26970.n2 a_26390_26970.t0 727.09
R8008 a_26390_26970.n1 a_26390_26970.t4 343.949
R8009 a_26390_26970.t3 a_26390_26970.n2 270.334
R8010 a_26390_26970.n1 a_26390_26970.n0 212.733
R8011 a_26390_26970.n0 a_26390_26970.t1 48.0005
R8012 a_26390_26970.n0 a_26390_26970.t2 48.0005
R8013 a_26390_26970.n2 a_26390_26970.n1 35.2005
R8014 a_25350_8708.t0 a_25350_8708.t1 127.201
R8015 a_13742_34050.t20 a_13742_34050.t11 178.589
R8016 a_13742_34050.t12 a_13742_34050.t5 0.1603
R8017 a_13742_34050.t6 a_13742_34050.t12 0.1603
R8018 a_13742_34050.t14 a_13742_34050.t6 0.1603
R8019 a_13742_34050.t18 a_13742_34050.t14 0.1603
R8020 a_13742_34050.t1 a_13742_34050.t18 0.1603
R8021 a_13742_34050.t19 a_13742_34050.t1 0.1603
R8022 a_13742_34050.t3 a_13742_34050.t19 0.1603
R8023 a_13742_34050.t9 a_13742_34050.t3 0.1603
R8024 a_13742_34050.t8 a_13742_34050.t15 0.1603
R8025 a_13742_34050.t2 a_13742_34050.t8 0.1603
R8026 a_13742_34050.t7 a_13742_34050.t2 0.1603
R8027 a_13742_34050.t0 a_13742_34050.t7 0.1603
R8028 a_13742_34050.t17 a_13742_34050.t0 0.1603
R8029 a_13742_34050.t13 a_13742_34050.t17 0.1603
R8030 a_13742_34050.t16 a_13742_34050.t13 0.1603
R8031 a_13742_34050.t11 a_13742_34050.t16 0.1603
R8032 a_13742_34050.t10 a_13742_34050.n0 0.159278
R8033 a_13742_34050.t15 a_13742_34050.t10 0.137822
R8034 a_13742_34050.n0 a_13742_34050.t9 0.1368
R8035 a_13742_34050.n0 a_13742_34050.t4 0.00152174
R8036 a_23020_29890.t4 a_23020_29890.t3 835.467
R8037 a_23020_29890.n0 a_23020_29890.t7 517.347
R8038 a_23020_29890.n1 a_23020_29890.t5 490.034
R8039 a_23020_29890.n2 a_23020_29890.n1 429.932
R8040 a_23020_29890.n2 a_23020_29890.t4 394.267
R8041 a_23020_29890.n1 a_23020_29890.t6 345.433
R8042 a_23020_29890.n5 a_23020_29890.n4 244.715
R8043 a_23020_29890.n0 a_23020_29890.t8 228.148
R8044 a_23020_29890.t0 a_23020_29890.n5 221.411
R8045 a_23020_29890.n3 a_23020_29890.n0 209.601
R8046 a_23020_29890.n5 a_23020_29890.n3 207.974
R8047 a_23020_29890.n3 a_23020_29890.n2 123.35
R8048 a_23020_29890.n4 a_23020_29890.t1 24.0005
R8049 a_23020_29890.n4 a_23020_29890.t2 24.0005
R8050 a_23130_29970.t0 a_23130_29970.t1 48.0005
R8051 a_26300_23710.n4 a_26300_23710.t0 758.734
R8052 a_26300_23710.t1 a_26300_23710.n5 758.734
R8053 a_26300_23710.n0 a_26300_23710.t4 538.234
R8054 a_26300_23710.n3 a_26300_23710.n2 342.757
R8055 a_26300_23710.n5 a_26300_23710.t2 260.733
R8056 a_26300_23710.n3 a_26300_23710.t6 190.123
R8057 a_26300_23710.n4 a_26300_23710.n3 180.8
R8058 a_26300_23710.n0 a_26300_23710.t5 136.567
R8059 a_26300_23710.n1 a_26300_23710.t3 136.567
R8060 a_26300_23710.n2 a_26300_23710.t7 136.567
R8061 a_26300_23710.n1 a_26300_23710.n0 128.534
R8062 a_26300_23710.n2 a_26300_23710.n1 128.534
R8063 a_26300_23710.n5 a_26300_23710.n4 57.6005
R8064 a_13532_33810.t0 a_13532_33810.t1 258.591
R8065 a_14610_33690.t0 a_14610_33690.t1 258.591
R8066 a_24310_31910.t0 a_24310_31910.t1 39.4005
R8067 a_24310_27960.n0 a_24310_27960.t3 605.311
R8068 a_24310_27960.t1 a_24310_27960.n1 458.818
R8069 a_24310_27960.t1 a_24310_27960.n1 429.281
R8070 a_24310_27960.t3 a_24310_27960.t0 423.983
R8071 a_24310_27960.n0 a_24310_27960.t2 148.775
R8072 a_24310_27960.n1 a_24310_27960.n0 65.048
R8073 a_26390_29240.t1 a_26390_29240.n2 749.134
R8074 a_26390_29240.n2 a_26390_29240.t0 691.534
R8075 a_26390_29240.n1 a_26390_29240.n0 359.233
R8076 a_26390_29240.n1 a_26390_29240.t2 346.601
R8077 a_26390_29240.n0 a_26390_29240.t3 345.433
R8078 a_26390_29240.n0 a_26390_29240.t4 168.701
R8079 a_26390_29240.n2 a_26390_29240.n1 6.4005
R8080 a_19940_24230.t0 a_19940_24230.n6 1026.49
R8081 a_19940_24230.n3 a_19940_24230.n2 398.401
R8082 a_19940_24230.n2 a_19940_24230.n0 328.447
R8083 a_19940_24230.n2 a_19940_24230.n1 322.601
R8084 a_19940_24230.n4 a_19940_24230.t8 313.3
R8085 a_19940_24230.n5 a_19940_24230.t5 313.3
R8086 a_19940_24230.n6 a_19940_24230.t6 313.3
R8087 a_19940_24230.n3 a_19940_24230.t7 232.968
R8088 a_19940_24230.n4 a_19940_24230.n3 175.73
R8089 a_19940_24230.n5 a_19940_24230.n4 160.667
R8090 a_19940_24230.n6 a_19940_24230.n5 160.667
R8091 a_19940_24230.n1 a_19940_24230.t4 60.0005
R8092 a_19940_24230.n1 a_19940_24230.t3 60.0005
R8093 a_19940_24230.n0 a_19940_24230.t2 49.2505
R8094 a_19940_24230.n0 a_19940_24230.t1 49.2505
R8095 a_23550_31390.t0 a_23550_31390.t1 39.4005
R8096 a_26420_27330.t0 a_26420_27330.t1 96.0005
R8097 a_14610_33930.n6 a_14610_33930.t10 287.764
R8098 a_14610_33930.n5 a_14610_33930.t8 287.764
R8099 a_14610_33930.n5 a_14610_33930.t7 287.591
R8100 a_14610_33930.n8 a_14610_33930.t11 287.012
R8101 a_14610_33930.n7 a_14610_33930.t9 287.012
R8102 a_14610_33930.t0 a_14610_33930.n9 155.326
R8103 a_14610_33930.n2 a_14610_33930.n0 107.266
R8104 a_14610_33930.n4 a_14610_33930.n3 105.016
R8105 a_14610_33930.n2 a_14610_33930.n1 105.016
R8106 a_14610_33930.n3 a_14610_33930.t6 13.1338
R8107 a_14610_33930.n3 a_14610_33930.t4 13.1338
R8108 a_14610_33930.n1 a_14610_33930.t2 13.1338
R8109 a_14610_33930.n1 a_14610_33930.t3 13.1338
R8110 a_14610_33930.n0 a_14610_33930.t1 13.1338
R8111 a_14610_33930.n0 a_14610_33930.t5 13.1338
R8112 a_14610_33930.n9 a_14610_33930.n4 9.0005
R8113 a_14610_33930.n9 a_14610_33930.n8 6.78086
R8114 a_14610_33930.n4 a_14610_33930.n2 2.2505
R8115 a_14610_33930.n7 a_14610_33930.n6 0.579071
R8116 a_14610_33930.n8 a_14610_33930.n7 0.282643
R8117 a_14610_33930.n6 a_14610_33930.n5 0.2755
R8118 a_26420_29270.t0 a_26420_29270.t1 96.0005
R8119 a_26330_22330.t0 a_26330_22330.t1 96.0005
R8120 a_26390_27410.n1 a_26390_27410.t0 691
R8121 a_26390_27410.n1 a_26390_27410.n0 674.168
R8122 a_26390_27410.n0 a_26390_27410.t2 345.433
R8123 a_26390_27410.t1 a_26390_27410.n1 330.601
R8124 a_26390_27410.n0 a_26390_27410.t3 168.701
R8125 a_26420_29380.n0 a_26420_29380.t1 663.801
R8126 a_26420_29380.t0 a_26420_29380.n0 406.334
R8127 a_26420_29380.n0 a_26420_29380.t2 348.851
R8128 a_26330_23630.t0 a_26330_23630.t1 96.0005
R8129 a_26330_22440.n0 a_26330_22440.t0 713.933
R8130 a_26330_22440.t1 a_26330_22440.n0 337
R8131 a_26330_22440.n0 a_26330_22440.t2 314.233
R8132 a_23130_27960.n0 a_23130_27960.t2 496.889
R8133 a_23130_27960.t0 a_23130_27960.n2 458.818
R8134 a_23130_27960.t0 a_23130_27960.n2 429.281
R8135 a_23130_27960.n0 a_23130_27960.t3 393.634
R8136 a_23130_27960.n1 a_23130_27960.n0 384.967
R8137 a_23130_27960.n1 a_23130_27960.t1 177.576
R8138 a_23130_27960.n2 a_23130_27960.n1 34.648
R8139 a_26330_24930.t0 a_26330_24930.t1 96.0005
R8140 a_26330_23740.n0 a_26330_23740.t1 713.933
R8141 a_26330_23740.t0 a_26330_23740.n0 337
R8142 a_26330_23740.n0 a_26330_23740.t2 314.233
R8143 a_18460_22530.t0 a_18460_22530.t1 286.111
R8144 a_21386_22530.t0 a_21386_22530.t1 364.192
R8145 a_26420_31640.t0 a_26420_31640.t1 96.0005
R8146 a_23100_28450.t0 a_23100_28450.n2 458.818
R8147 a_23100_28450.n0 a_23100_28450.t2 441.834
R8148 a_23100_28450.t0 a_23100_28450.n2 429.281
R8149 a_23100_28450.n0 a_23100_28450.t3 313.3
R8150 a_23100_28450.n1 a_23100_28450.n0 228.8
R8151 a_23100_28450.n1 a_23100_28450.t1 174.375
R8152 a_23100_28450.n2 a_23100_28450.n1 50.648
R8153 a_23550_31010.t0 a_23550_31010.t1 39.4005
R8154 a_26330_25040.n0 a_26330_25040.t0 713.933
R8155 a_26330_25040.t1 a_26330_25040.n0 337
R8156 a_26330_25040.n0 a_26330_25040.t2 314.233
R8157 a_26420_31750.n0 a_26420_31750.t1 663.801
R8158 a_26420_31750.t0 a_26420_31750.n0 406.334
R8159 a_26420_31750.n0 a_26420_31750.t2 355.378
R8160 a_26420_30310.t0 a_26420_30310.t1 96.0005
R8161 a_25860_20560.n0 a_25860_20560.t0 284.2
R8162 a_25860_20560.n0 a_25860_20560.t2 233
R8163 a_25860_20560.t1 a_25860_20560.n0 184.191
R8164 a_24310_28480.t0 a_24310_28480.n2 458.818
R8165 a_24310_28480.t0 a_24310_28480.n2 429.281
R8166 a_24310_28480.n0 a_24310_28480.t3 256.428
R8167 a_24310_28480.n1 a_24310_28480.t1 190.375
R8168 a_24310_28480.n0 a_24310_28480.t2 190.375
R8169 a_24310_28480.n1 a_24310_28480.n0 70.4005
R8170 a_24310_28480.n2 a_24310_28480.n1 34.648
R8171 a_13382_33380.t0 a_13382_33380.t1 258.591
R8172 a_17540_28930.t0 a_17540_28930.t1 178.194
R8173 a_25860_21160.n0 a_25860_21160.t1 284.2
R8174 a_25860_21160.n0 a_25860_21160.t2 233
R8175 a_25860_21160.t0 a_25860_21160.n0 184.191
R8176 a_13382_28490.t0 a_13382_28490.t1 258.591
R8177 a_14990_28610.t0 a_14990_28610.t1 258.591
R8178 a_14990_33260.t0 a_14990_33260.t1 258.591
C0 uio_oe[6] uio_oe[5] 0.031023f
C1 uio_in[2] uio_in[1] 0.031023f
C2 uio_out[5] uio_out[4] 0.031023f
C3 uo_out[2] uo_out[1] 0.031023f
C4 uio_oe[0] uio_out[7] 0.031023f
C5 uio_in[7] uio_in[6] 0.031023f
C6 VGND ua[0] 0.410436f
C7 uo_out[7] uo_out[6] 0.031023f
C8 rst_n clk 0.031023f
C9 uio_oe[5] uio_oe[4] 0.031023f
C10 ui_in[4] ui_in[3] 0.031023f
C11 uio_in[1] uio_in[0] 0.031023f
C12 uio_out[4] uio_out[3] 0.031023f
C13 VGND ua[1] 0.708002f
C14 uio_out[7] uio_out[6] 0.031023f
C15 uio_in[6] uio_in[5] 0.031023f
C16 uo_out[6] uo_out[5] 0.031023f
C17 clk ena 0.031023f
C18 uio_oe[4] uio_oe[3] 0.031023f
C19 uio_in[0] ui_in[7] 0.031023f
C20 uio_out[3] uio_out[2] 0.031023f
C21 ui_in[3] ui_in[2] 0.031023f
C22 uio_in[5] uio_in[4] 0.031023f
C23 uo_out[0] uo_out[1] 0.031023f
C24 uo_out[5] uo_out[4] 0.031023f
C25 uio_oe[3] uio_oe[2] 0.031023f
C26 ui_in[7] ui_in[6] 0.031023f
C27 uio_out[2] uio_out[1] 0.031023f
C28 ui_in[2] ui_in[1] 0.031023f
C29 uio_in[4] uio_in[3] 0.031023f
C30 uio_out[6] uio_out[5] 0.031023f
C31 uo_out[4] uo_out[3] 0.031023f
C32 uio_oe[2] uio_oe[1] 0.031023f
C33 ui_in[6] ui_in[5] 0.031023f
C34 uio_out[1] uio_out[0] 0.031023f
C35 ui_in[1] ui_in[0] 0.031023f
C36 uio_oe[7] uio_oe[6] 0.031023f
C37 uio_in[3] uio_in[2] 0.031023f
C38 uo_out[3] uo_out[2] 0.031023f
C39 uio_oe[1] uio_oe[0] 0.031023f
C40 uo_out[0] uio_in[7] 0.031023f
C41 ui_in[5] ui_in[4] 0.031023f
C42 uio_out[0] uo_out[7] 0.031023f
C43 ui_in[0] rst_n 0.031023f
C44 ua[2] VDPWR 0.146962f
C45 ua[3] VDPWR 0.146962f
C46 ua[4] VDPWR 0.146962f
C47 ua[5] VDPWR 0.146962f
C48 ua[6] VDPWR 0.146962f
C49 ua[7] VDPWR 0.146962f
C50 ena VDPWR 0.070385f
C51 clk VDPWR 0.042875f
C52 rst_n VDPWR 0.042875f
C53 ui_in[0] VDPWR 0.042875f
C54 ui_in[1] VDPWR 0.042875f
C55 ui_in[2] VDPWR 0.042875f
C56 ui_in[3] VDPWR 0.042875f
C57 ui_in[4] VDPWR 0.042875f
C58 ui_in[5] VDPWR 0.042875f
C59 ui_in[6] VDPWR 0.042875f
C60 ui_in[7] VDPWR 0.042875f
C61 uio_in[0] VDPWR 0.042875f
C62 uio_in[1] VDPWR 0.042875f
C63 uio_in[2] VDPWR 0.042875f
C64 uio_in[3] VDPWR 0.042875f
C65 uio_in[4] VDPWR 0.042875f
C66 uio_in[5] VDPWR 0.042875f
C67 uio_in[6] VDPWR 0.042875f
C68 uio_in[7] VDPWR 0.042875f
C69 uo_out[0] VDPWR 0.042875f
C70 uo_out[1] VDPWR 0.042875f
C71 uo_out[2] VDPWR 0.042875f
C72 uo_out[3] VDPWR 0.042875f
C73 uo_out[4] VDPWR 0.042875f
C74 uo_out[5] VDPWR 0.042875f
C75 uo_out[6] VDPWR 0.042875f
C76 uo_out[7] VDPWR 0.042875f
C77 uio_out[0] VDPWR 0.042875f
C78 uio_out[1] VDPWR 0.042875f
C79 uio_out[2] VDPWR 0.042875f
C80 uio_out[3] VDPWR 0.042875f
C81 uio_out[4] VDPWR 0.042875f
C82 uio_out[5] VDPWR 0.042875f
C83 uio_out[6] VDPWR 0.042875f
C84 uio_out[7] VDPWR 0.042875f
C85 uio_oe[0] VDPWR 0.042875f
C86 uio_oe[1] VDPWR 0.042875f
C87 uio_oe[2] VDPWR 0.042875f
C88 uio_oe[3] VDPWR 0.042875f
C89 uio_oe[4] VDPWR 0.042875f
C90 uio_oe[5] VDPWR 0.042875f
C91 uio_oe[6] VDPWR 0.042875f
C92 uio_oe[7] VDPWR 0.070385f
C93 ua[1] VDPWR 11.0531f
C94 ua[0] VDPWR 17.6488f
C95 VGND VDPWR 0.134561p
C96 a_23130_27960.t1 VDPWR 0.026996f
C97 a_23130_27960.t2 VDPWR 2.01377f
C98 a_23130_27960.t3 VDPWR 0.010471f
C99 a_23130_27960.n0 VDPWR 0.029667f
C100 a_23130_27960.n1 VDPWR 0.037413f
C101 a_23130_27960.n2 VDPWR 0.046542f
C102 a_23130_27960.t0 VDPWR 0.03514f
C103 a_14610_33930.t1 VDPWR 0.10095f
C104 a_14610_33930.t5 VDPWR 0.10095f
C105 a_14610_33930.n0 VDPWR 0.2816f
C106 a_14610_33930.t2 VDPWR 0.10095f
C107 a_14610_33930.t3 VDPWR 0.10095f
C108 a_14610_33930.n1 VDPWR 0.253459f
C109 a_14610_33930.n2 VDPWR 3.1126f
C110 a_14610_33930.t6 VDPWR 0.10095f
C111 a_14610_33930.t4 VDPWR 0.10095f
C112 a_14610_33930.n3 VDPWR 0.253459f
C113 a_14610_33930.n4 VDPWR 2.34993f
C114 a_14610_33930.t7 VDPWR 0.055705f
C115 a_14610_33930.t8 VDPWR 0.05457f
C116 a_14610_33930.n5 VDPWR 0.425181f
C117 a_14610_33930.t10 VDPWR 0.05457f
C118 a_14610_33930.n6 VDPWR 0.226996f
C119 a_14610_33930.t9 VDPWR 0.055305f
C120 a_14610_33930.n7 VDPWR 0.228617f
C121 a_14610_33930.t11 VDPWR 0.055305f
C122 a_14610_33930.n8 VDPWR 0.780841f
C123 a_14610_33930.n9 VDPWR 4.14023f
C124 a_14610_33930.t0 VDPWR 0.365925f
C125 a_13742_34050.t5 VDPWR 0.293845f
C126 a_13742_34050.t12 VDPWR 0.309615f
C127 a_13742_34050.t6 VDPWR 0.309615f
C128 a_13742_34050.t14 VDPWR 0.309615f
C129 a_13742_34050.t18 VDPWR 0.309615f
C130 a_13742_34050.t1 VDPWR 0.309615f
C131 a_13742_34050.t19 VDPWR 0.309615f
C132 a_13742_34050.t3 VDPWR 0.309615f
C133 a_13742_34050.t9 VDPWR 0.29491f
C134 a_13742_34050.t4 VDPWR 0.14206f
C135 a_13742_34050.n0 VDPWR 0.183237f
C136 a_13742_34050.t10 VDPWR 0.322105f
C137 a_13742_34050.t15 VDPWR 0.296149f
C138 a_13742_34050.t8 VDPWR 0.309615f
C139 a_13742_34050.t2 VDPWR 0.309615f
C140 a_13742_34050.t7 VDPWR 0.309615f
C141 a_13742_34050.t0 VDPWR 0.309615f
C142 a_13742_34050.t17 VDPWR 0.309615f
C143 a_13742_34050.t13 VDPWR 0.309615f
C144 a_13742_34050.t16 VDPWR 0.309615f
C145 a_13742_34050.t11 VDPWR 1.1782f
C146 a_13742_34050.t20 VDPWR 0.154879f
C147 a_25350_8708.t1 VDPWR 2.39855f
C148 a_14140_28370.t8 VDPWR 0.021628f
C149 a_14140_28370.t2 VDPWR 0.021628f
C150 a_14140_28370.n0 VDPWR 0.047663f
C151 a_14140_28370.t10 VDPWR 0.021628f
C152 a_14140_28370.t3 VDPWR 0.021628f
C153 a_14140_28370.n1 VDPWR 0.047367f
C154 a_14140_28370.n2 VDPWR 0.55165f
C155 a_14140_28370.t12 VDPWR 0.021628f
C156 a_14140_28370.t6 VDPWR 0.021628f
C157 a_14140_28370.n3 VDPWR 0.047367f
C158 a_14140_28370.n4 VDPWR 0.291113f
C159 a_14140_28370.t4 VDPWR 0.021628f
C160 a_14140_28370.t9 VDPWR 0.021628f
C161 a_14140_28370.n5 VDPWR 0.047367f
C162 a_14140_28370.n6 VDPWR 0.291113f
C163 a_14140_28370.t7 VDPWR 0.021628f
C164 a_14140_28370.t11 VDPWR 0.021628f
C165 a_14140_28370.n7 VDPWR 0.047367f
C166 a_14140_28370.n8 VDPWR 0.291113f
C167 a_14140_28370.t1 VDPWR 0.021628f
C168 a_14140_28370.t5 VDPWR 0.021628f
C169 a_14140_28370.n9 VDPWR 0.047367f
C170 a_14140_28370.n10 VDPWR 1.14445f
C171 a_14140_28370.t13 VDPWR 0.033253f
C172 a_14140_28370.t14 VDPWR 0.033188f
C173 a_14140_28370.n11 VDPWR 0.233433f
C174 a_14140_28370.t16 VDPWR 0.033188f
C175 a_14140_28370.n12 VDPWR 0.145136f
C176 a_14140_28370.t15 VDPWR 0.033188f
C177 a_14140_28370.n13 VDPWR 0.145136f
C178 a_14140_28370.t17 VDPWR 0.033188f
C179 a_14140_28370.n14 VDPWR 0.4804f
C180 a_14140_28370.n15 VDPWR 5.4833f
C181 a_14140_28370.t0 VDPWR 0.533116f
C182 a_22190_29430.n0 VDPWR 0.156934f
C183 a_22190_29430.n1 VDPWR 0.118238f
C184 a_22190_29430.t4 VDPWR 0.029882f
C185 a_22190_29430.t5 VDPWR 0.031397f
C186 a_22190_29430.n2 VDPWR 0.067221f
C187 a_22190_29430.t3 VDPWR 0.010639f
C188 a_22190_29430.t1 VDPWR 0.010639f
C189 a_22190_29430.n3 VDPWR 0.041426f
C190 a_22190_29430.t2 VDPWR 0.049455f
C191 a_22190_29430.t19 VDPWR 0.062085f
C192 a_22190_29430.t18 VDPWR 0.04628f
C193 a_22190_29430.n4 VDPWR 0.046455f
C194 a_22190_29430.n5 VDPWR 0.048543f
C195 a_22190_29430.t0 VDPWR 0.03365f
C196 a_22190_29430.n6 VDPWR 0.040235f
C197 a_22190_29430.n7 VDPWR 0.04416f
C198 a_22190_29430.n8 VDPWR 1.61807f
C199 a_22190_29430.n9 VDPWR 1.98317f
C200 a_22190_29430.n11 VDPWR 0.060082f
C201 a_22190_29430.n12 VDPWR 0.018725f
C202 a_22190_29430.n14 VDPWR 0.062631f
C203 a_22190_29430.n16 VDPWR 0.030586f
C204 a_22190_29430.n17 VDPWR 0.059176f
C205 a_22190_29430.n19 VDPWR 0.059176f
C206 a_22190_29430.n21 VDPWR 0.059176f
C207 a_22190_29430.n22 VDPWR 0.018725f
C208 a_22190_29430.n23 VDPWR 0.030586f
C209 a_22190_29430.n24 VDPWR 0.059176f
C210 a_14558_34050.t25 VDPWR 0.049701f
C211 a_14558_34050.t12 VDPWR 0.049641f
C212 a_14558_34050.n0 VDPWR 0.259633f
C213 a_14558_34050.t19 VDPWR 0.049641f
C214 a_14558_34050.n1 VDPWR 0.136128f
C215 a_14558_34050.t28 VDPWR 0.049641f
C216 a_14558_34050.n2 VDPWR 0.136128f
C217 a_14558_34050.t15 VDPWR 0.049641f
C218 a_14558_34050.n3 VDPWR 0.136128f
C219 a_14558_34050.t13 VDPWR 0.049641f
C220 a_14558_34050.n4 VDPWR 0.136128f
C221 a_14558_34050.t22 VDPWR 0.049641f
C222 a_14558_34050.n5 VDPWR 0.136128f
C223 a_14558_34050.t10 VDPWR 0.049641f
C224 a_14558_34050.n6 VDPWR 0.136128f
C225 a_14558_34050.t17 VDPWR 0.049641f
C226 a_14558_34050.n7 VDPWR 0.136128f
C227 a_14558_34050.t21 VDPWR 0.049641f
C228 a_14558_34050.n8 VDPWR 0.337114f
C229 a_14558_34050.t20 VDPWR 0.049641f
C230 a_14558_34050.n9 VDPWR 0.337114f
C231 a_14558_34050.t29 VDPWR 0.049641f
C232 a_14558_34050.n10 VDPWR 0.136128f
C233 a_14558_34050.t16 VDPWR 0.049641f
C234 a_14558_34050.n11 VDPWR 0.136128f
C235 a_14558_34050.t24 VDPWR 0.049641f
C236 a_14558_34050.n12 VDPWR 0.136128f
C237 a_14558_34050.t11 VDPWR 0.049641f
C238 a_14558_34050.n13 VDPWR 0.136128f
C239 a_14558_34050.t18 VDPWR 0.049641f
C240 a_14558_34050.n14 VDPWR 0.136128f
C241 a_14558_34050.t27 VDPWR 0.049641f
C242 a_14558_34050.n15 VDPWR 0.136128f
C243 a_14558_34050.t14 VDPWR 0.049641f
C244 a_14558_34050.n16 VDPWR 0.136128f
C245 a_14558_34050.t23 VDPWR 0.049641f
C246 a_14558_34050.n17 VDPWR 0.136128f
C247 a_14558_34050.t26 VDPWR 0.049641f
C248 a_14558_34050.n18 VDPWR 0.992373f
C249 a_14558_34050.t2 VDPWR 0.434311f
C250 a_14558_34050.t3 VDPWR 0.028712f
C251 a_14558_34050.t0 VDPWR 0.028712f
C252 a_14558_34050.n19 VDPWR 0.062021f
C253 a_14558_34050.n20 VDPWR 1.41734f
C254 a_14558_34050.t7 VDPWR 0.028712f
C255 a_14558_34050.t8 VDPWR 0.028712f
C256 a_14558_34050.n21 VDPWR 0.062021f
C257 a_14558_34050.n22 VDPWR 0.627074f
C258 a_14558_34050.t5 VDPWR 0.028712f
C259 a_14558_34050.t6 VDPWR 0.028712f
C260 a_14558_34050.n23 VDPWR 0.062021f
C261 a_14558_34050.n24 VDPWR 0.614154f
C262 a_14558_34050.t1 VDPWR 0.028712f
C263 a_14558_34050.t4 VDPWR 0.028712f
C264 a_14558_34050.n25 VDPWR 0.062021f
C265 a_14558_34050.n26 VDPWR 0.715576f
C266 a_14558_34050.n27 VDPWR 4.21165f
C267 a_14558_34050.t9 VDPWR 0.341077f
C268 a_19910_24460.n5 VDPWR 0.058699f
C269 a_19910_24460.n9 VDPWR 0.017948f
C270 a_19910_24460.n10 VDPWR 0.014992f
C271 a_19910_24460.n11 VDPWR 0.082942f
C272 a_19910_24460.n12 VDPWR 0.02022f
C273 a_19910_24460.t7 VDPWR 6.66862f
C274 a_19910_24460.n13 VDPWR 0.162298f
C275 a_19910_24460.t0 VDPWR 0.019038f
C276 a_23100_30050.t2 VDPWR 0.027951f
C277 a_23100_30050.t0 VDPWR 0.027951f
C278 a_23100_30050.n0 VDPWR 0.149246f
C279 a_23100_30050.t3 VDPWR 0.030633f
C280 a_23100_30050.t8 VDPWR 0.069862f
C281 a_23100_30050.n1 VDPWR 0.179221f
C282 a_23100_30050.t7 VDPWR 0.034065f
C283 a_23100_30050.t6 VDPWR 0.070751f
C284 a_23100_30050.n2 VDPWR 0.099239f
C285 a_23100_30050.t5 VDPWR 0.069179f
C286 a_23100_30050.t4 VDPWR 0.104293f
C287 a_23100_30050.n3 VDPWR 1.26639f
C288 a_23100_30050.n4 VDPWR 0.267564f
C289 a_23100_30050.n5 VDPWR 0.256539f
C290 a_23100_30050.t1 VDPWR 0.147114f
C291 a_14990_33500.t5 VDPWR 0.051177f
C292 a_14990_33500.t4 VDPWR 0.051177f
C293 a_14990_33500.n0 VDPWR 0.127305f
C294 a_14990_33500.t3 VDPWR 0.051177f
C295 a_14990_33500.t2 VDPWR 0.051177f
C296 a_14990_33500.n1 VDPWR 0.122339f
C297 a_14990_33500.n2 VDPWR 1.74488f
C298 a_14990_33500.t6 VDPWR 0.026228f
C299 a_14990_33500.t10 VDPWR 0.026177f
C300 a_14990_33500.n3 VDPWR 0.184117f
C301 a_14990_33500.t8 VDPWR 0.026177f
C302 a_14990_33500.n4 VDPWR 0.114474f
C303 a_14990_33500.t9 VDPWR 0.026177f
C304 a_14990_33500.n5 VDPWR 0.114474f
C305 a_14990_33500.t7 VDPWR 0.026177f
C306 a_14990_33500.n6 VDPWR 0.383297f
C307 a_14990_33500.n7 VDPWR 0.903315f
C308 a_14990_33500.t1 VDPWR 0.191955f
C309 a_14990_33500.n8 VDPWR 2.2109f
C310 a_14990_33500.t0 VDPWR 0.267299f
C311 a_17540_31010.t4 VDPWR 0.04324f
C312 a_17540_31010.t0 VDPWR 1.74484f
C313 a_17540_31010.t1 VDPWR 0.045667f
C314 a_17540_31010.n0 VDPWR 1.57161f
C315 a_17540_31010.t7 VDPWR 0.016248f
C316 a_17540_31010.t6 VDPWR 0.016248f
C317 a_17540_31010.n1 VDPWR 0.053414f
C318 a_17540_31010.t3 VDPWR 0.04324f
C319 a_17540_31010.t2 VDPWR 0.04324f
C320 a_17540_31010.n2 VDPWR 0.106515f
C321 a_17540_31010.n3 VDPWR 1.2172f
C322 a_17540_31010.n4 VDPWR 2.04879f
C323 a_17540_31010.n5 VDPWR 0.106515f
C324 a_17540_31010.t5 VDPWR 0.04324f
C325 a_19190_29290.t9 VDPWR 0.018056f
C326 a_19190_29290.t1 VDPWR 0.018056f
C327 a_19190_29290.t7 VDPWR 0.018056f
C328 a_19190_29290.n0 VDPWR 0.036969f
C329 a_19190_29290.t0 VDPWR 0.021667f
C330 a_19190_29290.t20 VDPWR 0.021667f
C331 a_19190_29290.t21 VDPWR 0.034973f
C332 a_19190_29290.n1 VDPWR 0.039055f
C333 a_19190_29290.n2 VDPWR 0.02668f
C334 a_19190_29290.t6 VDPWR 0.027505f
C335 a_19190_29290.n3 VDPWR 0.043175f
C336 a_19190_29290.n4 VDPWR 0.191386f
C337 a_19190_29290.t3 VDPWR 0.018056f
C338 a_19190_29290.t5 VDPWR 0.018056f
C339 a_19190_29290.n5 VDPWR 0.036969f
C340 a_19190_29290.t2 VDPWR 0.021667f
C341 a_19190_29290.t22 VDPWR 0.021667f
C342 a_19190_29290.t17 VDPWR 0.034973f
C343 a_19190_29290.n6 VDPWR 0.039055f
C344 a_19190_29290.n7 VDPWR 0.02668f
C345 a_19190_29290.t4 VDPWR 0.027505f
C346 a_19190_29290.n8 VDPWR 0.043175f
C347 a_19190_29290.n9 VDPWR 0.191386f
C348 a_19190_29290.n10 VDPWR 0.26218f
C349 a_19190_29290.n11 VDPWR 0.019256f
C350 a_19190_29290.t15 VDPWR 0.034183f
C351 a_19190_29290.n12 VDPWR 0.021429f
C352 a_19190_29290.n13 VDPWR 0.554666f
C353 a_19190_29290.n14 VDPWR 0.186578f
C354 a_19190_29290.t8 VDPWR 0.021667f
C355 a_19190_29290.t19 VDPWR 0.021667f
C356 a_19190_29290.t18 VDPWR 0.034973f
C357 a_19190_29290.n15 VDPWR 0.039055f
C358 a_19190_29290.n16 VDPWR 0.02668f
C359 a_19190_29290.t10 VDPWR 0.027505f
C360 a_19190_29290.n17 VDPWR 0.043175f
C361 a_19190_29290.n18 VDPWR 0.239421f
C362 a_19190_29290.n19 VDPWR 0.036969f
C363 a_19190_29290.t11 VDPWR 0.018056f
C364 a_19940_23090.n3 VDPWR 0.01467f
C365 a_19940_23090.t13 VDPWR 1.08371f
C366 a_19940_23090.t3 VDPWR 0.011718f
C367 a_19940_23090.n5 VDPWR 0.020093f
C368 a_19940_23090.t14 VDPWR 0.014564f
C369 a_19940_23090.t15 VDPWR 0.01094f
C370 a_19940_23090.n11 VDPWR 0.103723f
C371 a_19940_23090.n12 VDPWR 0.053506f
C372 a_19940_23090.t12 VDPWR 1.08411f
C373 a_19940_23090.n14 VDPWR 0.010922f
C374 a_13532_27710.t10 VDPWR 0.31433f
C375 a_13532_27710.t17 VDPWR 0.331199f
C376 a_13532_27710.t11 VDPWR 0.331199f
C377 a_13532_27710.t19 VDPWR 0.331199f
C378 a_13532_27710.t3 VDPWR 0.331199f
C379 a_13532_27710.t6 VDPWR 0.331199f
C380 a_13532_27710.t4 VDPWR 0.331199f
C381 a_13532_27710.t8 VDPWR 0.331199f
C382 a_13532_27710.t14 VDPWR 0.315469f
C383 a_13532_27710.t9 VDPWR 0.151964f
C384 a_13532_27710.n0 VDPWR 0.19601f
C385 a_13532_27710.t15 VDPWR 0.344559f
C386 a_13532_27710.t20 VDPWR 0.316794f
C387 a_13532_27710.t13 VDPWR 0.331199f
C388 a_13532_27710.t7 VDPWR 0.331199f
C389 a_13532_27710.t12 VDPWR 0.331199f
C390 a_13532_27710.t5 VDPWR 0.331199f
C391 a_13532_27710.t2 VDPWR 0.331199f
C392 a_13532_27710.t18 VDPWR 0.331199f
C393 a_13532_27710.t1 VDPWR 0.331199f
C394 a_13532_27710.t16 VDPWR 0.743991f
C395 a_13532_27710.t0 VDPWR 0.080098f
C396 a_17884_25798.t3 VDPWR 0.019014f
C397 a_17884_25798.t7 VDPWR 0.019014f
C398 a_17884_25798.n0 VDPWR 0.052203f
C399 a_17884_25798.t1 VDPWR 0.019014f
C400 a_17884_25798.t5 VDPWR 0.019014f
C401 a_17884_25798.n1 VDPWR 0.053666f
C402 a_17884_25798.n2 VDPWR 0.065336f
C403 a_17884_25798.t2 VDPWR 0.052478f
C404 a_17884_25798.t12 VDPWR 0.052478f
C405 a_17884_25798.t10 VDPWR 0.072156f
C406 a_17884_25798.n3 VDPWR 0.040407f
C407 a_17884_25798.n4 VDPWR 0.028673f
C408 a_17884_25798.t6 VDPWR 0.052478f
C409 a_17884_25798.t0 VDPWR 0.052478f
C410 a_17884_25798.t4 VDPWR 0.052478f
C411 a_17884_25798.t9 VDPWR 0.052478f
C412 a_17884_25798.t11 VDPWR 0.072156f
C413 a_17884_25798.n5 VDPWR 0.040407f
C414 a_17884_25798.n6 VDPWR 0.028673f
C415 a_17884_25798.n7 VDPWR 0.012378f
C416 a_17884_25798.n8 VDPWR 0.028673f
C417 a_17884_25798.n9 VDPWR 0.028673f
C418 a_17884_25798.n10 VDPWR 0.012321f
C419 a_17884_25798.n11 VDPWR 0.209105f
C420 a_17884_25798.t8 VDPWR 1.66425f
C421 w_20440_23530.n1 VDPWR 0.069381f
C422 w_20440_23530.n2 VDPWR 0.067052f
C423 w_20440_23530.n4 VDPWR 0.0681f
C424 w_20440_23530.n6 VDPWR 0.0681f
C425 w_20440_23530.n8 VDPWR 0.0681f
C426 w_20440_23530.n13 VDPWR 0.013149f
C427 w_20440_23530.n14 VDPWR 0.013149f
C428 w_20440_23530.t48 VDPWR 0.013103f
C429 w_20440_23530.n16 VDPWR 0.03259f
C430 w_20440_23530.t57 VDPWR 0.013103f
C431 w_20440_23530.n17 VDPWR 0.03259f
C432 w_20440_23530.t52 VDPWR 0.013103f
C433 w_20440_23530.n18 VDPWR 0.03259f
C434 w_20440_23530.t41 VDPWR 0.013103f
C435 w_20440_23530.n21 VDPWR 0.0161f
C436 w_20440_23530.n23 VDPWR 0.019123f
C437 w_20440_23530.n25 VDPWR 0.019123f
C438 w_20440_23530.n27 VDPWR 0.019123f
C439 w_20440_23530.n29 VDPWR 0.019123f
C440 w_20440_23530.n30 VDPWR 0.01395f
C441 w_20440_23530.t42 VDPWR 0.036185f
C442 w_20440_23530.n31 VDPWR 0.014871f
C443 w_20440_23530.n32 VDPWR 0.019123f
C444 w_20440_23530.n49 VDPWR 0.0161f
C445 w_20440_23530.n53 VDPWR 0.0161f
C446 w_20440_23530.n54 VDPWR 0.020191f
C447 w_20440_23530.n60 VDPWR 0.066005f
C448 w_20440_23530.n61 VDPWR 0.066111f
C449 w_20440_23530.n63 VDPWR 0.021967f
C450 w_20440_23530.n65 VDPWR 0.0161f
C451 w_20440_23530.n67 VDPWR 0.100347f
C452 w_20440_23530.t39 VDPWR 0.245913f
C453 w_20440_23530.t22 VDPWR 0.124407f
C454 w_20440_23530.t20 VDPWR 0.124407f
C455 w_20440_23530.t6 VDPWR 0.124407f
C456 w_20440_23530.t10 VDPWR 0.124407f
C457 w_20440_23530.t51 VDPWR 0.141154f
C458 w_20440_23530.n68 VDPWR 0.091173f
C459 w_20440_23530.n72 VDPWR 0.013149f
C460 w_20440_23530.n74 VDPWR 0.013149f
C461 w_20440_23530.n77 VDPWR 0.013149f
C462 w_20440_23530.t58 VDPWR 0.036926f
C463 w_20440_23530.n78 VDPWR 0.025802f
C464 w_20440_23530.n79 VDPWR 0.027394f
C465 w_20440_23530.n80 VDPWR 0.011613f
C466 w_20440_23530.n82 VDPWR 0.075462f
C467 w_20440_23530.n83 VDPWR 0.093273f
C468 w_20440_23530.t59 VDPWR 0.07895f
C469 w_20440_23530.t55 VDPWR 0.095697f
C470 w_20440_23530.t36 VDPWR 0.062203f
C471 w_20440_23530.t0 VDPWR 0.083735f
C472 w_20440_23530.t24 VDPWR 0.074165f
C473 w_20440_23530.t32 VDPWR 0.062203f
C474 w_20440_23530.t30 VDPWR 0.095697f
C475 w_20440_23530.t2 VDPWR 0.062203f
C476 w_20440_23530.t8 VDPWR 0.07895f
C477 w_20440_23530.t47 VDPWR 0.07895f
C478 w_20440_23530.t16 VDPWR 0.07895f
C479 w_20440_23530.n84 VDPWR 0.103135f
C480 w_20440_23530.t14 VDPWR 0.129191f
C481 w_20440_23530.t18 VDPWR 0.122014f
C482 w_20440_23530.t26 VDPWR 0.08852f
C483 w_20440_23530.t28 VDPWR 0.069381f
C484 w_20440_23530.t12 VDPWR 0.062203f
C485 w_20440_23530.t29 VDPWR 0.095697f
C486 w_20440_23530.t34 VDPWR 0.062203f
C487 w_20440_23530.t4 VDPWR 0.083735f
C488 w_20440_23530.t5 VDPWR 0.074165f
C489 w_20440_23530.t43 VDPWR 0.062203f
C490 w_20440_23530.t27 VDPWR 0.095697f
C491 w_20440_23530.n85 VDPWR 0.198572f
C492 w_20440_23530.n88 VDPWR 0.013149f
C493 w_20440_23530.n89 VDPWR 0.013271f
C494 w_20440_23530.n90 VDPWR 0.027394f
C495 a_20480_25210.t5 VDPWR 0.078785f
C496 a_20480_25210.t3 VDPWR 0.030346f
C497 a_20480_25210.n0 VDPWR 0.120193f
C498 a_20480_25210.t9 VDPWR 0.020046f
C499 a_20480_25210.t4 VDPWR 0.020046f
C500 a_20480_25210.n1 VDPWR 0.046f
C501 a_20480_25210.n2 VDPWR 0.087576f
C502 a_20480_25210.t11 VDPWR 0.050114f
C503 a_20480_25210.t13 VDPWR 0.050114f
C504 a_20480_25210.n3 VDPWR 0.291421f
C505 a_20480_25210.t12 VDPWR 0.050114f
C506 a_20480_25210.t2 VDPWR 0.050114f
C507 a_20480_25210.n4 VDPWR 0.1426f
C508 a_20480_25210.n5 VDPWR 0.355827f
C509 a_20480_25210.n6 VDPWR 0.128581f
C510 a_20480_25210.t0 VDPWR 0.020046f
C511 a_20480_25210.t10 VDPWR 0.020046f
C512 a_20480_25210.n7 VDPWR 0.045548f
C513 a_20480_25210.n8 VDPWR 0.08916f
C514 a_20480_25210.t8 VDPWR 0.020046f
C515 a_20480_25210.t1 VDPWR 0.020046f
C516 a_20480_25210.n9 VDPWR 0.045548f
C517 a_20480_25210.n10 VDPWR 0.088358f
C518 a_20480_25210.t6 VDPWR 0.030346f
C519 a_20480_25210.n11 VDPWR 0.120193f
C520 a_20480_25210.t7 VDPWR 0.078785f
C521 a_14730_30630.t7 VDPWR 3.38919f
C522 a_14730_30630.t6 VDPWR 0.044358f
C523 a_14730_30630.t5 VDPWR 0.044358f
C524 a_14730_30630.n0 VDPWR 0.118669f
C525 a_14730_30630.t3 VDPWR 0.044358f
C526 a_14730_30630.t4 VDPWR 0.044358f
C527 a_14730_30630.n1 VDPWR 0.107634f
C528 a_14730_30630.n2 VDPWR 1.21683f
C529 a_14730_30630.t1 VDPWR 0.014786f
C530 a_14730_30630.t2 VDPWR 0.014786f
C531 a_14730_30630.n3 VDPWR 0.041682f
C532 a_14730_30630.n4 VDPWR 0.860437f
C533 a_14730_30630.t8 VDPWR 0.024477f
C534 a_14730_30630.t12 VDPWR 0.023979f
C535 a_14730_30630.n5 VDPWR 0.186829f
C536 a_14730_30630.t10 VDPWR 0.023979f
C537 a_14730_30630.n6 VDPWR 0.099745f
C538 a_14730_30630.t11 VDPWR 0.024302f
C539 a_14730_30630.n7 VDPWR 0.100457f
C540 a_14730_30630.t9 VDPWR 0.024302f
C541 a_14730_30630.n8 VDPWR 0.343109f
C542 a_14730_30630.n9 VDPWR 0.545948f
C543 a_14730_30630.n10 VDPWR 3.51458f
C544 a_14730_30630.t0 VDPWR 0.146843f
C545 a_25860_20180.t2 VDPWR 0.104706f
C546 a_25860_20180.n0 VDPWR 0.184398f
C547 a_25860_20180.t4 VDPWR 0.298444f
C548 a_25860_20180.t5 VDPWR 0.298444f
C549 a_25860_20180.t3 VDPWR 0.497217f
C550 a_25860_20180.n1 VDPWR 0.243367f
C551 a_25860_20180.n2 VDPWR 0.217957f
C552 a_25860_20180.t1 VDPWR 0.298444f
C553 a_25860_20180.n3 VDPWR 0.169192f
C554 a_25860_20180.n4 VDPWR 0.045341f
C555 a_25860_20180.n5 VDPWR 0.177419f
C556 a_25860_20180.t0 VDPWR 0.165068f
C557 a_19190_31850.n0 VDPWR 0.454298f
C558 a_19190_31850.n1 VDPWR 0.360667f
C559 a_19190_31850.n2 VDPWR 0.360667f
C560 a_19190_31850.n3 VDPWR 0.541f
C561 a_19190_31850.n4 VDPWR 0.360667f
C562 a_19190_31850.n5 VDPWR 0.360667f
C563 a_19190_31850.n6 VDPWR 0.360667f
C564 a_19190_31850.n7 VDPWR 0.360667f
C565 a_19190_31850.n8 VDPWR 1.23776f
C566 a_19190_31850.t8 VDPWR 0.010305f
C567 a_19190_31850.t25 VDPWR 0.0244f
C568 a_19190_31850.t31 VDPWR 0.41219f
C569 a_19190_31850.t23 VDPWR 0.419031f
C570 a_19190_31850.t16 VDPWR 0.41219f
C571 a_19190_31850.t21 VDPWR 0.41219f
C572 a_19190_31850.t15 VDPWR 0.41219f
C573 a_19190_31850.t36 VDPWR 0.41219f
C574 a_19190_31850.t28 VDPWR 0.41219f
C575 a_19190_31850.t34 VDPWR 0.41219f
C576 a_19190_31850.t27 VDPWR 0.41219f
C577 a_19190_31850.t18 VDPWR 0.41219f
C578 a_19190_31850.t24 VDPWR 0.41219f
C579 a_19190_31850.t26 VDPWR 0.41219f
C580 a_19190_31850.t33 VDPWR 0.41219f
C581 a_19190_31850.t13 VDPWR 0.41219f
C582 a_19190_31850.t35 VDPWR 0.41219f
C583 a_19190_31850.t14 VDPWR 0.41219f
C584 a_19190_31850.t20 VDPWR 0.41219f
C585 a_19190_31850.t29 VDPWR 0.41219f
C586 a_19190_31850.t22 VDPWR 0.41219f
C587 a_19190_31850.t30 VDPWR 0.41219f
C588 a_19190_31850.n9 VDPWR 0.949842f
C589 a_19190_31850.t4 VDPWR 0.010305f
C590 a_19190_31850.t5 VDPWR 0.010305f
C591 a_19190_31850.n10 VDPWR 0.022597f
C592 a_19190_31850.n11 VDPWR 0.215358f
C593 a_19190_31850.t19 VDPWR 0.015954f
C594 a_19190_31850.t17 VDPWR 0.015954f
C595 a_19190_31850.n12 VDPWR 0.029642f
C596 a_19190_31850.t3 VDPWR 0.018148f
C597 a_19190_31850.n13 VDPWR 0.013021f
C598 a_19190_31850.n14 VDPWR 0.012563f
C599 a_19190_31850.n15 VDPWR 0.335083f
C600 a_19190_31850.n16 VDPWR 0.110146f
C601 a_19190_31850.n17 VDPWR 0.06623f
C602 a_19190_31850.n18 VDPWR 0.074194f
C603 a_19190_31850.t7 VDPWR 0.010305f
C604 a_19190_31850.t6 VDPWR 0.010305f
C605 a_19190_31850.n19 VDPWR 0.022597f
C606 a_19190_31850.n20 VDPWR 0.169072f
C607 a_19190_31850.t12 VDPWR 0.015954f
C608 a_19190_31850.t11 VDPWR 0.015954f
C609 a_19190_31850.n21 VDPWR 0.030906f
C610 a_19190_31850.n22 VDPWR 0.119581f
C611 a_19190_31850.t32 VDPWR 0.024727f
C612 a_19190_31850.n23 VDPWR 0.245331f
C613 a_19190_31850.n24 VDPWR 0.022597f
C614 a_19190_31850.t9 VDPWR 0.010305f
C615 a_19190_31610.t13 VDPWR 0.016667f
C616 a_19190_31610.t9 VDPWR 0.016667f
C617 a_19190_31610.t11 VDPWR 0.016667f
C618 a_19190_31610.n0 VDPWR 0.034125f
C619 a_19190_31610.t8 VDPWR 0.025389f
C620 a_19190_31610.t10 VDPWR 0.02f
C621 a_19190_31610.t22 VDPWR 0.02f
C622 a_19190_31610.t21 VDPWR 0.032283f
C623 a_19190_31610.n1 VDPWR 0.036051f
C624 a_19190_31610.n2 VDPWR 0.024627f
C625 a_19190_31610.n3 VDPWR 0.039854f
C626 a_19190_31610.n4 VDPWR 0.176664f
C627 a_19190_31610.t5 VDPWR 0.016667f
C628 a_19190_31610.t7 VDPWR 0.016667f
C629 a_19190_31610.n5 VDPWR 0.034125f
C630 a_19190_31610.t4 VDPWR 0.025389f
C631 a_19190_31610.t6 VDPWR 0.02f
C632 a_19190_31610.t18 VDPWR 0.02f
C633 a_19190_31610.t17 VDPWR 0.032283f
C634 a_19190_31610.n6 VDPWR 0.036051f
C635 a_19190_31610.n7 VDPWR 0.024627f
C636 a_19190_31610.n8 VDPWR 0.039854f
C637 a_19190_31610.n9 VDPWR 0.176664f
C638 a_19190_31610.n10 VDPWR 0.242013f
C639 a_19190_31610.n11 VDPWR 0.017774f
C640 a_19190_31610.t1 VDPWR 0.031554f
C641 a_19190_31610.n12 VDPWR 0.019781f
C642 a_19190_31610.n13 VDPWR 0.511999f
C643 a_19190_31610.n14 VDPWR 0.172226f
C644 a_19190_31610.t12 VDPWR 0.025389f
C645 a_19190_31610.t14 VDPWR 0.02f
C646 a_19190_31610.t19 VDPWR 0.02f
C647 a_19190_31610.t20 VDPWR 0.032283f
C648 a_19190_31610.n15 VDPWR 0.036051f
C649 a_19190_31610.n16 VDPWR 0.024627f
C650 a_19190_31610.n17 VDPWR 0.039854f
C651 a_19190_31610.n18 VDPWR 0.221004f
C652 a_19190_31610.n19 VDPWR 0.034125f
C653 a_19190_31610.t15 VDPWR 0.016667f
C654 VGND.n7 VDPWR 0.010041f
C655 VGND.n11 VDPWR 0.010041f
C656 VGND.t304 VDPWR 0.067284f
C657 VGND.n22 VDPWR 0.029746f
C658 VGND.t149 VDPWR 0.030725f
C659 VGND.t126 VDPWR 0.052116f
C660 VGND.t20 VDPWR 0.052116f
C661 VGND.t330 VDPWR 0.034225f
C662 VGND.t315 VDPWR 0.034225f
C663 VGND.t66 VDPWR 0.017113f
C664 VGND.t192 VDPWR 0.056783f
C665 VGND.t40 VDPWR 0.058728f
C666 VGND.t135 VDPWR 0.024502f
C667 VGND.n47 VDPWR 0.010041f
C668 VGND.n54 VDPWR 0.011523f
C669 VGND.n56 VDPWR 0.010586f
C670 VGND.n62 VDPWR 0.010586f
C671 VGND.n70 VDPWR 0.010041f
C672 VGND.n77 VDPWR 0.010041f
C673 VGND.n97 VDPWR 0.010041f
C674 VGND.n100 VDPWR 0.011523f
C675 VGND.t87 VDPWR 0.028003f
C676 VGND.t104 VDPWR 0.028003f
C677 VGND.t168 VDPWR 0.046671f
C678 VGND.t13 VDPWR 0.048616f
C679 VGND.n106 VDPWR 0.023523f
C680 VGND.t102 VDPWR 0.024502f
C681 VGND.t68 VDPWR 0.028003f
C682 VGND.t0 VDPWR 0.028003f
C683 VGND.t30 VDPWR 0.046671f
C684 VGND.t128 VDPWR 0.048616f
C685 VGND.t82 VDPWR 0.024502f
C686 VGND.n117 VDPWR 0.010041f
C687 VGND.n125 VDPWR 0.011523f
C688 VGND.n140 VDPWR 0.104803f
C689 VGND.t317 VDPWR 0.351034f
C690 VGND.n142 VDPWR 0.234023f
C691 VGND.t17 VDPWR 0.010479f
C692 VGND.n148 VDPWR 0.025216f
C693 VGND.t318 VDPWR 0.015633f
C694 VGND.n150 VDPWR 0.016298f
C695 VGND.n151 VDPWR 0.016298f
C696 VGND.n154 VDPWR 0.029117f
C697 VGND.n155 VDPWR 0.078798f
C698 VGND.t311 VDPWR 0.181444f
C699 VGND.t16 VDPWR 0.143014f
C700 VGND.n156 VDPWR 0.20152f
C701 VGND.t6 VDPWR 0.010479f
C702 VGND.t158 VDPWR 0.028003f
C703 VGND.t166 VDPWR 0.028003f
C704 VGND.t80 VDPWR 0.043311f
C705 VGND.t7 VDPWR 0.203769f
C706 VGND.t119 VDPWR 0.181444f
C707 VGND.t8 VDPWR 0.010479f
C708 VGND.n160 VDPWR 0.077311f
C709 VGND.t120 VDPWR 0.015625f
C710 VGND.n162 VDPWR 0.01401f
C711 VGND.n164 VDPWR 0.010371f
C712 VGND.n165 VDPWR 0.010371f
C713 VGND.n167 VDPWR 0.019958f
C714 VGND.n169 VDPWR 0.20152f
C715 VGND.t5 VDPWR 0.143014f
C716 VGND.t313 VDPWR 0.181444f
C717 VGND.n170 VDPWR 0.077311f
C718 VGND.n172 VDPWR 0.019958f
C719 VGND.t314 VDPWR 0.015625f
C720 VGND.n174 VDPWR 0.010371f
C721 VGND.n175 VDPWR 0.010371f
C722 VGND.n178 VDPWR 0.01401f
C723 VGND.n188 VDPWR 0.107498f
C724 VGND.n189 VDPWR 0.079284f
C725 VGND.n191 VDPWR 0.012547f
C726 VGND.n197 VDPWR 0.010041f
C727 VGND.n205 VDPWR 0.023523f
C728 VGND.t36 VDPWR 0.048616f
C729 VGND.t97 VDPWR 0.046671f
C730 VGND.t309 VDPWR 0.028003f
C731 VGND.t42 VDPWR 0.028003f
C732 VGND.t44 VDPWR 0.024502f
C733 VGND.n206 VDPWR 0.023523f
C734 VGND.n237 VDPWR 0.011523f
C735 VGND.n243 VDPWR 0.010041f
C736 VGND.n251 VDPWR 0.023523f
C737 VGND.t156 VDPWR 0.050172f
C738 VGND.t323 VDPWR 0.048227f
C739 VGND.t46 VDPWR 0.034225f
C740 VGND.t93 VDPWR 0.034225f
C741 VGND.t174 VDPWR 0.045116f
C742 VGND.t133 VDPWR 0.045116f
C743 VGND.t300 VDPWR 0.028003f
C744 VGND.t188 VDPWR 0.028003f
C745 VGND.t34 VDPWR 0.035003f
C746 VGND.t106 VDPWR 0.035003f
C747 VGND.t115 VDPWR 0.030725f
C748 VGND.n252 VDPWR 0.029746f
C749 VGND.n265 VDPWR 0.012059f
C750 VGND.n291 VDPWR 0.071032f
C751 VGND.n305 VDPWR 0.010371f
C752 VGND.n307 VDPWR 0.010371f
C753 VGND.n308 VDPWR 0.01443f
C754 VGND.t63 VDPWR 0.015625f
C755 VGND.n310 VDPWR 0.014954f
C756 VGND.n314 VDPWR 0.010371f
C757 VGND.n315 VDPWR 0.014954f
C758 VGND.n317 VDPWR 0.010371f
C759 VGND.t121 VDPWR 0.015625f
C760 VGND.n319 VDPWR 0.01443f
C761 VGND.n321 VDPWR 0.135495f
C762 VGND.t62 VDPWR 0.112529f
C763 VGND.t308 VDPWR 0.238838f
C764 VGND.t2 VDPWR 0.238838f
C765 VGND.t95 VDPWR 0.112529f
C766 VGND.n326 VDPWR 0.019506f
C767 VGND.t191 VDPWR 0.015633f
C768 VGND.n329 VDPWR 0.016298f
C769 VGND.n330 VDPWR 0.016298f
C770 VGND.n332 VDPWR 0.016247f
C771 VGND.t59 VDPWR 0.015633f
C772 VGND.n336 VDPWR 0.016298f
C773 VGND.n337 VDPWR 0.016298f
C774 VGND.n339 VDPWR 0.019506f
C775 VGND.n369 VDPWR 0.013335f
C776 VGND.n380 VDPWR 0.010371f
C777 VGND.n383 VDPWR 0.010371f
C778 VGND.n384 VDPWR 0.01443f
C779 VGND.t322 VDPWR 0.015625f
C780 VGND.n386 VDPWR 0.014646f
C781 VGND.n387 VDPWR 0.010371f
C782 VGND.n390 VDPWR 0.010371f
C783 VGND.n391 VDPWR 0.01443f
C784 VGND.t65 VDPWR 0.015625f
C785 VGND.n393 VDPWR 0.014646f
C786 VGND.n396 VDPWR 0.010371f
C787 VGND.n399 VDPWR 0.010371f
C788 VGND.n400 VDPWR 0.01443f
C789 VGND.t25 VDPWR 0.015625f
C790 VGND.n402 VDPWR 0.014646f
C791 VGND.n403 VDPWR 0.010371f
C792 VGND.n406 VDPWR 0.010371f
C793 VGND.n407 VDPWR 0.01443f
C794 VGND.t329 VDPWR 0.015625f
C795 VGND.n409 VDPWR 0.014646f
C796 VGND.t53 VDPWR 0.022954f
C797 VGND.n410 VDPWR 0.024755f
C798 VGND.n428 VDPWR 0.010371f
C799 VGND.n431 VDPWR 0.010371f
C800 VGND.n432 VDPWR 0.01443f
C801 VGND.t146 VDPWR 0.015625f
C802 VGND.n434 VDPWR 0.014954f
C803 VGND.n435 VDPWR 0.010371f
C804 VGND.n438 VDPWR 0.010371f
C805 VGND.n439 VDPWR 0.01443f
C806 VGND.t327 VDPWR 0.015625f
C807 VGND.n441 VDPWR 0.014954f
C808 VGND.n447 VDPWR 0.010371f
C809 VGND.n450 VDPWR 0.010371f
C810 VGND.n451 VDPWR 0.01443f
C811 VGND.t307 VDPWR 0.015548f
C812 VGND.n453 VDPWR 0.014678f
C813 VGND.n455 VDPWR 0.010371f
C814 VGND.n458 VDPWR 0.010371f
C815 VGND.n459 VDPWR 0.01443f
C816 VGND.t123 VDPWR 0.015625f
C817 VGND.n461 VDPWR 0.014954f
C818 VGND.n483 VDPWR 0.013335f
C819 VGND.n486 VDPWR 0.013335f
C820 VGND.n487 VDPWR 0.017594f
C821 VGND.t303 VDPWR 0.020832f
C822 VGND.n489 VDPWR 0.017895f
C823 VGND.n490 VDPWR 0.013335f
C824 VGND.n493 VDPWR 0.013335f
C825 VGND.n494 VDPWR 0.017594f
C826 VGND.t71 VDPWR 0.020832f
C827 VGND.n496 VDPWR 0.017895f
C828 VGND.n503 VDPWR 0.013335f
C829 VGND.n506 VDPWR 0.013335f
C830 VGND.n507 VDPWR 0.017594f
C831 VGND.t84 VDPWR 0.020832f
C832 VGND.n509 VDPWR 0.017895f
C833 VGND.n513 VDPWR 0.057055f
C834 VGND.n517 VDPWR 0.013335f
C835 VGND.n520 VDPWR 0.013335f
C836 VGND.n521 VDPWR 0.017594f
C837 VGND.t316 VDPWR 0.020832f
C838 VGND.n523 VDPWR 0.017895f
C839 VGND.n524 VDPWR 0.013335f
C840 VGND.n527 VDPWR 0.013335f
C841 VGND.n528 VDPWR 0.017594f
C842 VGND.t112 VDPWR 0.020832f
C843 VGND.n530 VDPWR 0.017895f
C844 VGND.t334 VDPWR 0.33257f
C845 VGND.t336 VDPWR 0.350056f
C846 VGND.n541 VDPWR 0.643773f
C847 VGND.t335 VDPWR 0.350056f
C848 VGND.n542 VDPWR 0.339817f
C849 VGND.t340 VDPWR 0.328516f
C850 VGND.n543 VDPWR 0.403278f
C851 VGND.t210 VDPWR 0.165646f
C852 VGND.t217 VDPWR 0.174535f
C853 VGND.t213 VDPWR 0.174535f
C854 VGND.t218 VDPWR 0.174535f
C855 VGND.t219 VDPWR 0.174535f
C856 VGND.t247 VDPWR 0.174535f
C857 VGND.t220 VDPWR 0.174535f
C858 VGND.t256 VDPWR 0.174535f
C859 VGND.t216 VDPWR 0.166246f
C860 VGND.t259 VDPWR 0.080082f
C861 VGND.n544 VDPWR 0.103294f
C862 VGND.t244 VDPWR 0.181576f
C863 VGND.t214 VDPWR 0.166944f
C864 VGND.t243 VDPWR 0.174535f
C865 VGND.t239 VDPWR 0.174535f
C866 VGND.t242 VDPWR 0.174535f
C867 VGND.t238 VDPWR 0.174535f
C868 VGND.t229 VDPWR 0.174535f
C869 VGND.t246 VDPWR 0.174535f
C870 VGND.t215 VDPWR 0.174535f
C871 VGND.t245 VDPWR 0.269587f
C872 VGND.n545 VDPWR 0.410227f
C873 VGND.n547 VDPWR 0.079217f
C874 VGND.n548 VDPWR 0.011522f
C875 VGND.t273 VDPWR 0.010307f
C876 VGND.n549 VDPWR 0.011434f
C877 VGND.n551 VDPWR 0.079217f
C878 VGND.n552 VDPWR 0.011522f
C879 VGND.t276 VDPWR 0.010307f
C880 VGND.n553 VDPWR 0.011522f
C881 VGND.t279 VDPWR 0.010307f
C882 VGND.n555 VDPWR 0.079217f
C883 VGND.n557 VDPWR 0.079217f
C884 VGND.n559 VDPWR 0.079217f
C885 VGND.n561 VDPWR 0.079217f
C886 VGND.n563 VDPWR 0.079217f
C887 VGND.n565 VDPWR 0.079217f
C888 VGND.n567 VDPWR 0.079217f
C889 VGND.n569 VDPWR 0.107944f
C890 VGND.n570 VDPWR 0.034643f
C891 VGND.n572 VDPWR 0.011434f
C892 VGND.n573 VDPWR 0.036527f
C893 VGND.t278 VDPWR 0.030752f
C894 VGND.t143 VDPWR 0.024891f
C895 VGND.t3 VDPWR 0.024891f
C896 VGND.t54 VDPWR 0.024891f
C897 VGND.t151 VDPWR 0.024891f
C898 VGND.t180 VDPWR 0.024891f
C899 VGND.t176 VDPWR 0.024891f
C900 VGND.t160 VDPWR 0.024891f
C901 VGND.t11 VDPWR 0.024891f
C902 VGND.t109 VDPWR 0.024891f
C903 VGND.t74 VDPWR 0.024891f
C904 VGND.t178 VDPWR 0.024891f
C905 VGND.t325 VDPWR 0.024891f
C906 VGND.t48 VDPWR 0.024891f
C907 VGND.t164 VDPWR 0.024891f
C908 VGND.t85 VDPWR 0.024891f
C909 VGND.t72 VDPWR 0.024891f
C910 VGND.t124 VDPWR 0.024891f
C911 VGND.t78 VDPWR 0.024891f
C912 VGND.t275 VDPWR 0.037822f
C913 VGND.n574 VDPWR 0.031531f
C914 VGND.n575 VDPWR 0.011434f
C915 VGND.n577 VDPWR 0.024465f
C916 VGND.n578 VDPWR 0.08053f
C917 VGND.n580 VDPWR 0.079217f
C918 VGND.n582 VDPWR 0.079217f
C919 VGND.n584 VDPWR 0.079217f
C920 VGND.n586 VDPWR 0.079217f
C921 VGND.n588 VDPWR 0.079217f
C922 VGND.n590 VDPWR 0.079217f
C923 VGND.n592 VDPWR 0.079217f
C924 VGND.n594 VDPWR 0.079217f
C925 VGND.n595 VDPWR 0.08053f
C926 VGND.n596 VDPWR 0.032623f
C927 VGND.t297 VDPWR 0.010307f
C928 VGND.n598 VDPWR 0.011522f
C929 VGND.n599 VDPWR 0.038349f
C930 VGND.t296 VDPWR 0.031005f
C931 VGND.t198 VDPWR 0.024891f
C932 VGND.t137 VDPWR 0.024891f
C933 VGND.t91 VDPWR 0.024891f
C934 VGND.t117 VDPWR 0.024891f
C935 VGND.t22 VDPWR 0.024891f
C936 VGND.t204 VDPWR 0.024891f
C937 VGND.t206 VDPWR 0.024891f
C938 VGND.t89 VDPWR 0.024891f
C939 VGND.t162 VDPWR 0.024891f
C940 VGND.t153 VDPWR 0.024891f
C941 VGND.t28 VDPWR 0.024891f
C942 VGND.t208 VDPWR 0.024891f
C943 VGND.t200 VDPWR 0.024891f
C944 VGND.t50 VDPWR 0.024891f
C945 VGND.t76 VDPWR 0.024891f
C946 VGND.t99 VDPWR 0.024891f
C947 VGND.t319 VDPWR 0.024891f
C948 VGND.t202 VDPWR 0.024891f
C949 VGND.t272 VDPWR 0.037246f
C950 VGND.n600 VDPWR 0.030033f
C951 VGND.n601 VDPWR 0.011434f
C952 VGND.n603 VDPWR 0.018358f
C953 VGND.n604 VDPWR 0.221781f
C954 VGND.n605 VDPWR 0.159089f
C955 VGND.n606 VDPWR 0.034589f
C956 VGND.n607 VDPWR 0.118908f
C957 VGND.t268 VDPWR 0.04239f
C958 VGND.n611 VDPWR 0.010371f
C959 VGND.n618 VDPWR 0.010371f
C960 VGND.n619 VDPWR 0.034589f
C961 VGND.n620 VDPWR 0.118908f
C962 VGND.n621 VDPWR 0.034589f
C963 VGND.n622 VDPWR 0.118908f
C964 VGND.n623 VDPWR 0.034589f
C965 VGND.n624 VDPWR 0.118908f
C966 VGND.n625 VDPWR 0.034589f
C967 VGND.n626 VDPWR 0.118908f
C968 VGND.n627 VDPWR 0.034589f
C969 VGND.n628 VDPWR 0.118908f
C970 VGND.n629 VDPWR 0.034589f
C971 VGND.n630 VDPWR 0.118908f
C972 VGND.n631 VDPWR 0.034589f
C973 VGND.n632 VDPWR 0.169411f
C974 VGND.t283 VDPWR 0.04239f
C975 VGND.n633 VDPWR 0.01712f
C976 VGND.n634 VDPWR 0.013168f
C977 VGND.n639 VDPWR 0.010371f
C978 VGND.n641 VDPWR 0.010309f
C979 VGND.n642 VDPWR 0.010309f
C980 VGND.n644 VDPWR 0.010371f
C981 VGND.n645 VDPWR 0.010371f
C982 VGND.n647 VDPWR 0.012504f
C983 VGND.n649 VDPWR 0.083119f
C984 VGND.t284 VDPWR 0.088157f
C985 VGND.t248 VDPWR 0.090675f
C986 VGND.t240 VDPWR 0.090675f
C987 VGND.t260 VDPWR 0.090675f
C988 VGND.t257 VDPWR 0.090675f
C989 VGND.t254 VDPWR 0.090675f
C990 VGND.t252 VDPWR 0.090675f
C991 VGND.t250 VDPWR 0.090675f
C992 VGND.t227 VDPWR 0.090675f
C993 VGND.t234 VDPWR 0.090675f
C994 VGND.t232 VDPWR 0.090675f
C995 VGND.t221 VDPWR 0.090675f
C996 VGND.t230 VDPWR 0.090675f
C997 VGND.t236 VDPWR 0.090675f
C998 VGND.t225 VDPWR 0.090675f
C999 VGND.t223 VDPWR 0.090675f
C1000 VGND.t211 VDPWR 0.090675f
C1001 VGND.t269 VDPWR 0.088157f
C1002 VGND.n653 VDPWR 0.010309f
C1003 VGND.n654 VDPWR 0.010309f
C1004 VGND.n655 VDPWR 0.010371f
C1005 VGND.n656 VDPWR 0.010371f
C1006 VGND.n658 VDPWR 0.012504f
C1007 VGND.n660 VDPWR 0.083119f
C1008 VGND.n664 VDPWR 0.010371f
C1009 VGND.n666 VDPWR 0.013168f
C1010 VGND.n667 VDPWR 0.016248f
C1011 VGND.n668 VDPWR 0.100269f
C1012 VGND.n669 VDPWR 0.098876f
C1013 VGND.n670 VDPWR 0.011522f
C1014 VGND.t267 VDPWR 0.010307f
C1015 VGND.n671 VDPWR 0.012116f
C1016 VGND.n672 VDPWR 0.03773f
C1017 VGND.t294 VDPWR 0.011758f
C1018 VGND.n674 VDPWR 0.012203f
C1019 VGND.n675 VDPWR 0.037099f
C1020 VGND.t293 VDPWR 0.03018f
C1021 VGND.t101 VDPWR 0.022817f
C1022 VGND.t155 VDPWR 0.022817f
C1023 VGND.t266 VDPWR 0.035815f
C1024 VGND.n676 VDPWR 0.02939f
C1025 VGND.n677 VDPWR 0.011434f
C1026 VGND.n679 VDPWR 0.020303f
C1027 VGND.n680 VDPWR 0.244582f
C1028 VGND.n681 VDPWR 0.091811f
C1029 VGND.n683 VDPWR 0.035085f
C1030 VGND.n684 VDPWR 0.01161f
C1031 VGND.n685 VDPWR 0.011434f
C1032 VGND.t264 VDPWR 0.010307f
C1033 VGND.n688 VDPWR 0.035085f
C1034 VGND.n689 VDPWR 0.01161f
C1035 VGND.n690 VDPWR 0.011434f
C1036 VGND.t288 VDPWR 0.010307f
C1037 VGND.n693 VDPWR 0.035085f
C1038 VGND.n695 VDPWR 0.035085f
C1039 VGND.n697 VDPWR 0.035085f
C1040 VGND.n699 VDPWR 0.043343f
C1041 VGND.n700 VDPWR 0.014694f
C1042 VGND.n701 VDPWR 0.019513f
C1043 VGND.n702 VDPWR 0.01161f
C1044 VGND.n703 VDPWR 0.035951f
C1045 VGND.t287 VDPWR 0.029254f
C1046 VGND.t298 VDPWR 0.022817f
C1047 VGND.t139 VDPWR 0.022817f
C1048 VGND.t147 VDPWR 0.022817f
C1049 VGND.t32 VDPWR 0.022817f
C1050 VGND.t38 VDPWR 0.022817f
C1051 VGND.t26 VDPWR 0.022817f
C1052 VGND.t141 VDPWR 0.022817f
C1053 VGND.t184 VDPWR 0.022817f
C1054 VGND.t170 VDPWR 0.022817f
C1055 VGND.t332 VDPWR 0.022817f
C1056 VGND.t290 VDPWR 0.035815f
C1057 VGND.n704 VDPWR 0.02939f
C1058 VGND.t291 VDPWR 0.010307f
C1059 VGND.n705 VDPWR 0.011434f
C1060 VGND.n706 VDPWR 0.019513f
C1061 VGND.n707 VDPWR 0.014063f
C1062 VGND.n708 VDPWR 0.023706f
C1063 VGND.n710 VDPWR 0.035085f
C1064 VGND.n712 VDPWR 0.035085f
C1065 VGND.n714 VDPWR 0.035085f
C1066 VGND.n716 VDPWR 0.035085f
C1067 VGND.n717 VDPWR 0.023706f
C1068 VGND.n718 VDPWR 0.014063f
C1069 VGND.n719 VDPWR 0.019513f
C1070 VGND.n720 VDPWR 0.01161f
C1071 VGND.n721 VDPWR 0.035951f
C1072 VGND.t263 VDPWR 0.029254f
C1073 VGND.t113 VDPWR 0.022817f
C1074 VGND.t9 VDPWR 0.022817f
C1075 VGND.t18 VDPWR 0.022817f
C1076 VGND.t172 VDPWR 0.022817f
C1077 VGND.t131 VDPWR 0.022817f
C1078 VGND.t56 VDPWR 0.022817f
C1079 VGND.t186 VDPWR 0.022817f
C1080 VGND.t196 VDPWR 0.022817f
C1081 VGND.t194 VDPWR 0.022817f
C1082 VGND.t60 VDPWR 0.022817f
C1083 VGND.t281 VDPWR 0.035815f
C1084 VGND.n722 VDPWR 0.02939f
C1085 VGND.t282 VDPWR 0.010307f
C1086 VGND.n723 VDPWR 0.011434f
C1087 VGND.n724 VDPWR 0.019513f
C1088 VGND.n725 VDPWR 0.014063f
C1089 VGND.n726 VDPWR 0.112477f
C1090 VGND.n727 VDPWR 0.139739f
C1091 VGND.n728 VDPWR 0.054347f
C1092 VGND.n730 VDPWR 0.017895f
C1093 VGND.n732 VDPWR 0.013335f
C1094 VGND.t183 VDPWR 0.020832f
C1095 VGND.n734 VDPWR 0.017594f
C1096 VGND.t182 VDPWR 0.218169f
C1097 VGND.n736 VDPWR 0.179129f
C1098 VGND.t108 VDPWR 0.236542f
C1099 VGND.t111 VDPWR 0.208983f
C1100 VGND.n737 VDPWR 0.179129f
C1101 VGND.t15 VDPWR 0.179129f
C1102 VGND.n738 VDPWR 0.179129f
C1103 VGND.t70 VDPWR 0.179129f
C1104 VGND.n739 VDPWR 0.195204f
C1105 VGND.n740 VDPWR 0.126309f
C1106 VGND.t321 VDPWR 0.062006f
C1107 VGND.t64 VDPWR 0.062006f
C1108 VGND.n741 VDPWR 0.089564f
C1109 VGND.n742 VDPWR 0.089564f
C1110 VGND.t24 VDPWR 0.062006f
C1111 VGND.t328 VDPWR 0.062006f
C1112 VGND.n743 VDPWR 0.089564f
C1113 VGND.n744 VDPWR 0.089564f
C1114 VGND.t52 VDPWR 0.057413f
C1115 VGND.t306 VDPWR 0.055117f
C1116 VGND.t122 VDPWR 0.062006f
C1117 VGND.n745 VDPWR 0.121716f
C1118 VGND.n746 VDPWR 0.126309f
C1119 VGND.t145 VDPWR 0.112529f
C1120 VGND.t190 VDPWR 0.238838f
C1121 VGND.t130 VDPWR 0.238838f
C1122 VGND.t58 VDPWR 0.112529f
C1123 VGND.n747 VDPWR 0.124012f
C1124 VGND.n749 VDPWR 0.016247f
C1125 VGND.n761 VDPWR 0.047025f
C1126 VGND.n762 VDPWR 2.38943f
C1127 VGND.n763 VDPWR 0.029632f
C1128 VGND.n764 VDPWR 2.5638f
C1129 VGND.n765 VDPWR 0.029632f
C1130 VGND.n767 VDPWR 0.029632f
C1131 VGND.n769 VDPWR 0.029632f
C1132 VGND.n770 VDPWR 0.029632f
C1133 VGND.n771 VDPWR 4.91738f
C1134 VGND.n772 VDPWR 5.08938f
C1135 a_14348_27710.t37 VDPWR 0.176337f
C1136 a_14348_27710.n0 VDPWR 0.064494f
C1137 a_14348_27710.t38 VDPWR 0.1754f
C1138 a_14348_27710.n1 VDPWR 0.073075f
C1139 a_14348_27710.t27 VDPWR 0.177279f
C1140 a_14348_27710.t28 VDPWR 0.176515f
C1141 a_14348_27710.n2 VDPWR 0.219612f
C1142 a_14348_27710.t15 VDPWR 0.176515f
C1143 a_14348_27710.n3 VDPWR 0.121656f
C1144 a_14348_27710.t16 VDPWR 0.176515f
C1145 a_14348_27710.n4 VDPWR 0.121656f
C1146 a_14348_27710.t18 VDPWR 0.176515f
C1147 a_14348_27710.n5 VDPWR 0.121656f
C1148 a_14348_27710.t19 VDPWR 0.176515f
C1149 a_14348_27710.n6 VDPWR 0.121656f
C1150 a_14348_27710.t20 VDPWR 0.176515f
C1151 a_14348_27710.n7 VDPWR 0.121656f
C1152 a_14348_27710.t42 VDPWR 0.177201f
C1153 a_14348_27710.n8 VDPWR 0.113324f
C1154 a_14348_27710.n9 VDPWR 0.034404f
C1155 a_14348_27710.t48 VDPWR 0.177779f
C1156 a_14348_27710.t47 VDPWR 0.176515f
C1157 a_14348_27710.n10 VDPWR 0.220068f
C1158 a_14348_27710.t46 VDPWR 0.176515f
C1159 a_14348_27710.n11 VDPWR 0.121656f
C1160 a_14348_27710.t33 VDPWR 0.176515f
C1161 a_14348_27710.n12 VDPWR 0.121656f
C1162 a_14348_27710.t40 VDPWR 0.176515f
C1163 a_14348_27710.n13 VDPWR 0.121656f
C1164 a_14348_27710.t39 VDPWR 0.176515f
C1165 a_14348_27710.n14 VDPWR 0.121656f
C1166 a_14348_27710.n15 VDPWR 0.034404f
C1167 a_14348_27710.n16 VDPWR 0.022936f
C1168 a_14348_27710.n17 VDPWR 0.127424f
C1169 a_14348_27710.t7 VDPWR 0.174413f
C1170 a_14348_27710.n18 VDPWR 0.48222f
C1171 a_14348_27710.t2 VDPWR 0.012742f
C1172 a_14348_27710.t11 VDPWR 0.012742f
C1173 a_14348_27710.n19 VDPWR 0.027525f
C1174 a_14348_27710.n20 VDPWR 0.259414f
C1175 a_14348_27710.t8 VDPWR 0.012742f
C1176 a_14348_27710.t9 VDPWR 0.012742f
C1177 a_14348_27710.n21 VDPWR 0.027525f
C1178 a_14348_27710.n22 VDPWR 0.278292f
C1179 a_14348_27710.t10 VDPWR 0.012742f
C1180 a_14348_27710.t12 VDPWR 0.012742f
C1181 a_14348_27710.n23 VDPWR 0.027525f
C1182 a_14348_27710.n24 VDPWR 0.270646f
C1183 a_14348_27710.t6 VDPWR 0.012742f
C1184 a_14348_27710.t0 VDPWR 0.012742f
C1185 a_14348_27710.n25 VDPWR 0.02609f
C1186 a_14348_27710.t4 VDPWR 0.012742f
C1187 a_14348_27710.t3 VDPWR 0.012742f
C1188 a_14348_27710.n26 VDPWR 0.029654f
C1189 a_14348_27710.n27 VDPWR 0.349463f
C1190 a_14348_27710.t13 VDPWR 0.012742f
C1191 a_14348_27710.t1 VDPWR 0.012742f
C1192 a_14348_27710.n28 VDPWR 0.02609f
C1193 a_14348_27710.n29 VDPWR 0.216014f
C1194 a_14348_27710.n30 VDPWR 0.654381f
C1195 a_14348_27710.t14 VDPWR 0.509694f
C1196 a_14348_27710.t23 VDPWR 0.518153f
C1197 a_14348_27710.t43 VDPWR 0.509694f
C1198 a_14348_27710.n31 VDPWR 0.338771f
C1199 a_14348_27710.t22 VDPWR 0.509694f
C1200 a_14348_27710.n32 VDPWR 0.222991f
C1201 a_14348_27710.t41 VDPWR 0.509694f
C1202 a_14348_27710.n33 VDPWR 0.222991f
C1203 a_14348_27710.t32 VDPWR 0.509694f
C1204 a_14348_27710.n34 VDPWR 0.222991f
C1205 a_14348_27710.t26 VDPWR 0.509694f
C1206 a_14348_27710.n35 VDPWR 0.222991f
C1207 a_14348_27710.t31 VDPWR 0.509694f
C1208 a_14348_27710.n36 VDPWR 0.222991f
C1209 a_14348_27710.t25 VDPWR 0.509694f
C1210 a_14348_27710.n37 VDPWR 0.222991f
C1211 a_14348_27710.t44 VDPWR 0.509694f
C1212 a_14348_27710.n38 VDPWR 0.215027f
C1213 a_14348_27710.t24 VDPWR 0.509694f
C1214 a_14348_27710.n39 VDPWR 0.230955f
C1215 a_14348_27710.n40 VDPWR 0.230955f
C1216 a_14348_27710.t36 VDPWR 0.509694f
C1217 a_14348_27710.n41 VDPWR 0.215027f
C1218 a_14348_27710.t17 VDPWR 0.509694f
C1219 a_14348_27710.n42 VDPWR 0.222991f
C1220 a_14348_27710.t29 VDPWR 0.509694f
C1221 a_14348_27710.n43 VDPWR 0.222991f
C1222 a_14348_27710.t21 VDPWR 0.509694f
C1223 a_14348_27710.n44 VDPWR 0.222991f
C1224 a_14348_27710.t30 VDPWR 0.509694f
C1225 a_14348_27710.n45 VDPWR 0.222991f
C1226 a_14348_27710.t34 VDPWR 0.509694f
C1227 a_14348_27710.n46 VDPWR 0.222991f
C1228 a_14348_27710.t45 VDPWR 0.509694f
C1229 a_14348_27710.n47 VDPWR 0.222991f
C1230 a_14348_27710.t35 VDPWR 0.509694f
C1231 a_14348_27710.n48 VDPWR 0.221398f
C1232 a_14348_27710.t49 VDPWR 0.509694f
C1233 a_14348_27710.n49 VDPWR 0.391094f
C1234 a_14348_27710.n50 VDPWR 1.23441f
C1235 a_14348_27710.t5 VDPWR 0.111663f
C1236 a_19190_29050.n0 VDPWR 1.02458f
C1237 a_19190_29050.n1 VDPWR 1.10014f
C1238 a_19190_29050.n2 VDPWR 1.33269f
C1239 a_19190_29050.n3 VDPWR 0.153679f
C1240 a_19190_29050.n4 VDPWR 3.88852f
C1241 a_19190_29050.t36 VDPWR 0.021247f
C1242 a_19190_29050.n5 VDPWR 0.019024f
C1243 a_19190_29050.t17 VDPWR 0.013904f
C1244 a_19190_29050.t13 VDPWR 0.013904f
C1245 a_19190_29050.n6 VDPWR 0.026482f
C1246 a_19190_29050.n7 VDPWR 0.019024f
C1247 a_19190_29050.t8 VDPWR 0.015816f
C1248 a_19190_29050.n8 VDPWR 0.011348f
C1249 a_19190_29050.n9 VDPWR 0.010949f
C1250 a_19190_29050.n10 VDPWR 0.292028f
C1251 a_19190_29050.t11 VDPWR 0.013904f
C1252 a_19190_29050.t34 VDPWR 0.013904f
C1253 a_19190_29050.n11 VDPWR 0.025867f
C1254 a_19190_29050.t25 VDPWR 0.359229f
C1255 a_19190_29050.t18 VDPWR 0.36519f
C1256 a_19190_29050.t35 VDPWR 0.359229f
C1257 a_19190_29050.t15 VDPWR 0.359229f
C1258 a_19190_29050.t33 VDPWR 0.359229f
C1259 a_19190_29050.t29 VDPWR 0.359229f
C1260 a_19190_29050.t22 VDPWR 0.359229f
C1261 a_19190_29050.t27 VDPWR 0.359229f
C1262 a_19190_29050.t21 VDPWR 0.359229f
C1263 a_19190_29050.t12 VDPWR 0.359229f
C1264 a_19190_29050.t19 VDPWR 0.359229f
C1265 a_19190_29050.t20 VDPWR 0.359229f
C1266 a_19190_29050.t26 VDPWR 0.359229f
C1267 a_19190_29050.t31 VDPWR 0.359229f
C1268 a_19190_29050.t28 VDPWR 0.359229f
C1269 a_19190_29050.t32 VDPWR 0.359229f
C1270 a_19190_29050.t14 VDPWR 0.359229f
C1271 a_19190_29050.t23 VDPWR 0.359229f
C1272 a_19190_29050.t16 VDPWR 0.359229f
C1273 a_19190_29050.t24 VDPWR 0.359229f
C1274 a_19190_29050.t30 VDPWR 0.021589f
C1275 a_19190_29050.n12 VDPWR 0.019024f
.ends

