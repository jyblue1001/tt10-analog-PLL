* PEX produced on Tue Sep  2 04:44:30 AM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from project_5.ext - technology: sky130A

.subckt project_5 ua[0] VDPWR VGND
X0 VGND.t300 V_CONT.t5 sky130_fd_pr__cap_mim_m3_1 l=60 w=13.8
X1 a_14930_6670.t1 a_11860_6640.t3 VGND.t124 VGND.t123 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X2 VDPWR.t106 a_17714_9374.t9 a_18160_10940.t6 VDPWR.t105 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X3 a_19550_2800.t0 a_18930_3150.t3 a_19250_3100.t0 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X4 a_11200_9430.t14 VDPWR.t211 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5 a_12300_6670.t0 a_11780_7290.t3 a_11860_6640.t1 VDPWR.t379 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X6 a_12290_3150.t2 a_12070_2860.t3 a_12870_2890.t0 VGND.t85 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X7 a_19250_3100.t1 a_18330_3180.t2 VDPWR.t202 VDPWR.t201 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X8 VDPWR.t213 a_11200_9430.t15 a_9570_16200.t3 VDPWR.t212 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X9 VDPWR.t321 VDPWR.t319 a_9450_16252.t5 VDPWR.t320 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X10 VDPWR.t132 a_11200_9430.t16 a_10480_13480.t5 VDPWR.t131 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X11 a_9450_17070.t6 a_9450_16252.t2 VGND.t143 sky130_fd_pr__res_high_po_0p35 l=2.05
X12 a_11200_9430.t17 VDPWR.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X13 VDPWR.t189 a_13200_10990.t10 a_13200_10990.t11 VDPWR.t188 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X14 a_13070_11250.t10 a_10000_15820.t6 a_13360_11960.t4 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X15 a_20140_2930.t2 a_20230_3150.t3 VGND.t249 VGND.t248 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X16 VDPWR.t64 a_17950_3100.t2 a_17540_2930.t0 VDPWR.t63 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X17 a_16000_6670.t1 a_15320_6670.t2 a_12960_8860.t17 VDPWR.t200 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X18 VGND.t163 pll_bgr_magic_3_0.VV1.t5 a_15870_5490.t8 VGND.t162 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X19 a_12380_5460.t0 a_12760_5460.t3 a_12680_5910.t0 VDPWR.t175 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X20 VGND.t106 a_11040_2860.t2 a_10910_3020.t2 VGND.t105 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X21 VGND.t178 a_16240_3020.t4 a_15820_2860.t0 VGND.t177 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X22 a_17630_3150.t1 a_18330_3180.t3 VDPWR.t338 VDPWR.t337 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X23 VDPWR.t413 a_13200_10990.t17 a_13070_11250.t5 VDPWR.t412 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X24 a_13070_11250.t9 a_10000_15820.t7 a_13360_11960.t2 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X25 VGND.t72 a_12070_2860.t4 a_11960_2860.t2 VGND.t71 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X26 VGND.t253 a_12960_8860.t18 a_18390_5940.t5 VGND.t252 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X27 VGND.t60 VDPWR.t423 a_11200_9430.t10 VGND.t58 sky130_fd_pr__nfet_01v8 ad=1.01 pd=6.15 as=1 ps=5.8 w=2.5 l=5
X28 a_13070_11250.t11 a_15790_17280.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X29 VDPWR.t358 a_10160_10990.t17 a_10030_11260.t8 VDPWR.t357 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X30 a_10751_12090.t10 a_9450_16252.t10 VDPWR.t52 VDPWR.t51 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X31 a_18160_10940.t5 a_18160_10940.t3 a_18160_10940.t4 VDPWR.t83 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X32 a_20850_2800.t0 a_20230_3150.t4 a_20550_3100.t1 VGND.t34 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X33 a_18390_5940.t3 a_15870_5490.t10 VDPWR.t340 VDPWR.t339 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X34 VGND.t242 VGND.t240 VGND.t242 VGND.t241 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X35 a_20550_3100.t0 a_19630_3180.t2 VDPWR.t1 VDPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X36 a_9450_16252.t6 VDPWR.t424 VGND.t61 VGND.t58 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X37 a_13070_11250.t12 a_15790_17280.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 a_15320_5490.t0 a_14930_5490.t2 VDPWR.t191 VDPWR.t190 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X39 a_12380_6640.t0 a_12760_6640.t3 a_12680_6670.t0 VDPWR.t175 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X40 VDPWR.t404 a_10160_10990.t15 a_10160_10990.t16 VDPWR.t403 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X41 a_12540_2890.t2 a_12700_3340.t2 VGND.t158 VGND.t157 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X42 VGND.t239 VGND.t236 VGND.t238 VGND.t237 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X43 a_11200_9430.t18 VDPWR.t359 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X44 a_10060_12570.t9 a_9570_16200.t7 a_10160_10990.t4 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X45 VDPWR.t116 a_14010_6640.t2 a_13680_6640.t0 VDPWR.t115 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X46 a_10030_11260.t11 a_9450_17070.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X47 a_13200_5910.t0 a_12380_5460.t3 a_12760_5460.t0 VDPWR.t2 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X48 a_18510_9670.t7 V_CONT.t8 a_19530_10890.t5 VGND.t175 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X49 VDPWR.t128 a_10160_10990.t13 a_10160_10990.t14 VDPWR.t127 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X50 a_11200_9430.t19 VDPWR.t360 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X51 VGND.t193 VGND.t235 a_10900_14480.t8 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X52 VGND.t295 a_10120_15820.t1 VGND.t27 sky130_fd_pr__res_xhigh_po_0p35 l=6
X53 a_22240_2700.t1 a_21720_2700.t2 a_22130_3360.t0 VDPWR.t328 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X54 a_12960_8860.t16 VDPWR.t316 VDPWR.t318 VDPWR.t317 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X55 VGND.t234 VGND.t232 VGND.t234 VGND.t233 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X56 a_18160_10940.t10 a_18390_5940.t6 pll_bgr_magic_3_0.VV1.t4 VDPWR.t248 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X57 a_12960_8860.t10 a_9450_16252.t11 VDPWR.t54 VDPWR.t53 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X58 a_9570_16200.t2 a_11200_9430.t20 VDPWR.t348 VDPWR.t347 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X59 VDPWR.t402 a_13200_10990.t8 a_13200_10990.t9 VDPWR.t401 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X60 a_10030_11260.t12 a_9450_17070.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X61 VDPWR.t90 a_12070_2860.t5 a_11040_2860.t0 VDPWR.t89 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X62 a_15320_6670.t1 VGND.t301 a_14930_6670.t0 VDPWR.t190 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X63 VDPWR.t215 a_18930_3150.t4 a_18330_3180.t0 VDPWR.t214 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X64 ua1.t0 a_22240_2700.t2 a_22650_1940.t0 VGND.t46 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X65 a_18390_5940.t4 a_12960_8860.t19 VGND.t265 VGND.t264 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X66 VDPWR.t344 a_10030_11260.t13 a_9450_16252.t8 VDPWR.t343 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X67 VGND.t251 V_CONT.t9 a_22130_1940.t2 VGND.t159 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X68 a_10751_12090.t9 a_9450_16252.t12 VDPWR.t172 VDPWR.t171 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X69 VGND.t74 a_10751_12090.t0 VGND.t73 sky130_fd_pr__res_xhigh_po_0p35 l=1
X70 a_13070_11250.t13 a_15790_17280.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X71 a_13200_6670.t0 a_12380_6640.t3 a_12760_6640.t1 VDPWR.t2 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X72 a_10000_15820.t4 a_11200_9430.t21 VDPWR.t350 VDPWR.t349 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X73 VDPWR.t104 a_17714_9374.t2 a_17714_9374.t3 VDPWR.t103 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X74 VDPWR.t245 a_11040_2860.t3 a_10780_3220.t0 VDPWR.t244 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X75 VGND.t277 a_18840_2930.t4 a_18330_3180.t1 VGND.t276 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X76 a_14930_5490.t0 a_11860_5460.t3 VDPWR.t110 VDPWR.t109 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X77 VDPWR.t150 a_12700_3340.t3 a_12650_3210.t1 VDPWR.t149 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X78 VGND.t180 a_11860_5460.t4 a_11780_5490.t2 VGND.t179 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X79 VDPWR.t112 a_13200_10990.t18 a_13070_11250.t4 VDPWR.t111 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X80 VGND.t193 VGND.t230 a_10900_14480.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X81 a_18160_10940.t7 a_17714_9374.t10 VDPWR.t102 VDPWR.t101 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X82 VGND.t193 VGND.t231 a_10900_14480.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X83 a_11200_9430.t22 VDPWR.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X84 VGND.t174 a_18390_10330.t2 a_18390_10330.t3 VGND.t173 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X85 a_12960_8860.t9 a_9450_16252.t13 VDPWR.t174 VDPWR.t173 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X86 a_10030_11260.t14 a_9450_17070.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X87 VGND.t16 a_16000_6670.t3 V_CONT.t0 VGND.t15 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X88 VDPWR.t187 a_13070_11250.t14 a_11200_9430.t5 VDPWR.t186 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X89 a_13360_11960.t9 a_11840_9460.t8 a_13200_10990.t15 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X90 a_21690_4400.t0 V_CONT.t10 VGND.t170 VGND.t169 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X91 VDPWR.t179 a_10160_10990.t11 a_10160_10990.t12 VDPWR.t178 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X92 a_14160_5490.t0 a_13720_5910.t3 VDPWR.t25 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X93 a_13070_11250.t15 a_15790_17280.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X94 a_14930_6670.t2 a_11860_6640.t4 VDPWR.t336 VDPWR.t109 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X95 VGND.t229 VGND.t228 VGND.t229 VGND.t162 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X96 a_10030_11260.t15 a_9450_17070.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X97 VDPWR.t331 VGND.t302 a_21610_3360.t0 VDPWR.t330 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X98 VDPWR.t315 VDPWR.t313 VDPWR.t315 VDPWR.t314 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X99 VDPWR.t422 a_13070_11250.t16 a_11200_9430.t13 VDPWR.t421 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X100 a_10751_12090.t8 a_9450_16252.t14 VDPWR.t135 VDPWR.t134 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X101 a_16000_6670.t4 a_15710_6670.t0 sky130_fd_pr__cap_mim_m3_1 l=3.8 w=2.7
X102 a_18930_3150.t0 a_19630_3180.t3 VDPWR.t243 VDPWR.t242 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X103 a_13070_11250.t17 a_15790_17280.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X104 a_11860_5460.t1 a_11780_5490.t3 VGND.t32 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X105 VDPWR.t312 VDPWR.t310 VDPWR.t312 VDPWR.t311 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X106 a_15710_6670.t2 a_15320_6670.t3 VGND.t152 VGND.t151 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X107 a_10030_11260.t16 a_9450_17070.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X108 VGND.t50 a_12380_6640.t4 a_11860_6640.t0 VGND.t49 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X109 a_13280_3020.t2 a_12070_2860.t6 VGND.t101 VGND.t100 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X110 a_18390_10330.t5 V_CONT.t11 a_18160_10940.t11 VDPWR.t333 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X111 a_9450_16252.t9 a_10030_11260.t17 VDPWR.t346 VDPWR.t345 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X112 a_13070_11250.t18 a_15790_17280.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X113 a_18410_9620.t7 a_18410_9620.t6 VGND.t70 VGND.t69 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X114 a_10060_12570.t4 a_10751_12090.t13 a_10030_11260.t2 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X115 a_11200_9430.t23 VDPWR.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X116 VGND.t62 VDPWR.t425 a_10060_12570.t10 VGND.t58 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X117 VGND.t56 a_14340_6640.t2 a_14010_6640.t0 VGND.t55 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X118 a_11780_7290.t0 a_10780_3220.t2 VGND.t115 VGND.t114 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X119 VDPWR.t4 a_13200_10990.t6 a_13200_10990.t7 VDPWR.t3 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X120 a_13910_2890.t0 a_12070_2860.t7 a_13800_2890.t0 VGND.t102 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X121 a_16000_5490.t0 a_15320_5490.t2 a_15870_5490.t1 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X122 VDPWR.t181 a_10030_11260.t18 a_9450_16252.t1 VDPWR.t180 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X123 a_14890_17428.t1 a_14770_15820.t1 VGND.t168 sky130_fd_pr__res_xhigh_po_0p35 l=6
X124 a_11540_2890.t0 a_11040_2860.t4 a_11430_2890.t0 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X125 a_10000_17428.t0 a_10000_15820.t0 VGND.t27 sky130_fd_pr__res_xhigh_po_0p35 l=6
X126 a_15870_5490.t7 pll_bgr_magic_3_0.VV1.t6 VGND.t126 VGND.t125 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X127 a_11200_9430.t24 VDPWR.t207 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X128 a_18510_9670.t1 a_18410_9620.t9 VGND.t18 VGND.t17 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X129 VGND.t145 a_17030_3180.t2 a_18250_2800.t0 VGND.t144 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X130 a_10060_12570.t3 a_10751_12090.t14 a_10030_11260.t0 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X131 a_11200_9430.t25 VDPWR.t208 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X132 a_12960_8860.t8 a_9450_16252.t15 VDPWR.t137 VDPWR.t136 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X133 pll_bgr_magic_3_0.VV3.t1 a_18390_5940.t7 a_18510_9670.t3 VGND.t150 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X134 V_CONT.t7 a_16000_6670.t5 VGND.t286 VGND.t285 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X135 a_15050_2860.t3 a_15160_2860.t3 VGND.t292 VGND.t291 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X136 a_13720_5910.t0 a_11860_6640.t5 VDPWR.t335 VDPWR.t334 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.805 ps=5 w=2 l=0.15
X137 VDPWR.t13 a_10160_10990.t18 a_10030_11260.t7 VDPWR.t12 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X138 VGND.t188 VDPWR.t426 a_21610_1940.t0 VGND.t94 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X139 a_10030_11260.t19 a_9450_17070.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X140 a_18510_9670.t12 a_18510_9670.t11 a_18510_9670.t12 VGND.t91 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X141 ua1.t1 a_22240_2700.t3 a_22650_3360.t0 VDPWR.t238 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X142 VDPWR.t118 a_16000_5490.t3 V_CONT.t1 VDPWR.t117 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X143 a_16650_3100.t1 a_12070_2860.t8 VDPWR.t73 VDPWR.t72 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X144 a_10751_12090.t7 a_9450_16252.t16 VDPWR.t142 VDPWR.t141 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X145 VDPWR.t240 a_11200_9430.t26 a_10000_15820.t3 VDPWR.t239 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X146 VGND.t193 VGND.t227 a_11840_9460.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X147 VDPWR.t309 VDPWR.t306 VDPWR.t308 VDPWR.t307 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X148 a_9570_17278.t1 a_9570_16200.t6 VGND.t95 sky130_fd_pr__res_xhigh_po_0p35 l=3.35
X149 VGND.t193 VGND.t218 a_10900_14480.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X150 VGND.t128 a_12760_5460.t4 a_12380_5460.t1 VGND.t127 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X151 a_20230_3150.t0 ua1.t2 VGND.t42 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X152 VGND.t303 a_15288_18640.t1 sky130_fd_pr__cap_mim_m3_1 l=60 w=69.8
X153 a_13280_3020.t1 a_12070_2860.t9 VGND.t45 VGND.t44 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X154 VDPWR.t144 a_9450_16252.t17 a_12960_8860.t7 VDPWR.t143 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X155 a_13070_11250.t19 a_15790_17280.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X156 a_10060_12570.t2 a_10751_12090.t15 a_10030_11260.t9 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X157 VGND.t47 V_CONT.t12 a_22650_1940.t2 VGND.t46 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X158 a_15380_3150.t1 a_15160_2860.t4 a_15850_2890.t1 VGND.t120 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X159 VGND.t24 a_12070_2860.t10 a_16950_2890.t1 VGND.t23 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X160 VGND.t30 a_11040_2860.t5 a_13990_2860.t2 VGND.t29 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X161 VDPWR.t368 a_13800_2890.t2 a_13280_3020.t3 VDPWR.t367 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X162 VGND.t226 VGND.t223 VGND.t225 VGND.t224 sky130_fd_pr__nfet_01v8 ad=0.625 pd=3.5 as=0 ps=0 w=1.25 l=0.5
X163 a_17714_9374.t5 a_17714_9374.t4 VDPWR.t100 VDPWR.t99 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X164 VDPWR.t370 a_11430_2890.t2 a_10910_3020.t3 VDPWR.t369 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X165 a_13070_11250.t20 a_15790_17280.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X166 a_13070_11250.t21 a_15790_17280.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X167 VDPWR.t164 a_9450_16252.t18 a_10751_12090.t6 VDPWR.t163 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X168 pll_bgr_magic_3_0.VV1.t3 pll_bgr_magic_3_0.VV2.t1 VGND.t182 sky130_fd_pr__res_xhigh_po_0p35 l=0.86
X169 VDPWR.t160 pll_bgr_magic_3_0.VV3.t5 a_15870_5490.t3 VDPWR.t159 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X170 a_17540_2930.t1 a_17630_3150.t3 VGND.t78 VGND.t77 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X171 a_13360_11960.t5 a_10000_15820.t8 a_13070_11250.t8 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X172 VDPWR.t305 VDPWR.t302 VDPWR.t304 VDPWR.t303 sky130_fd_pr__pfet_01v8 ad=1.25 pd=6 as=0 ps=0 w=2.5 l=0.5
X173 a_13070_11250.t22 a_15790_17280.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X174 a_11200_9430.t27 VDPWR.t241 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X175 a_15320_5490.t1 a_14930_5490.t3 VGND.t244 VGND.t243 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X176 VGND.t165 a_18410_9620.t10 a_18510_9670.t5 VGND.t164 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X177 a_10480_13480.t4 a_11200_9430.t28 VDPWR.t45 VDPWR.t44 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X178 a_12560_13480.t0 a_10480_13480.t0 a_10480_13480.t1 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X179 a_15050_2860.t0 a_15380_3150.t3 VDPWR.t37 VDPWR.t36 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X180 a_12960_8860.t6 a_9450_16252.t19 VDPWR.t166 VDPWR.t165 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X181 pll_bgr_magic_3_0.VV1.t2 a_18390_10330.t6 VGND.t136 VGND.t135 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X182 VGND.t222 VGND.t219 VGND.t221 VGND.t220 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X183 VDPWR.t68 a_19530_10890.t6 pll_bgr_magic_3_0.VV3.t4 VDPWR.t67 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X184 a_11200_9430.t29 VDPWR.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X185 a_15050_2860.t2 a_15160_2860.t5 VGND.t267 VGND.t266 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X186 a_11200_9430.t30 VDPWR.t392 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X187 a_12760_5460.t1 a_12380_5460.t4 VGND.t2 VGND.t1 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X188 V_CONT.t2 a_16000_5490.t4 VDPWR.t139 VDPWR.t138 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X189 VGND.t54 a_13280_5460.t2 a_12760_6640.t0 VGND.t53 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X190 a_10751_12090.t12 VDPWR.t299 VDPWR.t301 VDPWR.t300 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X191 a_11200_9430.t31 VDPWR.t393 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X192 a_10060_12570.t8 a_9570_16200.t8 a_10160_10990.t0 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X193 VDPWR.t23 a_21690_4400.t1 a_21690_4400.t2 VDPWR.t22 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X194 VDPWR.t342 a_15870_5490.t11 a_18390_5940.t2 VDPWR.t341 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X195 a_12380_6640.t2 a_11780_7290.t4 VGND.t271 VGND.t270 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X196 a_15710_5490.t0 a_15320_5490.t3 VDPWR.t56 VDPWR.t16 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X197 VDPWR.t364 a_9450_16252.t20 a_12960_8860.t5 VDPWR.t363 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X198 VDPWR.t237 a_13200_10990.t19 a_13070_11250.t3 VDPWR.t236 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X199 VDPWR.t324 a_12380_5460.t5 a_12300_5910.t0 VDPWR.t151 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X200 VDPWR.t210 a_17030_3180.t3 a_15160_2860.t1 VDPWR.t209 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X201 a_13990_2860.t1 a_11040_2860.t6 VDPWR.t183 VDPWR.t182 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X202 a_15740_2890.t1 a_14690_3160.t2 VGND.t149 VGND.t148 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X203 a_16240_3020.t2 a_15160_2860.t6 VGND.t279 VGND.t278 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X204 VDPWR.t199 a_21690_4400.t3 a_21610_3360.t1 VDPWR.t198 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X205 VGND.t147 a_18930_3150.t5 a_18840_2930.t2 VGND.t146 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X206 a_15870_5490.t12 pll_bgr_magic_3_0.VV2.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X207 VGND.t288 a_13680_6640.t2 a_13280_5460.t1 VGND.t287 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X208 VDPWR.t298 VDPWR.t296 a_11200_9430.t9 VDPWR.t297 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X209 a_11780_5910.t0 ua[0].t0 VDPWR.t140 VDPWR.t69 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X210 a_12070_2860.t2 a_14690_3160.t3 VDPWR.t410 VDPWR.t409 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X211 VDPWR.t185 a_13070_11250.t23 a_11200_9430.t4 VDPWR.t184 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X212 a_17540_2930.t2 a_17630_3150.t4 VGND.t80 VGND.t79 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X213 a_13360_11960.t6 a_10000_15820.t9 a_13070_11250.t7 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X214 a_14930_5490.t1 a_11860_5460.t5 VGND.t138 VGND.t137 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X215 VGND.t217 VGND.t215 VGND.t217 VGND.t216 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X216 VGND.t110 a_18330_3180.t4 a_19550_2800.t1 VGND.t109 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X217 a_15710_6670.t1 a_15320_6670.t4 VDPWR.t17 VDPWR.t16 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X218 VDPWR.t152 a_12380_6640.t5 a_12300_6670.t1 VDPWR.t151 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X219 VDPWR.t156 a_16000_5490.t5 V_CONT.t3 VDPWR.t155 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X220 a_16000_6670.t2 a_15320_6670.t5 VGND.t263 VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X221 a_13200_10990.t5 a_13200_10990.t4 VDPWR.t204 VDPWR.t203 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X222 a_10030_11260.t20 a_9450_17070.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X223 VDPWR.t389 a_14340_6640.t3 a_14010_6640.t1 VDPWR.t388 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X224 a_11780_6670.t1 a_10780_3220.t3 VDPWR.t70 VDPWR.t69 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X225 a_9450_16252.t7 a_10030_11260.t21 VDPWR.t326 VDPWR.t325 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X226 VDPWR.t120 a_11200_9430.t32 a_10480_13480.t3 VDPWR.t119 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X227 VGND.t130 a_20230_3150.t5 a_20140_2930.t1 VGND.t129 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X228 a_18390_5940.t1 a_15870_5490.t13 VDPWR.t124 VDPWR.t123 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X229 a_10030_11260.t22 a_9450_17070.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X230 VDPWR.t170 a_14690_3160.t4 a_15380_3150.t2 VDPWR.t169 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X231 VDPWR.t329 VGND.t304 a_22130_3360.t2 VDPWR.t328 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X232 a_14160_5490.t1 a_13720_5910.t4 VGND.t52 VGND.t51 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X233 VGND.t214 VGND.t211 VGND.t213 VGND.t212 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X234 a_19530_10890.t3 a_19530_10890.t2 VDPWR.t219 VDPWR.t218 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X235 a_13070_11250.t24 a_15790_17280.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X236 a_10910_3020.t1 a_11040_2860.t7 VGND.t191 VGND.t190 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X237 VDPWR.t406 a_11860_5460.t6 a_13720_5910.t2 VDPWR.t405 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X238 a_16240_3020.t3 a_15160_2860.t7 VGND.t290 VGND.t289 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X239 VGND.t176 a_9690_16200.t1 VGND.t95 sky130_fd_pr__res_xhigh_po_0p35 l=3.35
X240 a_11960_2860.t1 a_12070_2860.t11 VGND.t26 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X241 a_11840_9460.t2 a_10480_13480.t6 a_11200_9430.t11 VDPWR.t397 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X242 a_10030_11260.t6 a_10160_10990.t19 VDPWR.t21 VDPWR.t20 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X243 a_13070_11250.t25 a_15790_17280.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X244 VDPWR.t295 VDPWR.t293 a_10751_12090.t11 VDPWR.t294 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X245 VDPWR.t122 a_11200_9430.t33 a_10000_15820.t2 VDPWR.t121 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X246 VDPWR.t98 a_17714_9374.t0 a_17714_9374.t1 VDPWR.t97 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X247 VGND.t38 a_19630_3180.t4 a_20850_2800.t1 VGND.t37 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X248 VGND.t210 VGND.t208 VGND.t210 VGND.t209 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0 ps=0 w=1.25 l=0.5
X249 a_11200_9430.t34 VDPWR.t373 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X250 a_15870_5490.t0 pll_bgr_magic_3_0.VV3.t6 VDPWR.t7 VDPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X251 a_16950_2890.t0 a_15160_2860.t8 a_16650_3100.t0 VGND.t104 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X252 VDPWR.t400 a_20230_3150.t6 a_19630_3180.t0 VDPWR.t399 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X253 a_11200_9430.t0 a_13070_11250.t26 VDPWR.t9 VDPWR.t8 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X254 a_12870_2890.t1 a_11040_2860.t8 a_12540_2890.t0 VGND.t187 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X255 VDPWR.t81 a_19250_3100.t2 a_18840_2930.t3 VDPWR.t80 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X256 VGND.t112 a_18390_10330.t7 pll_bgr_magic_3_0.VV1.t1 VGND.t111 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X257 a_11200_9430.t35 VDPWR.t374 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X258 VGND.t269 a_14690_3160.t5 a_12070_2860.t0 VGND.t268 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X259 a_10160_10990.t10 a_10160_10990.t9 VDPWR.t148 VDPWR.t147 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X260 VDPWR.t35 a_13280_5460.t3 a_13200_5910.t1 VDPWR.t34 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X261 a_10030_11260.t23 a_9450_17070.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X262 VGND.t257 a_20140_2930.t4 a_19630_3180.t1 VGND.t256 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X263 VGND.t189 VDPWR.t427 a_22130_1940.t1 VGND.t159 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X264 VDPWR.t292 VDPWR.t289 VDPWR.t291 VDPWR.t290 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X265 a_13720_5490.t0 a_11860_6640.t6 VGND.t184 VGND.t183 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X266 a_12680_5910.t1 a_11780_5490.t4 VDPWR.t378 VDPWR.t377 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X267 VDPWR.t288 VDPWR.t286 a_12960_8860.t15 VDPWR.t287 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X268 a_10030_11260.t24 a_9450_17070.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X269 a_10910_3020.t0 a_11040_2860.t9 VGND.t167 VGND.t166 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X270 V_CONT.t6 a_16000_5490.t6 VDPWR.t362 VDPWR.t361 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X271 a_11960_2860.t3 a_12290_3150.t3 VDPWR.t15 VDPWR.t14 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X272 a_14340_6640.t0 a_14160_5490.t2 VDPWR.t247 VDPWR.t246 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X273 VDPWR.t66 a_18330_3180.t5 a_17630_3150.t0 VDPWR.t65 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X274 a_11840_9460.t6 a_11200_9430.t36 VDPWR.t227 VDPWR.t226 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X275 a_11960_2860.t0 a_12070_2860.t12 VGND.t119 VGND.t118 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X276 a_13200_10990.t3 a_13200_10990.t2 VDPWR.t19 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X277 a_13360_11960.t10 a_11840_9460.t9 a_13200_10990.t16 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X278 a_13070_11250.t27 a_15790_17280.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X279 VDPWR.t366 a_9450_16252.t21 a_10751_12090.t5 VDPWR.t365 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X280 VDPWR.t50 pll_bgr_magic_3_0.VV3.t7 a_15870_5490.t2 VDPWR.t49 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X281 a_13070_11250.t28 a_15790_17280.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X282 VDPWR.t394 a_13280_5460.t4 a_13200_6670.t1 VDPWR.t34 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X283 VDPWR.t381 a_20550_3100.t2 a_20140_2930.t3 VDPWR.t380 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X284 VGND.t207 VGND.t204 VGND.t206 VGND.t205 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X285 a_18840_2930.t1 a_18930_3150.t6 VGND.t140 VGND.t139 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X286 a_12290_3150.t1 a_11040_2860.t10 VDPWR.t75 VDPWR.t74 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X287 a_12680_6670.t1 a_11780_7290.t5 VDPWR.t411 VDPWR.t377 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X288 a_13070_11250.t2 a_13200_10990.t20 VDPWR.t195 VDPWR.t194 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X289 a_13360_11960.t1 a_11840_9460.t10 a_13200_10990.t13 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X290 a_13070_11250.t29 a_15790_17280.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X291 VGND.t66 a_10780_3220.t4 a_12540_2890.t1 VGND.t65 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X292 a_9570_16200.t1 a_11200_9430.t37 VDPWR.t229 VDPWR.t228 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X293 a_11200_9430.t38 VDPWR.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X294 a_10030_11260.t5 a_10160_10990.t20 VDPWR.t77 VDPWR.t76 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X295 a_20230_3150.t2 ua1.t3 VDPWR.t177 VDPWR.t176 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X296 VDPWR.t396 a_14690_3160.t6 a_12070_2860.t1 VDPWR.t395 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X297 VDPWR.t130 a_13680_6640.t3 a_13280_5460.t0 VDPWR.t129 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X298 a_18160_10940.t2 a_18160_10940.t1 a_18160_10940.t2 VDPWR.t82 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X299 a_16000_5490.t1 a_15320_5490.t4 VDPWR.t231 VDPWR.t230 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X300 a_11200_9430.t39 VDPWR.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X301 a_15870_5490.t14 pll_bgr_magic_3_0.VV4.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X302 VDPWR.t285 VDPWR.t282 VDPWR.t284 VDPWR.t283 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X303 a_10030_11260.t25 a_9450_17070.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X304 a_15790_17280.t20 a_11200_9430.t2 VGND.t33 sky130_fd_pr__res_high_po_0p35 l=2.05
X305 a_10160_10990.t8 a_10160_10990.t7 VDPWR.t193 VDPWR.t192 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X306 VDPWR.t281 VDPWR.t278 VDPWR.t280 VDPWR.t279 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X307 a_11200_9430.t40 VDPWR.t414 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X308 a_10160_10990.t1 a_9570_16200.t9 a_10060_12570.t7 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X309 a_11840_9460.t5 a_11200_9430.t41 VDPWR.t416 VDPWR.t415 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X310 a_18390_10330.t1 a_18390_10330.t0 VGND.t186 VGND.t185 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X311 VDPWR.t233 a_19530_10890.t0 a_19530_10890.t1 VDPWR.t232 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X312 a_21720_2700.t0 ua1.t4 a_21610_1940.t2 VGND.t94 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X313 a_11200_9430.t3 a_13070_11250.t30 VDPWR.t85 VDPWR.t84 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X314 VDPWR.t327 VGND.t305 a_22650_3360.t1 VDPWR.t238 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X315 a_10030_11260.t26 a_9450_17070.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X316 a_16000_5490.t7 a_15710_5490.t2 sky130_fd_pr__cap_mim_m3_1 l=6.3 w=5.2
X317 VDPWR.t39 a_9450_16252.t22 a_10751_12090.t4 VDPWR.t38 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X318 a_10160_10990.t6 a_10160_10990.t5 VDPWR.t60 VDPWR.t59 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X319 a_10000_17428.t1 a_10120_15820.t0 VGND.t27 sky130_fd_pr__res_xhigh_po_0p35 l=6
X320 VDPWR.t235 a_21690_4400.t4 a_22130_3360.t1 VDPWR.t234 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X321 a_15710_5490.t1 a_15320_5490.t5 VGND.t273 VGND.t272 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X322 a_13070_11250.t31 a_15790_17280.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X323 VGND.t297 a_12380_5460.t6 a_11860_5460.t0 VGND.t296 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X324 VGND.t193 VGND.t194 a_10900_14480.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X325 a_10160_10990.t3 a_9570_16200.t10 a_10060_12570.t6 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X326 VDPWR.t87 a_11200_9430.t42 a_11840_9460.t4 VDPWR.t86 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X327 a_12650_3210.t0 a_10780_3220.t5 a_12290_3150.t0 VDPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X328 a_11780_5490.t0 ua[0].t1 VGND.t117 VGND.t116 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X329 VGND.t90 a_11860_6640.t7 a_11780_7290.t2 VGND.t89 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X330 a_9450_16252.t3 a_10030_11260.t27 VDPWR.t221 VDPWR.t220 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X331 VGND.t282 a_13990_2860.t3 a_13910_2890.t1 VGND.t281 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X332 VGND.t280 a_12560_13480.t1 a_12560_13480.t0 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X333 VGND.t36 a_10780_3220.t6 a_11540_2890.t1 VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X334 a_10900_14480.t0 a_10000_15820.t5 VGND.t181 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X335 a_11200_9430.t43 VDPWR.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X336 VGND.t84 a_18410_9620.t4 a_18410_9620.t5 VGND.t83 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X337 a_17630_3150.t2 a_18330_3180.t6 VGND.t134 VGND.t133 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X338 a_9570_17278.t0 a_9690_16200.t0 VGND.t95 sky130_fd_pr__res_xhigh_po_0p35 l=3.35
X339 VDPWR.t41 a_9450_16252.t23 a_12960_8860.t4 VDPWR.t40 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X340 VDPWR.t31 a_11200_9430.t44 a_9570_16200.t0 VDPWR.t30 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X341 a_18510_9670.t10 a_18510_9670.t8 a_18510_9670.t9 VGND.t155 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X342 a_17714_9374.t8 a_18410_9620.t8 sky130_fd_pr__res_generic_po w=0.33 l=2.4
X343 a_10160_10990.t2 a_9570_16200.t11 a_10060_12570.t5 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X344 a_9450_16252.t4 VDPWR.t275 VDPWR.t277 VDPWR.t276 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X345 VGND.t57 VDPWR.t428 a_22650_1940.t1 VGND.t46 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X346 a_18160_10940.t12 V_CONT.t13 a_18390_10330.t4 VDPWR.t332 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X347 a_10030_11260.t28 a_9450_17070.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X348 VGND.t82 a_18410_9620.t2 a_18410_9620.t3 VGND.t81 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X349 a_13360_11960.t7 VDPWR.t429 VGND.t59 VGND.t58 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1.01 ps=6.15 w=2.5 l=5
X350 VDPWR.t223 a_9450_16252.t24 a_10751_12090.t3 VDPWR.t222 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X351 VDPWR.t323 a_19630_3180.t5 a_18930_3150.t1 VDPWR.t322 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X352 VDPWR.t162 a_15160_2860.t9 a_15820_2860.t1 VDPWR.t161 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X353 a_13720_5910.t1 a_11860_5460.t7 a_13720_5490.t1 VGND.t113 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X354 a_11860_6640.t2 a_11780_7290.t6 VGND.t294 VGND.t293 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X355 VDPWR.t274 VDPWR.t272 VDPWR.t274 VDPWR.t273 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X356 a_11200_9430.t1 a_13070_11250.t32 VDPWR.t43 VDPWR.t42 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X357 VGND.t284 a_12070_2860.t13 a_13280_3020.t0 VGND.t283 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X358 VDPWR.t33 a_11200_9430.t45 a_11840_9460.t3 VDPWR.t32 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X359 a_13200_10990.t14 a_11840_9460.t11 a_13360_11960.t8 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X360 VGND.t247 a_10910_3020.t4 a_10780_3220.t1 VGND.t246 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X361 VGND.t4 a_12960_8860.t13 a_12960_8860.t14 VGND.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X362 VGND.t76 pll_bgr_magic_3_0.VV1.t7 a_15870_5490.t6 VGND.t75 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X363 VGND.t8 a_18410_9620.t11 a_18510_9670.t0 VGND.t7 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X364 VDPWR.t96 a_17714_9374.t11 a_18160_10940.t8 VDPWR.t95 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X365 a_15160_2860.t2 a_17030_3180.t4 VGND.t97 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X366 a_13800_2890.t1 a_13990_2860.t4 VDPWR.t408 VDPWR.t407 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X367 VGND.t132 a_11960_2860.t4 a_11040_2860.t1 VGND.t131 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X368 a_11430_2890.t1 a_10780_3220.t7 VDPWR.t154 VDPWR.t153 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X369 a_10751_12090.t2 a_9450_16252.t25 VDPWR.t225 VDPWR.t224 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X370 a_18510_9670.t2 a_18390_5940.t8 pll_bgr_magic_3_0.VV3.t0 VGND.t93 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X371 a_16000_6670.t0 a_15710_6670.t3 a_12960_8860.t0 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X372 a_17714_9374.t7 a_17714_9374.t6 VDPWR.t94 VDPWR.t93 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X373 a_18250_2800.t1 a_17630_3150.t5 a_17950_3100.t1 VGND.t245 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X374 a_10030_11260.t29 a_9450_17070.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X375 a_10030_11260.t1 a_10751_12090.t16 a_10060_12570.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X376 a_17950_3100.t0 a_17030_3180.t5 VDPWR.t158 VDPWR.t157 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X377 VDPWR.t271 VDPWR.t269 a_9570_16200.t5 VDPWR.t270 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X378 VDPWR.t418 a_9450_16252.t26 a_12960_8860.t3 VDPWR.t417 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X379 a_13200_10990.t1 a_13200_10990.t0 VDPWR.t146 VDPWR.t145 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X380 VGND.t255 a_15160_2860.t10 a_15050_2860.t1 VGND.t254 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X381 a_15870_5490.t9 pll_bgr_magic_3_0.VV3.t8 VDPWR.t391 VDPWR.t390 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X382 a_21720_2700.t1 ua1.t5 a_21610_3360.t2 VDPWR.t330 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X383 VDPWR.t114 ua1.t6 a_20230_3150.t1 VDPWR.t113 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X384 VGND.t87 a_14770_15820.t0 VGND.t86 sky130_fd_pr__res_xhigh_po_0p35 l=6
X385 a_10030_11260.t30 a_9450_17070.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X386 VGND.t99 a_13280_5460.t5 a_12760_5460.t2 VGND.t98 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X387 VDPWR.t217 a_16650_3100.t2 a_16240_3020.t1 VDPWR.t216 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X388 VDPWR.t420 a_9450_16252.t27 a_10751_12090.t1 VDPWR.t419 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X389 a_18510_9670.t4 a_18410_9620.t12 VGND.t161 VGND.t160 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X390 a_10030_11260.t31 a_9450_17070.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X391 pll_bgr_magic_3_0.VV3.t3 a_19530_10890.t7 VDPWR.t387 VDPWR.t386 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X392 a_10030_11260.t10 a_10751_12090.t17 a_10060_12570.t0 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X393 a_10000_15820.t1 a_11200_9430.t46 VDPWR.t27 VDPWR.t26 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X394 a_12380_5460.t2 a_11780_5490.t5 VGND.t275 VGND.t274 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X395 a_13070_11250.t1 a_13200_10990.t21 VDPWR.t376 VDPWR.t375 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X396 a_14340_6640.t1 a_14160_5490.t3 VGND.t20 VGND.t19 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X397 VGND.t172 a_12760_6640.t4 a_12380_6640.t1 VGND.t171 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X398 a_12960_8860.t2 a_9450_16252.t28 VDPWR.t354 VDPWR.t353 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X399 a_13200_10990.t12 a_11840_9460.t12 a_13360_11960.t0 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X400 VGND.t103 V_CONT.t14 a_21610_1940.t1 VGND.t94 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X401 a_13070_11250.t33 a_15790_17280.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X402 VGND.t68 a_13280_3020.t4 a_12700_3340.t0 VGND.t67 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X403 VDPWR.t268 VDPWR.t266 VDPWR.t268 VDPWR.t267 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X404 a_10030_11260.t4 a_10160_10990.t21 VDPWR.t206 VDPWR.t205 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X405 a_15160_2860.t0 a_17030_3180.t6 VDPWR.t372 VDPWR.t371 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X406 a_12960_8860.t12 a_12960_8860.t11 VGND.t40 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X407 a_15850_2890.t0 a_15820_2860.t2 a_15740_2890.t0 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X408 a_18840_2930.t0 a_18930_3150.t7 VGND.t142 VGND.t141 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X409 VDPWR.t250 a_21690_4400.t5 a_22650_3360.t2 VDPWR.t249 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X410 VGND.t64 a_14010_6640.t3 a_13680_6640.t1 VGND.t63 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X411 VGND.t203 VGND.t200 VGND.t202 VGND.t201 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X412 a_18410_9620.t1 a_18410_9620.t0 VGND.t259 VGND.t258 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X413 a_13070_11250.t34 a_15790_17280.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X414 a_11780_5490.t1 a_11860_5460.t8 a_11780_5910.t1 VDPWR.t55 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X415 a_9570_16200.t4 VDPWR.t263 VDPWR.t265 VDPWR.t264 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X416 VGND.t193 VGND.t192 a_10900_14480.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X417 a_10480_13480.t2 a_11200_9430.t47 VDPWR.t29 VDPWR.t28 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X418 VGND.t108 a_17630_3150.t6 a_17540_2930.t3 VGND.t107 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X419 VGND.t193 VGND.t199 a_10900_14480.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X420 VDPWR.t11 a_10030_11260.t32 a_9450_16252.t0 VDPWR.t10 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X421 a_11200_9430.t48 VDPWR.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X422 VDPWR.t126 a_12070_2860.t14 a_12700_3340.t1 VDPWR.t125 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X423 a_15320_6670.t0 VDPWR.t430 a_14930_6670.t3 VGND.t250 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X424 VDPWR.t352 a_15160_2860.t11 a_14690_3160.t0 VDPWR.t351 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X425 a_14890_17428.t0 a_11840_9460.t0 VGND.t22 sky130_fd_pr__res_xhigh_po_0p35 l=6
X426 VDPWR.t356 a_9450_16252.t29 a_12960_8860.t1 VDPWR.t355 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X427 a_11200_9430.t8 VDPWR.t260 VDPWR.t262 VDPWR.t261 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X428 a_18930_3150.t2 a_19630_3180.t6 VGND.t299 VGND.t298 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X429 a_11200_9430.t49 VDPWR.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X430 VGND.t122 a_15050_2860.t4 a_14690_3160.t1 VGND.t121 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X431 a_19530_10890.t4 V_CONT.t15 a_18510_9670.t6 VGND.t48 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X432 VDPWR.t259 VDPWR.t257 VDPWR.t259 VDPWR.t258 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0 ps=0 w=2.5 l=0.5
X433 a_12760_6640.t2 a_12380_6640.t6 VGND.t261 VGND.t260 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X434 a_10030_11260.t33 a_9450_17070.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X435 a_11780_7290.t1 a_11860_6640.t8 a_11780_6670.t0 VDPWR.t55 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X436 VDPWR.t197 a_10160_10990.t22 a_10030_11260.t3 VDPWR.t196 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X437 pll_bgr_magic_3_0.VV1.t0 a_18390_5940.t9 a_18160_10940.t0 VDPWR.t5 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X438 a_20140_2930.t0 a_20230_3150.t7 VGND.t154 VGND.t153 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X439 a_15288_18640.t0 V_CONT.t4 VGND.t156 sky130_fd_pr__res_xhigh_po_0p35 l=7.52
X440 a_10030_11260.t34 a_9450_17070.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X441 pll_bgr_magic_3_0.VV4.t1 pll_bgr_magic_3_0.VV3.t2 VGND.t43 sky130_fd_pr__res_xhigh_po_0p35 l=1.14
X442 a_22240_2700.t0 a_21720_2700.t3 a_22130_1940.t0 VGND.t159 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X443 a_15380_3150.t0 a_15820_2860.t3 VDPWR.t385 VDPWR.t384 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X444 a_10030_11260.t35 a_9450_17070.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X445 VDPWR.t168 a_17630_3150.t7 a_17030_3180.t0 VDPWR.t167 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X446 a_12300_5910.t1 a_11780_5490.t6 a_11860_5460.t2 VDPWR.t379 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X447 VDPWR.t62 a_11040_2860.t11 a_13990_2860.t0 VDPWR.t61 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X448 VGND.t14 a_15160_2860.t12 a_16240_3020.t0 VGND.t13 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X449 a_13070_11250.t35 a_15790_17280.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X450 a_11200_9430.t7 VDPWR.t254 VDPWR.t256 VDPWR.t255 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.45 ps=2.9 w=1 l=0.15
X451 a_10030_11260.t36 a_9450_17070.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X452 VGND.t198 VGND.t196 VGND.t198 VGND.t197 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X453 a_11200_9430.t12 a_10480_13480.t7 a_11840_9460.t1 VDPWR.t398 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X454 a_15870_5490.t5 pll_bgr_magic_3_0.VV1.t8 VGND.t10 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X455 VDPWR.t253 VDPWR.t251 a_11200_9430.t6 VDPWR.t252 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X456 a_13070_11250.t6 a_10000_15820.t10 a_13360_11960.t3 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X457 a_18160_10940.t9 a_17714_9374.t12 VDPWR.t92 VDPWR.t91 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X458 a_13070_11250.t36 a_15790_17280.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X459 a_16000_5490.t2 a_15710_5490.t3 a_15870_5490.t4 VDPWR.t200 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X460 VGND.t193 VGND.t195 a_10900_14480.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X461 VDPWR.t383 a_15870_5490.t15 a_18390_5940.t0 VDPWR.t382 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X462 VGND.t6 a_17540_2930.t4 a_17030_3180.t1 VGND.t5 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X463 a_13070_11250.t0 a_13200_10990.t22 VDPWR.t58 VDPWR.t57 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
R0 VGND.n686 VGND.n586 1.28274e+06
R1 VGND.n687 VGND.n686 462138
R2 VGND.n950 VGND.n949 193700
R3 VGND.n687 VGND.t55 132039
R4 VGND.n710 VGND.n586 132000
R5 VGND.n949 VGND.n586 42900
R6 VGND.n739 VGND.t43 14832.4
R7 VGND.n710 VGND.n709 11603.1
R8 VGND.n898 VGND.n870 11250
R9 VGND.n950 VGND.n585 9511.11
R10 VGND.n712 VGND.n710 9155.25
R11 VGND.n896 VGND.n871 8618.75
R12 VGND.n896 VGND.n872 8323.25
R13 VGND.n952 VGND.n951 8289.79
R14 VGND.n882 VGND.n871 6796.5
R15 VGND.n870 VGND.n738 6739.68
R16 VGND.n882 VGND.n872 6501
R17 VGND.n686 VGND.n672 4738.46
R18 VGND.n951 VGND.n950 4657.55
R19 VGND.n685 VGND.n585 4106.67
R20 VGND.n953 VGND.n952 3870.38
R21 VGND.n682 VGND.n585 3748.15
R22 VGND.n845 VGND.n738 2923.95
R23 VGND.n952 VGND.n583 2834.83
R24 VGND.n881 VGND.n870 2777.59
R25 VGND.n739 VGND.n582 2623.32
R26 VGND.n949 VGND.t246 2620.22
R27 VGND.n949 VGND.n662 2351.73
R28 VGND.n738 VGND.t12 2080.51
R29 VGND.n870 VGND.n869 1503.36
R30 VGND.n923 VGND.n922 1217.93
R31 VGND.n911 VGND.n910 1217.93
R32 VGND.n909 VGND.n908 1217.93
R33 VGND.n954 VGND.n953 1192.53
R34 VGND.n868 VGND.n867 1192.53
R35 VGND.n759 VGND.n758 1186
R36 VGND.n857 VGND.n856 1186
R37 VGND.n772 VGND.n771 1186
R38 VGND.t162 VGND.n866 1186
R39 VGND.n948 VGND.n947 1182.8
R40 VGND.n925 VGND.n924 1182.8
R41 VGND.n2352 VGND.n2351 1182.66
R42 VGND.n961 VGND.n960 1182.66
R43 VGND.t260 VGND.t171 1054.97
R44 VGND.t89 VGND.t293 1054.97
R45 VGND.n582 VGND.t156 1019.28
R46 VGND.n492 VGND.n481 893.807
R47 VGND.n845 VGND.n760 871.141
R48 VGND.t169 VGND.t46 846.154
R49 VGND.n953 VGND.n582 833.124
R50 VGND.t159 VGND.t94 733.333
R51 VGND.t127 VGND.t1 724.499
R52 VGND.t31 VGND.t179 724.499
R53 VGND.n958 VGND.n957 686.717
R54 VGND.n958 VGND.n579 686.717
R55 VGND.n880 VGND.t159 683.975
R56 VGND.t123 VGND.t250 683.665
R57 VGND.n696 VGND.t287 681.871
R58 VGND.n841 VGND.n840 669.307
R59 VGND.n818 VGND.n817 669.307
R60 VGND.n820 VGND.n809 669.307
R61 VGND.n793 VGND.n745 669.307
R62 VGND.n789 VGND.n746 669.307
R63 VGND.n654 VGND.t88 656.367
R64 VGND.n963 VGND.n461 654.447
R65 VGND.t193 VGND.t88 628.787
R66 VGND.n619 VGND.n588 609.484
R67 VGND.n843 VGND.n583 596.899
R68 VGND.n715 VGND.n713 585.003
R69 VGND.n707 VGND.n706 585.003
R70 VGND.n709 VGND.n708 585.001
R71 VGND.n697 VGND.n696 585.001
R72 VGND.n695 VGND.n694 585.001
R73 VGND.n693 VGND.n692 585.001
R74 VGND.n689 VGND.n688 585.001
R75 VGND.n860 VGND.n858 585.001
R76 VGND.n847 VGND.n846 585.001
R77 VGND.n684 VGND.n683 585.001
R78 VGND.n737 VGND.n736 585.001
R79 VGND.n734 VGND.n733 585.001
R80 VGND.n732 VGND.n731 585.001
R81 VGND.n730 VGND.n729 585.001
R82 VGND.n726 VGND.n725 585.001
R83 VGND.n724 VGND.n723 585.001
R84 VGND.n722 VGND.n721 585.001
R85 VGND.n712 VGND.n711 585.001
R86 VGND.n677 VGND.n676 585.001
R87 VGND.n681 VGND.n680 585.001
R88 VGND.n797 VGND.n796 585
R89 VGND.n799 VGND.n798 585
R90 VGND.n813 VGND.n812 585
R91 VGND.n822 VGND.n821 585
R92 VGND.n780 VGND.n767 585
R93 VGND.n773 VGND.n767 585
R94 VGND.n769 VGND.n766 585
R95 VGND.n776 VGND.n775 585
R96 VGND.n768 VGND.n765 585
R97 VGND.n773 VGND.n768 585
R98 VGND.n2272 VGND.n2271 585
R99 VGND.n2273 VGND.n1685 585
R100 VGND.n2275 VGND.n2274 585
R101 VGND.n2277 VGND.n1683 585
R102 VGND.n2279 VGND.n2278 585
R103 VGND.n2280 VGND.n1682 585
R104 VGND.n2282 VGND.n2281 585
R105 VGND.n2284 VGND.n1680 585
R106 VGND.n2286 VGND.n2285 585
R107 VGND.n2287 VGND.n1679 585
R108 VGND.n2289 VGND.n2288 585
R109 VGND.n2291 VGND.n1672 585
R110 VGND.n1466 VGND.n1465 585
R111 VGND.n1463 VGND.n1300 585
R112 VGND.n1354 VGND.n1353 585
R113 VGND.n1458 VGND.n1457 585
R114 VGND.n1456 VGND.n1455 585
R115 VGND.n1382 VGND.n1358 585
R116 VGND.n1384 VGND.n1383 585
R117 VGND.n1389 VGND.n1388 585
R118 VGND.n1387 VGND.n1380 585
R119 VGND.n1395 VGND.n1394 585
R120 VGND.n1397 VGND.n1396 585
R121 VGND.n1378 VGND.n1377 585
R122 VGND.n1182 VGND.n102 585
R123 VGND.n1293 VGND.n1292 585
R124 VGND.n1184 VGND.n1181 585
R125 VGND.n1287 VGND.n1286 585
R126 VGND.n1285 VGND.n1284 585
R127 VGND.n1210 VGND.n1188 585
R128 VGND.n1212 VGND.n1211 585
R129 VGND.n1217 VGND.n1216 585
R130 VGND.n1215 VGND.n1208 585
R131 VGND.n1223 VGND.n1222 585
R132 VGND.n1225 VGND.n1224 585
R133 VGND.n1175 VGND.n109 585
R134 VGND.n108 VGND.n107 585
R135 VGND.n1545 VGND.n1482 585
R136 VGND.n1555 VGND.n1554 585
R137 VGND.n1557 VGND.n1480 585
R138 VGND.n1560 VGND.n1559 585
R139 VGND.n1561 VGND.n1476 585
R140 VGND.n1570 VGND.n1569 585
R141 VGND.n1572 VGND.n1475 585
R142 VGND.n1575 VGND.n1574 585
R143 VGND.n1576 VGND.n1469 585
R144 VGND.n1585 VGND.n1584 585
R145 VGND.n1587 VGND.n1174 585
R146 VGND.n2332 VGND.n2331 585
R147 VGND.n74 VGND.n72 585
R148 VGND.n1310 VGND.n1309 585
R149 VGND.n1312 VGND.n1311 585
R150 VGND.n1314 VGND.n1313 585
R151 VGND.n1316 VGND.n1315 585
R152 VGND.n1318 VGND.n1317 585
R153 VGND.n1320 VGND.n1319 585
R154 VGND.n1322 VGND.n1321 585
R155 VGND.n1324 VGND.n1323 585
R156 VGND.n1326 VGND.n1325 585
R157 VGND.n1327 VGND.n1308 585
R158 VGND.n143 VGND.n122 585
R159 VGND.n142 VGND.n141 585
R160 VGND.n140 VGND.n139 585
R161 VGND.n138 VGND.n137 585
R162 VGND.n136 VGND.n135 585
R163 VGND.n134 VGND.n133 585
R164 VGND.n132 VGND.n131 585
R165 VGND.n130 VGND.n129 585
R166 VGND.n128 VGND.n127 585
R167 VGND.n126 VGND.n125 585
R168 VGND.n124 VGND.n123 585
R169 VGND.n78 VGND.n75 585
R170 VGND.n1613 VGND.n1612 585
R171 VGND.n1615 VGND.n1614 585
R172 VGND.n1617 VGND.n1616 585
R173 VGND.n1619 VGND.n1618 585
R174 VGND.n1621 VGND.n1620 585
R175 VGND.n1623 VGND.n1622 585
R176 VGND.n1625 VGND.n1624 585
R177 VGND.n1627 VGND.n1626 585
R178 VGND.n1629 VGND.n1628 585
R179 VGND.n1631 VGND.n1630 585
R180 VGND.n1633 VGND.n1632 585
R181 VGND.n1635 VGND.n1634 585
R182 VGND.n1066 VGND.n1065 585
R183 VGND.n1090 VGND.n1068 585
R184 VGND.n1092 VGND.n1091 585
R185 VGND.n1088 VGND.n1087 585
R186 VGND.n1086 VGND.n1085 585
R187 VGND.n1081 VGND.n1080 585
R188 VGND.n1079 VGND.n1078 585
R189 VGND.n1074 VGND.n1073 585
R190 VGND.n1072 VGND.n360 585
R191 VGND.n1100 VGND.n1099 585
R192 VGND.n1102 VGND.n1101 585
R193 VGND.n1105 VGND.n1104 585
R194 VGND.n1116 VGND.n1115 585
R195 VGND.n1120 VGND.n1119 585
R196 VGND.n1118 VGND.n288 585
R197 VGND.n1127 VGND.n1126 585
R198 VGND.n1129 VGND.n1128 585
R199 VGND.n1132 VGND.n1131 585
R200 VGND.n1130 VGND.n284 585
R201 VGND.n1141 VGND.n1140 585
R202 VGND.n1143 VGND.n1142 585
R203 VGND.n1144 VGND.n278 585
R204 VGND.n1154 VGND.n1153 585
R205 VGND.n1151 VGND.n277 585
R206 VGND.n1158 VGND.n147 585
R207 VGND.n255 VGND.n148 585
R208 VGND.n264 VGND.n263 585
R209 VGND.n156 VGND.n154 585
R210 VGND.n181 VGND.n180 585
R211 VGND.n186 VGND.n185 585
R212 VGND.n184 VGND.n178 585
R213 VGND.n193 VGND.n192 585
R214 VGND.n191 VGND.n177 585
R215 VGND.n199 VGND.n198 585
R216 VGND.n201 VGND.n200 585
R217 VGND.n149 VGND.n21 585
R218 VGND.n541 VGND.n540 585
R219 VGND.n542 VGND.n538 585
R220 VGND.n543 VGND.n537 585
R221 VGND.n535 VGND.n532 585
R222 VGND.n549 VGND.n531 585
R223 VGND.n550 VGND.n529 585
R224 VGND.n551 VGND.n528 585
R225 VGND.n526 VGND.n524 585
R226 VGND.n556 VGND.n523 585
R227 VGND.n557 VGND.n521 585
R228 VGND.n520 VGND.n470 585
R229 VGND.n562 VGND.n468 585
R230 VGND.n1160 VGND.n145 585
R231 VGND.n145 VGND.n38 585
R232 VGND.n562 VGND.n561 585
R233 VGND.n559 VGND.n470 585
R234 VGND.n558 VGND.n557 585
R235 VGND.n556 VGND.n555 585
R236 VGND.n554 VGND.n524 585
R237 VGND.n552 VGND.n551 585
R238 VGND.n550 VGND.n525 585
R239 VGND.n549 VGND.n548 585
R240 VGND.n546 VGND.n532 585
R241 VGND.n544 VGND.n543 585
R242 VGND.n542 VGND.n534 585
R243 VGND.n541 VGND.n146 585
R244 VGND.n1160 VGND.n1159 585
R245 VGND.n1159 VGND.n38 585
R246 VGND.n1670 VGND.n1669 585
R247 VGND.n1667 VGND.n110 585
R248 VGND.n1666 VGND.n1665 585
R249 VGND.n1654 VGND.n112 585
R250 VGND.n1655 VGND.n115 585
R251 VGND.n1658 VGND.n1657 585
R252 VGND.n1653 VGND.n117 585
R253 VGND.n1651 VGND.n1650 585
R254 VGND.n119 VGND.n118 585
R255 VGND.n1644 VGND.n1643 585
R256 VGND.n1641 VGND.n121 585
R257 VGND.n1639 VGND.n1638 585
R258 VGND.n2302 VGND.n105 585
R259 VGND.n2304 VGND.n105 585
R260 VGND.n1638 VGND.n1637 585
R261 VGND.n121 VGND.n120 585
R262 VGND.n1645 VGND.n1644 585
R263 VGND.n1647 VGND.n119 585
R264 VGND.n1650 VGND.n1649 585
R265 VGND.n117 VGND.n116 585
R266 VGND.n1659 VGND.n1658 585
R267 VGND.n1661 VGND.n115 585
R268 VGND.n1662 VGND.n112 585
R269 VGND.n1665 VGND.n1664 585
R270 VGND.n114 VGND.n110 585
R271 VGND.n1670 VGND.n106 585
R272 VGND.n2303 VGND.n2302 585
R273 VGND.n2304 VGND.n2303 585
R274 VGND.n2193 VGND.n1778 585
R275 VGND.n2196 VGND.n2195 585
R276 VGND.n1807 VGND.n1780 585
R277 VGND.n1805 VGND.n1804 585
R278 VGND.n1782 VGND.n1781 585
R279 VGND.n1798 VGND.n1797 585
R280 VGND.n1795 VGND.n1784 585
R281 VGND.n1793 VGND.n1792 585
R282 VGND.n1787 VGND.n1786 585
R283 VGND.n1677 VGND.n1676 585
R284 VGND.n2296 VGND.n2295 585
R285 VGND.n2298 VGND.n1673 585
R286 VGND.n2292 VGND.n1673 585
R287 VGND.n2295 VGND.n2294 585
R288 VGND.n1678 VGND.n1677 585
R289 VGND.n1789 VGND.n1787 585
R290 VGND.n1792 VGND.n1791 585
R291 VGND.n1784 VGND.n1783 585
R292 VGND.n1799 VGND.n1798 585
R293 VGND.n1801 VGND.n1782 585
R294 VGND.n1804 VGND.n1803 585
R295 VGND.n1780 VGND.n1779 585
R296 VGND.n2197 VGND.n2196 585
R297 VGND.n2199 VGND.n1778 585
R298 VGND.n2300 VGND.n2299 585
R299 VGND.n2025 VGND.n1674 585
R300 VGND.n2027 VGND.n2026 585
R301 VGND.n2029 VGND.n2023 585
R302 VGND.n2031 VGND.n2030 585
R303 VGND.n2032 VGND.n2022 585
R304 VGND.n2034 VGND.n2033 585
R305 VGND.n2036 VGND.n2020 585
R306 VGND.n2038 VGND.n2037 585
R307 VGND.n2039 VGND.n2019 585
R308 VGND.n2041 VGND.n2040 585
R309 VGND.n2043 VGND.n2018 585
R310 VGND.n2052 VGND.n2051 585
R311 VGND.n2053 VGND.n1976 585
R312 VGND.n2055 VGND.n2054 585
R313 VGND.n2057 VGND.n1974 585
R314 VGND.n2059 VGND.n2058 585
R315 VGND.n2060 VGND.n1973 585
R316 VGND.n2062 VGND.n2061 585
R317 VGND.n2064 VGND.n1971 585
R318 VGND.n2066 VGND.n2065 585
R319 VGND.n2067 VGND.n1970 585
R320 VGND.n2069 VGND.n2068 585
R321 VGND.n2071 VGND.n1969 585
R322 VGND.n1998 VGND.n1886 585
R323 VGND.n1999 VGND.n1997 585
R324 VGND.n2004 VGND.n1995 585
R325 VGND.n2005 VGND.n1993 585
R326 VGND.n2006 VGND.n1992 585
R327 VGND.n1990 VGND.n1988 585
R328 VGND.n2012 VGND.n1987 585
R329 VGND.n2013 VGND.n1985 585
R330 VGND.n2014 VGND.n1984 585
R331 VGND.n1981 VGND.n1980 585
R332 VGND.n2048 VGND.n2047 585
R333 VGND.n2050 VGND.n1979 585
R334 VGND.n2044 VGND.n1979 585
R335 VGND.n2047 VGND.n2046 585
R336 VGND.n2017 VGND.n1981 585
R337 VGND.n2015 VGND.n2014 585
R338 VGND.n2013 VGND.n1982 585
R339 VGND.n2012 VGND.n2011 585
R340 VGND.n2009 VGND.n1988 585
R341 VGND.n2007 VGND.n2006 585
R342 VGND.n2005 VGND.n1989 585
R343 VGND.n2004 VGND.n2003 585
R344 VGND.n2001 VGND.n1999 585
R345 VGND.n1998 VGND.n1885 585
R346 VGND.n2308 VGND.n100 585
R347 VGND.n2309 VGND.n98 585
R348 VGND.n2310 VGND.n97 585
R349 VGND.n95 VGND.n93 585
R350 VGND.n2316 VGND.n92 585
R351 VGND.n2317 VGND.n90 585
R352 VGND.n2318 VGND.n89 585
R353 VGND.n87 VGND.n85 585
R354 VGND.n2323 VGND.n84 585
R355 VGND.n2324 VGND.n82 585
R356 VGND.n81 VGND.n77 585
R357 VGND.n2329 VGND.n73 585
R358 VGND.n104 VGND.n103 585
R359 VGND.n2304 VGND.n104 585
R360 VGND.n2329 VGND.n2328 585
R361 VGND.n2326 VGND.n77 585
R362 VGND.n2325 VGND.n2324 585
R363 VGND.n2323 VGND.n2322 585
R364 VGND.n2321 VGND.n85 585
R365 VGND.n2319 VGND.n2318 585
R366 VGND.n2317 VGND.n86 585
R367 VGND.n2316 VGND.n2315 585
R368 VGND.n2313 VGND.n93 585
R369 VGND.n2311 VGND.n2310 585
R370 VGND.n2309 VGND.n94 585
R371 VGND.n2308 VGND.n2307 585
R372 VGND.n2305 VGND.n103 585
R373 VGND.n2305 VGND.n2304 585
R374 VGND.n1106 VGND.n76 585
R375 VGND.n1106 VGND.n38 585
R376 VGND.n1114 VGND.n76 585
R377 VGND.n1114 VGND.n38 585
R378 VGND.n1107 VGND.n354 585
R379 VGND.n1110 VGND.n1109 585
R380 VGND.n357 VGND.n356 585
R381 VGND.n997 VGND.n996 585
R382 VGND.n1002 VGND.n994 585
R383 VGND.n1003 VGND.n992 585
R384 VGND.n1004 VGND.n991 585
R385 VGND.n989 VGND.n987 585
R386 VGND.n1009 VGND.n986 585
R387 VGND.n1010 VGND.n984 585
R388 VGND.n983 VGND.n453 585
R389 VGND.n1015 VGND.n451 585
R390 VGND.n1015 VGND.n1014 585
R391 VGND.n1012 VGND.n453 585
R392 VGND.n1011 VGND.n1010 585
R393 VGND.n1009 VGND.n1008 585
R394 VGND.n1007 VGND.n987 585
R395 VGND.n1005 VGND.n1004 585
R396 VGND.n1003 VGND.n988 585
R397 VGND.n1002 VGND.n1001 585
R398 VGND.n999 VGND.n997 585
R399 VGND.n356 VGND.n355 585
R400 VGND.n1111 VGND.n1110 585
R401 VGND.n1113 VGND.n354 585
R402 VGND.n1018 VGND.n1017 585
R403 VGND.n1018 VGND.n36 585
R404 VGND.n1019 VGND.n450 585
R405 VGND.n1020 VGND.n1019 585
R406 VGND.n1023 VGND.n1022 585
R407 VGND.n1022 VGND.n1021 585
R408 VGND.n1024 VGND.n449 585
R409 VGND.n449 VGND.n448 585
R410 VGND.n1026 VGND.n1025 585
R411 VGND.n1027 VGND.n1026 585
R412 VGND.n447 VGND.n446 585
R413 VGND.n1028 VGND.n447 585
R414 VGND.n1031 VGND.n1030 585
R415 VGND.n1030 VGND.n1029 585
R416 VGND.n1032 VGND.n445 585
R417 VGND.n445 VGND.n444 585
R418 VGND.n1034 VGND.n1033 585
R419 VGND.n1035 VGND.n1034 585
R420 VGND.n442 VGND.n441 585
R421 VGND.n1036 VGND.n442 585
R422 VGND.n1039 VGND.n1038 585
R423 VGND.n1038 VGND.n1037 585
R424 VGND.n1040 VGND.n440 585
R425 VGND.n443 VGND.n440 585
R426 VGND.n565 VGND.n564 585
R427 VGND.n566 VGND.n565 585
R428 VGND.n466 VGND.n465 585
R429 VGND.n567 VGND.n466 585
R430 VGND.n570 VGND.n569 585
R431 VGND.n569 VGND.n568 585
R432 VGND.n571 VGND.n463 585
R433 VGND.n463 VGND.n462 585
R434 VGND.n573 VGND.n572 585
R435 VGND.n574 VGND.n573 585
R436 VGND.n464 VGND.n460 585
R437 VGND.n575 VGND.n460 585
R438 VGND.n972 VGND.n971 585
R439 VGND.n971 VGND.n970 585
R440 VGND.n973 VGND.n457 585
R441 VGND.n457 VGND.n456 585
R442 VGND.n975 VGND.n974 585
R443 VGND.n976 VGND.n975 585
R444 VGND.n458 VGND.n454 585
R445 VGND.n977 VGND.n454 585
R446 VGND.n979 VGND.n455 585
R447 VGND.n979 VGND.n978 585
R448 VGND.n980 VGND.n452 585
R449 VGND.n980 VGND.n35 585
R450 VGND.n495 VGND.n482 585
R451 VGND.n482 VGND.n481 585
R452 VGND.n497 VGND.n496 585
R453 VGND.n498 VGND.n497 585
R454 VGND.n480 VGND.n479 585
R455 VGND.n499 VGND.n480 585
R456 VGND.n502 VGND.n501 585
R457 VGND.n501 VGND.n500 585
R458 VGND.n503 VGND.n478 585
R459 VGND.n478 VGND.n477 585
R460 VGND.n505 VGND.n504 585
R461 VGND.n506 VGND.n505 585
R462 VGND.n476 VGND.n475 585
R463 VGND.n507 VGND.n476 585
R464 VGND.n510 VGND.n509 585
R465 VGND.n509 VGND.n508 585
R466 VGND.n511 VGND.n473 585
R467 VGND.n473 VGND.n472 585
R468 VGND.n513 VGND.n512 585
R469 VGND.n514 VGND.n513 585
R470 VGND.n474 VGND.n471 585
R471 VGND.n515 VGND.n471 585
R472 VGND.n517 VGND.n469 585
R473 VGND.n517 VGND.n516 585
R474 VGND.n577 VGND.n576 585
R475 VGND.n969 VGND.n968 585
R476 VGND.t193 VGND.n969 585
R477 VGND.n2250 VGND.n2249 585
R478 VGND.n2253 VGND.n1697 585
R479 VGND.n1697 VGND.n1696 585
R480 VGND.n2255 VGND.n2254 585
R481 VGND.n2256 VGND.n2255 585
R482 VGND.n1698 VGND.n1694 585
R483 VGND.n2257 VGND.n1694 585
R484 VGND.n2259 VGND.n1695 585
R485 VGND.n2259 VGND.n2258 585
R486 VGND.n2260 VGND.n1693 585
R487 VGND.n2260 VGND.n41 585
R488 VGND.n2262 VGND.n2261 585
R489 VGND.n2261 VGND.n40 585
R490 VGND.n2263 VGND.n1691 585
R491 VGND.n1691 VGND.n1690 585
R492 VGND.n2265 VGND.n2264 585
R493 VGND.n2266 VGND.n2265 585
R494 VGND.n1692 VGND.n1688 585
R495 VGND.n2267 VGND.n1688 585
R496 VGND.n2269 VGND.n1689 585
R497 VGND.n2269 VGND.n2268 585
R498 VGND.n2270 VGND.n1686 585
R499 VGND.n2270 VGND.n46 585
R500 VGND.n2248 VGND.n2247 585
R501 VGND.n1173 VGND.n1172 585
R502 VGND.n1592 VGND.n1591 585
R503 VGND.n1593 VGND.n1592 585
R504 VGND.n1170 VGND.n1169 585
R505 VGND.n1594 VGND.n1170 585
R506 VGND.n1597 VGND.n1596 585
R507 VGND.n1596 VGND.n1595 585
R508 VGND.n1598 VGND.n1168 585
R509 VGND.n1171 VGND.n1168 585
R510 VGND.n1600 VGND.n1599 585
R511 VGND.n1600 VGND.n48 585
R512 VGND.n1601 VGND.n1167 585
R513 VGND.n1601 VGND.n49 585
R514 VGND.n1604 VGND.n1603 585
R515 VGND.n1603 VGND.n1602 585
R516 VGND.n1605 VGND.n1165 585
R517 VGND.n1165 VGND.n1164 585
R518 VGND.n1607 VGND.n1606 585
R519 VGND.n1608 VGND.n1607 585
R520 VGND.n1166 VGND.n1163 585
R521 VGND.n1609 VGND.n1163 585
R522 VGND.n1611 VGND.n1162 585
R523 VGND.n1611 VGND.n1610 585
R524 VGND.n1588 VGND.n45 585
R525 VGND.n2350 VGND.n2349 585
R526 VGND.n2346 VGND.n19 585
R527 VGND.n19 VGND.n17 585
R528 VGND.n2345 VGND.n2344 585
R529 VGND.n2344 VGND.n2343 585
R530 VGND.n23 VGND.n22 585
R531 VGND.n2342 VGND.n23 585
R532 VGND.n2340 VGND.n2339 585
R533 VGND.n2341 VGND.n2340 585
R534 VGND.n2338 VGND.n25 585
R535 VGND.n25 VGND.n24 585
R536 VGND.n2337 VGND.n2336 585
R537 VGND.n2336 VGND.n2335 585
R538 VGND.n27 VGND.n26 585
R539 VGND.n28 VGND.n27 585
R540 VGND.n487 VGND.n486 585
R541 VGND.n486 VGND.n485 585
R542 VGND.n489 VGND.n488 585
R543 VGND.n490 VGND.n489 585
R544 VGND.n484 VGND.n483 585
R545 VGND.n491 VGND.n484 585
R546 VGND.n494 VGND.n493 585
R547 VGND.n493 VGND.n492 585
R548 VGND.n20 VGND.n18 585
R549 VGND.n621 VGND.n620 585
R550 VGND.n620 VGND.n619 585
R551 VGND.n608 VGND.n605 585
R552 VGND.n609 VGND.n608 585
R553 VGND.n607 VGND.n606 585
R554 VGND.n607 VGND.n584 585
R555 VGND.n618 VGND.n617 585
R556 VGND.n619 VGND.n618 585
R557 VGND.n616 VGND.n610 585
R558 VGND.n610 VGND.n609 585
R559 VGND.n613 VGND.n612 585
R560 VGND.n612 VGND.n584 585
R561 VGND.n641 VGND.n639 585
R562 VGND.n654 VGND.n639 585
R563 VGND.n652 VGND.n651 585
R564 VGND.n653 VGND.n652 585
R565 VGND.n642 VGND.n640 585
R566 VGND.n640 VGND.t58 585
R567 VGND.n645 VGND.n587 585
R568 VGND.n661 VGND.n587 585
R569 VGND.n647 VGND.n646 585
R570 VGND.n646 VGND.n588 585
R571 VGND.n656 VGND.n655 585
R572 VGND.n655 VGND.n654 585
R573 VGND.n638 VGND.n637 585
R574 VGND.n653 VGND.n638 585
R575 VGND.n593 VGND.n589 585
R576 VGND.n589 VGND.t58 585
R577 VGND.n660 VGND.n659 585
R578 VGND.n661 VGND.n660 585
R579 VGND.n592 VGND.n590 585
R580 VGND.n590 VGND.n588 585
R581 VGND.n2144 VGND.n2143 585
R582 VGND.n2143 VGND.n42 585
R583 VGND.n2099 VGND.n2098 585
R584 VGND.n2100 VGND.n1900 585
R585 VGND.n2110 VGND.n2109 585
R586 VGND.n2112 VGND.n1899 585
R587 VGND.n2115 VGND.n2114 585
R588 VGND.n2116 VGND.n1895 585
R589 VGND.n2125 VGND.n2124 585
R590 VGND.n2127 VGND.n1894 585
R591 VGND.n2130 VGND.n2129 585
R592 VGND.n2131 VGND.n1888 585
R593 VGND.n2140 VGND.n2139 585
R594 VGND.n2142 VGND.n1887 585
R595 VGND.n2192 VGND.n1777 585
R596 VGND.n2192 VGND.n42 585
R597 VGND.n2145 VGND.n2144 585
R598 VGND.n2145 VGND.n42 585
R599 VGND.n2148 VGND.n2147 585
R600 VGND.n2149 VGND.n1821 585
R601 VGND.n2159 VGND.n2158 585
R602 VGND.n2161 VGND.n1820 585
R603 VGND.n2164 VGND.n2163 585
R604 VGND.n2165 VGND.n1816 585
R605 VGND.n2174 VGND.n2173 585
R606 VGND.n2176 VGND.n1815 585
R607 VGND.n2179 VGND.n2178 585
R608 VGND.n2180 VGND.n1809 585
R609 VGND.n2189 VGND.n2188 585
R610 VGND.n2191 VGND.n1808 585
R611 VGND.n2200 VGND.n1777 585
R612 VGND.n2200 VGND.n42 585
R613 VGND.n2203 VGND.n2202 585
R614 VGND.n2204 VGND.n1713 585
R615 VGND.n2214 VGND.n2213 585
R616 VGND.n2216 VGND.n1712 585
R617 VGND.n2219 VGND.n2218 585
R618 VGND.n2220 VGND.n1708 585
R619 VGND.n2229 VGND.n2228 585
R620 VGND.n2231 VGND.n1707 585
R621 VGND.n2234 VGND.n2233 585
R622 VGND.n2235 VGND.n1701 585
R623 VGND.n2244 VGND.n2243 585
R624 VGND.n2246 VGND.n1699 585
R625 VGND.n838 VGND.n837 585
R626 VGND.n837 VGND.n760 585
R627 VGND.n832 VGND.n762 585
R628 VGND.n834 VGND.n761 585
R629 VGND.n842 VGND.n761 585
R630 VGND.n2074 VGND.n2073 585
R631 VGND.n2075 VGND.n1968 585
R632 VGND.n2077 VGND.n2076 585
R633 VGND.n2079 VGND.n1967 585
R634 VGND.n2082 VGND.n2081 585
R635 VGND.n2083 VGND.n1966 585
R636 VGND.n2085 VGND.n2084 585
R637 VGND.n2087 VGND.n1965 585
R638 VGND.n2090 VGND.n2089 585
R639 VGND.n2091 VGND.n1964 585
R640 VGND.n2093 VGND.n2092 585
R641 VGND.n2093 VGND.n43 585
R642 VGND.n2094 VGND.n1963 585
R643 VGND.n2096 VGND.n1963 585
R644 VGND.n1329 VGND.n1328 585
R645 VGND.n1331 VGND.n1307 585
R646 VGND.n1334 VGND.n1333 585
R647 VGND.n1335 VGND.n1306 585
R648 VGND.n1337 VGND.n1336 585
R649 VGND.n1339 VGND.n1305 585
R650 VGND.n1342 VGND.n1341 585
R651 VGND.n1343 VGND.n1304 585
R652 VGND.n1345 VGND.n1344 585
R653 VGND.n1347 VGND.n1303 585
R654 VGND.n1348 VGND.n1302 585
R655 VGND.n1301 VGND.n43 585
R656 VGND.n1042 VGND.n1041 585
R657 VGND.n1044 VGND.n439 585
R658 VGND.n1045 VGND.n438 585
R659 VGND.n1045 VGND.n43 585
R660 VGND.n1048 VGND.n1047 585
R661 VGND.n1049 VGND.n437 585
R662 VGND.n1051 VGND.n1050 585
R663 VGND.n1053 VGND.n436 585
R664 VGND.n1056 VGND.n1055 585
R665 VGND.n1057 VGND.n435 585
R666 VGND.n1059 VGND.n1058 585
R667 VGND.n1061 VGND.n434 585
R668 VGND.n1062 VGND.n433 585
R669 VGND.n1064 VGND.n433 585
R670 VGND.n891 VGND.t302 575.92
R671 VGND.n875 VGND.t304 575.92
R672 VGND.n878 VGND.t305 575.92
R673 VGND.n678 VGND.t301 572.105
R674 VGND.n895 VGND.n873 560
R675 VGND.t12 VGND.t272 512.451
R676 VGND.n732 VGND.t19 503.615
R677 VGND.n693 VGND.t55 501.755
R678 VGND.n695 VGND.t63 501.755
R679 VGND.t268 VGND.t29 499.685
R680 VGND.t85 VGND.t67 485.805
R681 VGND.t35 VGND.t131 471.925
R682 VGND.t182 VGND.t162 471.825
R683 VGND.t181 VGND.t88 462.974
R684 VGND.t153 VGND.t34 458.045
R685 VGND.t141 VGND.t21 458.045
R686 VGND.t245 VGND.t77 458.045
R687 VGND.t278 VGND.t104 458.045
R688 VGND.t120 VGND.t177 458.045
R689 VGND.t25 VGND.t65 458.045
R690 VGND.n883 VGND.n873 441.601
R691 VGND.n948 VGND.t29 437.224
R692 VGND.t262 VGND.n583 426.358
R693 VGND.n737 VGND.t243 415.262
R694 VGND.n733 VGND.t137 415.262
R695 VGND.n685 VGND.n684 385.658
R696 VGND.t41 VGND.n898 381.704
R697 VGND.n467 VGND.n30 370.214
R698 VGND.n467 VGND.n29 365.957
R699 VGND.n960 VGND.t33 364.351
R700 VGND.t63 VGND.n693 347.368
R701 VGND.t287 VGND.n695 347.368
R702 VGND.n696 VGND.t53 347.368
R703 VGND.t49 VGND.n707 347.368
R704 VGND.n709 VGND.t114 347.368
R705 VGND.t121 VGND.t268 347.003
R706 VGND.t100 VGND.t102 347.003
R707 VGND.t190 VGND.t11 347.003
R708 VGND.n730 VGND.t51 344.579
R709 VGND.n725 VGND.t113 344.579
R710 VGND.t156 VGND.n443 338.411
R711 VGND.n808 VGND.t215 336.329
R712 VGND.n808 VGND.t200 336.329
R713 VGND.n788 VGND.t196 336.329
R714 VGND.n788 VGND.t219 336.329
R715 VGND.n830 VGND.t204 330
R716 VGND.n763 VGND.t232 330
R717 VGND.t92 VGND.t151 329.716
R718 VGND.t193 VGND.n29 327.661
R719 VGND.t193 VGND.n31 172.876
R720 VGND.t193 VGND.n33 172.876
R721 VGND.t193 VGND.n30 323.404
R722 VGND.t193 VGND.n32 172.615
R723 VGND.t193 VGND.n34 172.615
R724 VGND.t58 VGND.t88 317.781
R725 VGND.n952 VGND.t33 317.774
R726 VGND.t298 VGND.n909 312.303
R727 VGND.n910 VGND.t133 312.303
R728 VGND.t96 VGND.n923 312.303
R729 VGND.n935 VGND.t36 309.733
R730 VGND.n932 VGND.t30 309.733
R731 VGND.n931 VGND.t269 309.733
R732 VGND.n757 VGND.t211 304.634
R733 VGND.n855 VGND.t240 304.634
R734 VGND.n770 VGND.t236 304.634
R735 VGND.n865 VGND.t228 304.634
R736 VGND.n1700 VGND.t181 296.538
R737 VGND.n861 VGND.t208 292.584
R738 VGND.n848 VGND.t223 292.584
R739 VGND.n874 VGND.n872 292.5
R740 VGND.n880 VGND.n872 292.5
R741 VGND.n873 VGND.n871 292.5
R742 VGND.n880 VGND.n871 292.5
R743 VGND.n684 VGND.t123 289.243
R744 VGND.t53 VGND.t260 283.041
R745 VGND.t171 VGND.t270 283.041
R746 VGND.t293 VGND.t49 283.041
R747 VGND.t114 VGND.t89 283.041
R748 VGND.n2248 VGND.t88 280.567
R749 VGND.n898 VGND.n897 278.938
R750 VGND.t272 VGND.n737 273.897
R751 VGND.n733 VGND.t243 273.897
R752 VGND.t137 VGND.n732 273.897
R753 VGND.n909 VGND.t256 270.663
R754 VGND.n910 VGND.t276 270.663
R755 VGND.n923 VGND.t5 270.663
R756 VGND.n924 VGND.t291 270.663
R757 VGND.n1063 VGND.n43 264.301
R758 VGND.n2252 VGND.n2251 264.301
R759 VGND.n1590 VGND.n1589 264.301
R760 VGND.n2348 VGND.n2347 264.301
R761 VGND.n2095 VGND.n43 264.301
R762 VGND.n1351 VGND.n1350 264.301
R763 VGND.n4 VGND.n3 261.733
R764 VGND.n934 VGND.n933 261.733
R765 VGND.n937 VGND.n936 261.733
R766 VGND.n939 VGND.n938 261.733
R767 VGND.n941 VGND.n940 261.733
R768 VGND.n943 VGND.n942 261.733
R769 VGND.n945 VGND.n944 261.733
R770 VGND.n930 VGND.n929 261.733
R771 VGND.n928 VGND.n927 261.733
R772 VGND.n664 VGND.n663 261.733
R773 VGND.n919 VGND.n918 261.733
R774 VGND.n921 VGND.n920 260.514
R775 VGND.n957 VGND.t280 260
R776 VGND.t280 VGND.n579 260
R777 VGND.n1018 VGND.n451 259.416
R778 VGND.n2051 VGND.n2050 259.416
R779 VGND.n2299 VGND.n2298 259.416
R780 VGND.n493 VGND.n482 259.416
R781 VGND.n565 VGND.n468 259.416
R782 VGND.n1612 VGND.n1611 259.416
R783 VGND.n1639 VGND.n122 259.416
R784 VGND.n2332 VGND.n73 259.416
R785 VGND.n2271 VGND.n2270 259.416
R786 VGND.n1948 VGND.n1906 258.334
R787 VGND.n1869 VGND.n1827 258.334
R788 VGND.n336 VGND.n334 258.334
R789 VGND.n416 VGND.n415 258.334
R790 VGND.n1530 VGND.n1488 258.334
R791 VGND.n1262 VGND.n1205 258.334
R792 VGND.n1434 VGND.n1375 258.334
R793 VGND.n1761 VGND.n1719 258.334
R794 VGND.n240 VGND.n239 258.334
R795 VGND.t193 VGND.n461 257.779
R796 VGND.n676 VGND.t92 255.815
R797 VGND.n1687 VGND.n44 254.34
R798 VGND.n2276 VGND.n44 254.34
R799 VGND.n1684 VGND.n44 254.34
R800 VGND.n2283 VGND.n44 254.34
R801 VGND.n1681 VGND.n44 254.34
R802 VGND.n2290 VGND.n44 254.34
R803 VGND.n1468 VGND.n1467 254.34
R804 VGND.n1468 VGND.n1299 254.34
R805 VGND.n1468 VGND.n1298 254.34
R806 VGND.n1468 VGND.n1297 254.34
R807 VGND.n1468 VGND.n1296 254.34
R808 VGND.n1468 VGND.n1295 254.34
R809 VGND.n1468 VGND.n1294 254.34
R810 VGND.n1468 VGND.n1180 254.34
R811 VGND.n1468 VGND.n1179 254.34
R812 VGND.n1468 VGND.n1178 254.34
R813 VGND.n1468 VGND.n1177 254.34
R814 VGND.n1468 VGND.n1176 254.34
R815 VGND.n1481 VGND.n1468 254.34
R816 VGND.n1556 VGND.n1468 254.34
R817 VGND.n1558 VGND.n1468 254.34
R818 VGND.n1571 VGND.n1468 254.34
R819 VGND.n1573 VGND.n1468 254.34
R820 VGND.n1586 VGND.n1468 254.34
R821 VGND.n2334 VGND.n2333 254.34
R822 VGND.n2334 VGND.n71 254.34
R823 VGND.n2334 VGND.n70 254.34
R824 VGND.n2334 VGND.n69 254.34
R825 VGND.n2334 VGND.n68 254.34
R826 VGND.n2334 VGND.n67 254.34
R827 VGND.n2334 VGND.n66 254.34
R828 VGND.n2334 VGND.n65 254.34
R829 VGND.n2334 VGND.n64 254.34
R830 VGND.n2334 VGND.n63 254.34
R831 VGND.n2334 VGND.n62 254.34
R832 VGND.n2334 VGND.n61 254.34
R833 VGND.n2334 VGND.n60 254.34
R834 VGND.n2334 VGND.n59 254.34
R835 VGND.n2334 VGND.n58 254.34
R836 VGND.n2334 VGND.n57 254.34
R837 VGND.n2334 VGND.n56 254.34
R838 VGND.n2334 VGND.n55 254.34
R839 VGND.n1156 VGND.n266 254.34
R840 VGND.n1156 VGND.n267 254.34
R841 VGND.n1156 VGND.n268 254.34
R842 VGND.n1156 VGND.n269 254.34
R843 VGND.n1156 VGND.n270 254.34
R844 VGND.n1156 VGND.n271 254.34
R845 VGND.n1156 VGND.n272 254.34
R846 VGND.n1156 VGND.n273 254.34
R847 VGND.n1156 VGND.n274 254.34
R848 VGND.n1156 VGND.n275 254.34
R849 VGND.n1156 VGND.n276 254.34
R850 VGND.n1156 VGND.n1155 254.34
R851 VGND.n1157 VGND.n1156 254.34
R852 VGND.n1156 VGND.n265 254.34
R853 VGND.n1156 VGND.n153 254.34
R854 VGND.n1156 VGND.n152 254.34
R855 VGND.n1156 VGND.n151 254.34
R856 VGND.n1156 VGND.n150 254.34
R857 VGND.n539 VGND.n29 254.34
R858 VGND.n536 VGND.n29 254.34
R859 VGND.n530 VGND.n29 254.34
R860 VGND.n527 VGND.n29 254.34
R861 VGND.n522 VGND.n29 254.34
R862 VGND.n519 VGND.n29 254.34
R863 VGND.n560 VGND.n30 254.34
R864 VGND.n518 VGND.n30 254.34
R865 VGND.n553 VGND.n30 254.34
R866 VGND.n547 VGND.n30 254.34
R867 VGND.n545 VGND.n30 254.34
R868 VGND.n533 VGND.n30 254.34
R869 VGND.n1668 VGND.n52 254.34
R870 VGND.n111 VGND.n52 254.34
R871 VGND.n1656 VGND.n52 254.34
R872 VGND.n1652 VGND.n52 254.34
R873 VGND.n1642 VGND.n52 254.34
R874 VGND.n1640 VGND.n52 254.34
R875 VGND.n1636 VGND.n53 254.34
R876 VGND.n1646 VGND.n53 254.34
R877 VGND.n1648 VGND.n53 254.34
R878 VGND.n1660 VGND.n53 254.34
R879 VGND.n1663 VGND.n53 254.34
R880 VGND.n113 VGND.n53 254.34
R881 VGND.n2194 VGND.n33 254.34
R882 VGND.n1806 VGND.n33 254.34
R883 VGND.n1796 VGND.n33 254.34
R884 VGND.n1794 VGND.n33 254.34
R885 VGND.n1785 VGND.n33 254.34
R886 VGND.n2297 VGND.n33 254.34
R887 VGND.n2293 VGND.n34 254.34
R888 VGND.n1788 VGND.n34 254.34
R889 VGND.n1790 VGND.n34 254.34
R890 VGND.n1800 VGND.n34 254.34
R891 VGND.n1802 VGND.n34 254.34
R892 VGND.n2198 VGND.n34 254.34
R893 VGND.n1675 VGND.n44 254.34
R894 VGND.n2028 VGND.n44 254.34
R895 VGND.n2024 VGND.n44 254.34
R896 VGND.n2035 VGND.n44 254.34
R897 VGND.n2021 VGND.n44 254.34
R898 VGND.n2042 VGND.n44 254.34
R899 VGND.n1978 VGND.n44 254.34
R900 VGND.n2056 VGND.n44 254.34
R901 VGND.n1975 VGND.n44 254.34
R902 VGND.n2063 VGND.n44 254.34
R903 VGND.n1972 VGND.n44 254.34
R904 VGND.n2070 VGND.n44 254.34
R905 VGND.n1996 VGND.n31 254.34
R906 VGND.n1994 VGND.n31 254.34
R907 VGND.n1991 VGND.n31 254.34
R908 VGND.n1986 VGND.n31 254.34
R909 VGND.n1983 VGND.n31 254.34
R910 VGND.n2049 VGND.n31 254.34
R911 VGND.n2045 VGND.n32 254.34
R912 VGND.n2016 VGND.n32 254.34
R913 VGND.n2010 VGND.n32 254.34
R914 VGND.n2008 VGND.n32 254.34
R915 VGND.n2002 VGND.n32 254.34
R916 VGND.n2000 VGND.n32 254.34
R917 VGND.n99 VGND.n50 254.34
R918 VGND.n96 VGND.n50 254.34
R919 VGND.n91 VGND.n50 254.34
R920 VGND.n88 VGND.n50 254.34
R921 VGND.n83 VGND.n50 254.34
R922 VGND.n80 VGND.n50 254.34
R923 VGND.n2327 VGND.n51 254.34
R924 VGND.n79 VGND.n51 254.34
R925 VGND.n2320 VGND.n51 254.34
R926 VGND.n2314 VGND.n51 254.34
R927 VGND.n2312 VGND.n51 254.34
R928 VGND.n2306 VGND.n51 254.34
R929 VGND.n1108 VGND.n39 254.34
R930 VGND.n995 VGND.n39 254.34
R931 VGND.n993 VGND.n39 254.34
R932 VGND.n990 VGND.n39 254.34
R933 VGND.n985 VGND.n39 254.34
R934 VGND.n982 VGND.n39 254.34
R935 VGND.n1013 VGND.n37 254.34
R936 VGND.n981 VGND.n37 254.34
R937 VGND.n1006 VGND.n37 254.34
R938 VGND.n1000 VGND.n37 254.34
R939 VGND.n998 VGND.n37 254.34
R940 VGND.n1112 VGND.n37 254.34
R941 VGND.n2097 VGND.n1700 254.34
R942 VGND.n2111 VGND.n1700 254.34
R943 VGND.n2113 VGND.n1700 254.34
R944 VGND.n2126 VGND.n1700 254.34
R945 VGND.n2128 VGND.n1700 254.34
R946 VGND.n2141 VGND.n1700 254.34
R947 VGND.n2146 VGND.n1700 254.34
R948 VGND.n2160 VGND.n1700 254.34
R949 VGND.n2162 VGND.n1700 254.34
R950 VGND.n2175 VGND.n1700 254.34
R951 VGND.n2177 VGND.n1700 254.34
R952 VGND.n2190 VGND.n1700 254.34
R953 VGND.n2201 VGND.n1700 254.34
R954 VGND.n2215 VGND.n1700 254.34
R955 VGND.n2217 VGND.n1700 254.34
R956 VGND.n2230 VGND.n1700 254.34
R957 VGND.n2232 VGND.n1700 254.34
R958 VGND.n2245 VGND.n1700 254.34
R959 VGND.n2072 VGND.n43 254.34
R960 VGND.n2078 VGND.n43 254.34
R961 VGND.n2080 VGND.n43 254.34
R962 VGND.n2086 VGND.n43 254.34
R963 VGND.n2088 VGND.n43 254.34
R964 VGND.n1330 VGND.n43 254.34
R965 VGND.n1332 VGND.n43 254.34
R966 VGND.n1338 VGND.n43 254.34
R967 VGND.n1340 VGND.n43 254.34
R968 VGND.n1346 VGND.n43 254.34
R969 VGND.n1349 VGND.n43 254.34
R970 VGND.n1043 VGND.n43 254.34
R971 VGND.n1046 VGND.n43 254.34
R972 VGND.n1052 VGND.n43 254.34
R973 VGND.n1054 VGND.n43 254.34
R974 VGND.n1060 VGND.n43 254.34
R975 VGND.t250 VGND.n682 254.184
R976 VGND.t7 VGND.n745 250.349
R977 VGND.t7 VGND.n746 250.349
R978 VGND.n819 VGND.n818 250.349
R979 VGND.n820 VGND.n819 250.349
R980 VGND.n774 VGND.n773 250.349
R981 VGND.n842 VGND.n841 250.349
R982 VGND.n1042 VGND.n440 249.663
R983 VGND.n2073 VGND.n2071 249.663
R984 VGND.n2044 VGND.n2043 249.663
R985 VGND.n561 VGND.n517 249.663
R986 VGND.n1014 VGND.n980 249.663
R987 VGND.n1637 VGND.n1635 249.663
R988 VGND.n2328 VGND.n78 249.663
R989 VGND.n1329 VGND.n1308 249.663
R990 VGND.n2292 VGND.n2291 249.663
R991 VGND.n724 VGND.n722 247.391
R992 VGND.n881 VGND.t169 246.796
R993 VGND.n897 VGND.t94 246.796
R994 VGND.n655 VGND.n638 246.25
R995 VGND.n638 VGND.n589 246.25
R996 VGND.n660 VGND.n589 246.25
R997 VGND.n660 VGND.n590 246.25
R998 VGND.n652 VGND.n639 246.25
R999 VGND.n652 VGND.n640 246.25
R1000 VGND.n640 VGND.n587 246.25
R1001 VGND.n646 VGND.n587 246.25
R1002 VGND.n951 VGND.n584 246.137
R1003 VGND.n758 VGND.t214 245
R1004 VGND.n856 VGND.t242 245
R1005 VGND.n771 VGND.t239 245
R1006 VGND.n866 VGND.t229 245
R1007 VGND.n959 VGND.n958 241.643
R1008 VGND.t19 VGND.n730 238.554
R1009 VGND.n725 VGND.t51 238.554
R1010 VGND.t183 VGND.n724 238.554
R1011 VGND.n722 VGND.t98 238.554
R1012 VGND.n713 VGND.t274 238.554
R1013 VGND.n713 VGND.t296 238.554
R1014 VGND.t116 VGND.n712 238.554
R1015 VGND.n901 VGND.n899 233.793
R1016 VGND.n947 VGND.t282 233
R1017 VGND.n925 VGND.t149 233
R1018 VGND.n917 VGND.n916 232.934
R1019 VGND.n915 VGND.n914 232.934
R1020 VGND.n913 VGND.n912 232.934
R1021 VGND.n666 VGND.n665 232.934
R1022 VGND.n905 VGND.n904 232.934
R1023 VGND.n907 VGND.n906 232.934
R1024 VGND.n903 VGND.n902 232.934
R1025 VGND.n901 VGND.n900 232.934
R1026 VGND.n895 VGND.n894 230.4
R1027 VGND.n884 VGND.n883 230.4
R1028 VGND.t162 VGND.n739 222.036
R1029 VGND.n669 VGND.t180 211.857
R1030 VGND.n670 VGND.t32 211.857
R1031 VGND.n718 VGND.t128 211.857
R1032 VGND.n719 VGND.t2 211.857
R1033 VGND.n702 VGND.t90 211.857
R1034 VGND.n703 VGND.t294 211.857
R1035 VGND.n700 VGND.t172 211.857
R1036 VGND.n699 VGND.t261 211.857
R1037 VGND.n853 VGND.n748 204.201
R1038 VGND.n854 VGND.n747 204.201
R1039 VGND.n750 VGND.n749 204.201
R1040 VGND.n863 VGND.n741 204.201
R1041 VGND.n864 VGND.n740 204.201
R1042 VGND.n743 VGND.n742 204.201
R1043 VGND.n868 VGND.t182 203.532
R1044 VGND.n762 VGND.n761 197
R1045 VGND.n837 VGND.n761 197
R1046 VGND.n618 VGND.n610 197
R1047 VGND.n612 VGND.n610 197
R1048 VGND.n620 VGND.n608 197
R1049 VGND.n608 VGND.n607 197
R1050 VGND.n821 VGND.n812 197
R1051 VGND.n798 VGND.n797 197
R1052 VGND.n769 VGND.n767 197
R1053 VGND.n775 VGND.n768 197
R1054 VGND.n2143 VGND.n2142 197
R1055 VGND.n2192 VGND.n2191 197
R1056 VGND.n277 VGND.n145 197
R1057 VGND.n1106 VGND.n1105 197
R1058 VGND.n1588 VGND.n1587 197
R1059 VGND.n1175 VGND.n105 197
R1060 VGND.n1377 VGND.n104 197
R1061 VGND.n2247 VGND.n2246 197
R1062 VGND.n149 VGND.n20 197
R1063 VGND.t113 VGND.t183 194.379
R1064 VGND.t1 VGND.t98 194.379
R1065 VGND.t274 VGND.t127 194.379
R1066 VGND.t296 VGND.t31 194.379
R1067 VGND.t179 VGND.t116 194.379
R1068 VGND.n688 VGND.n687 192.829
R1069 VGND.n858 VGND.t220 189.57
R1070 VGND.n676 VGND.t262 187.597
R1071 VGND.n681 VGND.t151 187.597
R1072 VGND.n924 VGND.t148 187.382
R1073 VGND.t281 VGND.n948 187.382
R1074 VGND.n2098 VGND.n2096 187.249
R1075 VGND.n2147 VGND.n2145 187.249
R1076 VGND.n1115 VGND.n1114 187.249
R1077 VGND.n1065 VGND.n1064 187.249
R1078 VGND.n2303 VGND.n107 187.249
R1079 VGND.n2305 VGND.n102 187.249
R1080 VGND.n1466 VGND.n1301 187.249
R1081 VGND.n2202 VGND.n2200 187.249
R1082 VGND.n1159 VGND.n1158 187.249
R1083 VGND.n657 VGND.n656 185
R1084 VGND.n635 VGND.n592 185
R1085 VGND.n649 VGND.n641 185
R1086 VGND.n649 VGND.n642 185
R1087 VGND.n643 VGND.n641 185
R1088 VGND.n647 VGND.n643 185
R1089 VGND.n840 VGND.n839 185
R1090 VGND.n839 VGND.n838 185
R1091 VGND.n817 VGND.n816 185
R1092 VGND.n816 VGND.n809 185
R1093 VGND.n793 VGND.n792 185
R1094 VGND.n792 VGND.n789 185
R1095 VGND.n781 VGND.n780 185
R1096 VGND.n781 VGND.n765 185
R1097 VGND.n1948 VGND.n1947 185
R1098 VGND.n1950 VGND.n1905 185
R1099 VGND.n1953 VGND.n1952 185
R1100 VGND.n1954 VGND.n1904 185
R1101 VGND.n1956 VGND.n1955 185
R1102 VGND.n1958 VGND.n1903 185
R1103 VGND.n1961 VGND.n1960 185
R1104 VGND.n1962 VGND.n1902 185
R1105 VGND.n2103 VGND.n2102 185
R1106 VGND.n1930 VGND.n1910 185
R1107 VGND.n1932 VGND.n1931 185
R1108 VGND.n1934 VGND.n1909 185
R1109 VGND.n1937 VGND.n1936 185
R1110 VGND.n1938 VGND.n1908 185
R1111 VGND.n1940 VGND.n1939 185
R1112 VGND.n1942 VGND.n1907 185
R1113 VGND.n1945 VGND.n1944 185
R1114 VGND.n1946 VGND.n1906 185
R1115 VGND.n2137 VGND.n2136 185
R1116 VGND.n1915 VGND.n1890 185
R1117 VGND.n1917 VGND.n1916 185
R1118 VGND.n1919 VGND.n1913 185
R1119 VGND.n1921 VGND.n1920 185
R1120 VGND.n1922 VGND.n1912 185
R1121 VGND.n1924 VGND.n1923 185
R1122 VGND.n1926 VGND.n1911 185
R1123 VGND.n1929 VGND.n1928 185
R1124 VGND.n2135 VGND.n1889 185
R1125 VGND.n2133 VGND.n2132 185
R1126 VGND.n1893 VGND.n1892 185
R1127 VGND.n2123 VGND.n2122 185
R1128 VGND.n2120 VGND.n1896 185
R1129 VGND.n2118 VGND.n2117 185
R1130 VGND.n1898 VGND.n1897 185
R1131 VGND.n2108 VGND.n2107 185
R1132 VGND.n2105 VGND.n1901 185
R1133 VGND.n1869 VGND.n1868 185
R1134 VGND.n1871 VGND.n1826 185
R1135 VGND.n1874 VGND.n1873 185
R1136 VGND.n1875 VGND.n1825 185
R1137 VGND.n1877 VGND.n1876 185
R1138 VGND.n1879 VGND.n1824 185
R1139 VGND.n1882 VGND.n1881 185
R1140 VGND.n1883 VGND.n1823 185
R1141 VGND.n2152 VGND.n2151 185
R1142 VGND.n1851 VGND.n1831 185
R1143 VGND.n1853 VGND.n1852 185
R1144 VGND.n1855 VGND.n1830 185
R1145 VGND.n1858 VGND.n1857 185
R1146 VGND.n1859 VGND.n1829 185
R1147 VGND.n1861 VGND.n1860 185
R1148 VGND.n1863 VGND.n1828 185
R1149 VGND.n1866 VGND.n1865 185
R1150 VGND.n1867 VGND.n1827 185
R1151 VGND.n2186 VGND.n2185 185
R1152 VGND.n1836 VGND.n1811 185
R1153 VGND.n1838 VGND.n1837 185
R1154 VGND.n1840 VGND.n1834 185
R1155 VGND.n1842 VGND.n1841 185
R1156 VGND.n1843 VGND.n1833 185
R1157 VGND.n1845 VGND.n1844 185
R1158 VGND.n1847 VGND.n1832 185
R1159 VGND.n1850 VGND.n1849 185
R1160 VGND.n2184 VGND.n1810 185
R1161 VGND.n2182 VGND.n2181 185
R1162 VGND.n1814 VGND.n1813 185
R1163 VGND.n2172 VGND.n2171 185
R1164 VGND.n2169 VGND.n1817 185
R1165 VGND.n2167 VGND.n2166 185
R1166 VGND.n1819 VGND.n1818 185
R1167 VGND.n2157 VGND.n2156 185
R1168 VGND.n2154 VGND.n1822 185
R1169 VGND.n337 VGND.n336 185
R1170 VGND.n338 VGND.n293 185
R1171 VGND.n340 VGND.n339 185
R1172 VGND.n342 VGND.n292 185
R1173 VGND.n345 VGND.n344 185
R1174 VGND.n346 VGND.n291 185
R1175 VGND.n348 VGND.n347 185
R1176 VGND.n350 VGND.n290 185
R1177 VGND.n352 VGND.n351 185
R1178 VGND.n318 VGND.n298 185
R1179 VGND.n321 VGND.n320 185
R1180 VGND.n322 VGND.n297 185
R1181 VGND.n324 VGND.n323 185
R1182 VGND.n326 VGND.n296 185
R1183 VGND.n329 VGND.n328 185
R1184 VGND.n330 VGND.n295 185
R1185 VGND.n332 VGND.n331 185
R1186 VGND.n334 VGND.n294 185
R1187 VGND.n1150 VGND.n1149 185
R1188 VGND.n304 VGND.n280 185
R1189 VGND.n306 VGND.n305 185
R1190 VGND.n307 VGND.n302 185
R1191 VGND.n309 VGND.n308 185
R1192 VGND.n311 VGND.n300 185
R1193 VGND.n313 VGND.n312 185
R1194 VGND.n314 VGND.n299 185
R1195 VGND.n316 VGND.n315 185
R1196 VGND.n1148 VGND.n279 185
R1197 VGND.n1146 VGND.n1145 185
R1198 VGND.n283 VGND.n282 185
R1199 VGND.n1139 VGND.n1138 185
R1200 VGND.n1136 VGND.n285 185
R1201 VGND.n1134 VGND.n1133 185
R1202 VGND.n287 VGND.n286 185
R1203 VGND.n1125 VGND.n1124 185
R1204 VGND.n1122 VGND.n1121 185
R1205 VGND.n417 VGND.n416 185
R1206 VGND.n419 VGND.n418 185
R1207 VGND.n421 VGND.n420 185
R1208 VGND.n423 VGND.n422 185
R1209 VGND.n425 VGND.n424 185
R1210 VGND.n427 VGND.n426 185
R1211 VGND.n429 VGND.n428 185
R1212 VGND.n431 VGND.n430 185
R1213 VGND.n432 VGND.n380 185
R1214 VGND.n399 VGND.n398 185
R1215 VGND.n401 VGND.n400 185
R1216 VGND.n403 VGND.n402 185
R1217 VGND.n405 VGND.n404 185
R1218 VGND.n407 VGND.n406 185
R1219 VGND.n409 VGND.n408 185
R1220 VGND.n411 VGND.n410 185
R1221 VGND.n413 VGND.n412 185
R1222 VGND.n415 VGND.n414 185
R1223 VGND.n372 VGND.n358 185
R1224 VGND.n383 VGND.n382 185
R1225 VGND.n385 VGND.n384 185
R1226 VGND.n387 VGND.n386 185
R1227 VGND.n389 VGND.n388 185
R1228 VGND.n391 VGND.n390 185
R1229 VGND.n393 VGND.n392 185
R1230 VGND.n395 VGND.n394 185
R1231 VGND.n397 VGND.n396 185
R1232 VGND.n362 VGND.n359 185
R1233 VGND.n1098 VGND.n1097 185
R1234 VGND.n1071 VGND.n361 185
R1235 VGND.n1077 VGND.n1076 185
R1236 VGND.n1075 VGND.n1070 185
R1237 VGND.n1084 VGND.n1083 185
R1238 VGND.n1082 VGND.n1069 185
R1239 VGND.n1089 VGND.n381 185
R1240 VGND.n1094 VGND.n1093 185
R1241 VGND.n1530 VGND.n1529 185
R1242 VGND.n1532 VGND.n1487 185
R1243 VGND.n1535 VGND.n1534 185
R1244 VGND.n1536 VGND.n1486 185
R1245 VGND.n1538 VGND.n1537 185
R1246 VGND.n1540 VGND.n1485 185
R1247 VGND.n1543 VGND.n1542 185
R1248 VGND.n1544 VGND.n1484 185
R1249 VGND.n1548 VGND.n1547 185
R1250 VGND.n1512 VGND.n1492 185
R1251 VGND.n1514 VGND.n1513 185
R1252 VGND.n1516 VGND.n1491 185
R1253 VGND.n1519 VGND.n1518 185
R1254 VGND.n1520 VGND.n1490 185
R1255 VGND.n1522 VGND.n1521 185
R1256 VGND.n1524 VGND.n1489 185
R1257 VGND.n1527 VGND.n1526 185
R1258 VGND.n1528 VGND.n1488 185
R1259 VGND.n1582 VGND.n1581 185
R1260 VGND.n1497 VGND.n1471 185
R1261 VGND.n1499 VGND.n1498 185
R1262 VGND.n1501 VGND.n1495 185
R1263 VGND.n1503 VGND.n1502 185
R1264 VGND.n1504 VGND.n1494 185
R1265 VGND.n1506 VGND.n1505 185
R1266 VGND.n1508 VGND.n1493 185
R1267 VGND.n1511 VGND.n1510 185
R1268 VGND.n1580 VGND.n1470 185
R1269 VGND.n1578 VGND.n1577 185
R1270 VGND.n1474 VGND.n1473 185
R1271 VGND.n1568 VGND.n1567 185
R1272 VGND.n1565 VGND.n1477 185
R1273 VGND.n1563 VGND.n1562 185
R1274 VGND.n1479 VGND.n1478 185
R1275 VGND.n1553 VGND.n1552 185
R1276 VGND.n1550 VGND.n1483 185
R1277 VGND.n1264 VGND.n1205 185
R1278 VGND.n1279 VGND.n1278 185
R1279 VGND.n1277 VGND.n1206 185
R1280 VGND.n1276 VGND.n1275 185
R1281 VGND.n1274 VGND.n1273 185
R1282 VGND.n1272 VGND.n1271 185
R1283 VGND.n1270 VGND.n1269 185
R1284 VGND.n1268 VGND.n1267 185
R1285 VGND.n1266 VGND.n1265 185
R1286 VGND.n1247 VGND.n1246 185
R1287 VGND.n1249 VGND.n1248 185
R1288 VGND.n1251 VGND.n1250 185
R1289 VGND.n1253 VGND.n1252 185
R1290 VGND.n1255 VGND.n1254 185
R1291 VGND.n1257 VGND.n1256 185
R1292 VGND.n1259 VGND.n1258 185
R1293 VGND.n1261 VGND.n1260 185
R1294 VGND.n1263 VGND.n1262 185
R1295 VGND.n1229 VGND.n1228 185
R1296 VGND.n1231 VGND.n1230 185
R1297 VGND.n1233 VGND.n1232 185
R1298 VGND.n1235 VGND.n1234 185
R1299 VGND.n1237 VGND.n1236 185
R1300 VGND.n1239 VGND.n1238 185
R1301 VGND.n1241 VGND.n1240 185
R1302 VGND.n1243 VGND.n1242 185
R1303 VGND.n1245 VGND.n1244 185
R1304 VGND.n1227 VGND.n1226 185
R1305 VGND.n1221 VGND.n1220 185
R1306 VGND.n1219 VGND.n1218 185
R1307 VGND.n1214 VGND.n1213 185
R1308 VGND.n1209 VGND.n1190 185
R1309 VGND.n1283 VGND.n1282 185
R1310 VGND.n1189 VGND.n1187 185
R1311 VGND.n1289 VGND.n1288 185
R1312 VGND.n1291 VGND.n1290 185
R1313 VGND.n1436 VGND.n1375 185
R1314 VGND.n1450 VGND.n1449 185
R1315 VGND.n1448 VGND.n1376 185
R1316 VGND.n1447 VGND.n1446 185
R1317 VGND.n1445 VGND.n1444 185
R1318 VGND.n1443 VGND.n1442 185
R1319 VGND.n1441 VGND.n1440 185
R1320 VGND.n1439 VGND.n1438 185
R1321 VGND.n1437 VGND.n1352 185
R1322 VGND.n1419 VGND.n1418 185
R1323 VGND.n1421 VGND.n1420 185
R1324 VGND.n1423 VGND.n1422 185
R1325 VGND.n1425 VGND.n1424 185
R1326 VGND.n1427 VGND.n1426 185
R1327 VGND.n1429 VGND.n1428 185
R1328 VGND.n1431 VGND.n1430 185
R1329 VGND.n1433 VGND.n1432 185
R1330 VGND.n1435 VGND.n1434 185
R1331 VGND.n1401 VGND.n1400 185
R1332 VGND.n1403 VGND.n1402 185
R1333 VGND.n1405 VGND.n1404 185
R1334 VGND.n1407 VGND.n1406 185
R1335 VGND.n1409 VGND.n1408 185
R1336 VGND.n1411 VGND.n1410 185
R1337 VGND.n1413 VGND.n1412 185
R1338 VGND.n1415 VGND.n1414 185
R1339 VGND.n1417 VGND.n1416 185
R1340 VGND.n1399 VGND.n1398 185
R1341 VGND.n1393 VGND.n1392 185
R1342 VGND.n1391 VGND.n1390 185
R1343 VGND.n1386 VGND.n1385 185
R1344 VGND.n1381 VGND.n1360 185
R1345 VGND.n1454 VGND.n1453 185
R1346 VGND.n1359 VGND.n1357 185
R1347 VGND.n1460 VGND.n1459 185
R1348 VGND.n1462 VGND.n1461 185
R1349 VGND.n1761 VGND.n1760 185
R1350 VGND.n1763 VGND.n1718 185
R1351 VGND.n1766 VGND.n1765 185
R1352 VGND.n1767 VGND.n1717 185
R1353 VGND.n1769 VGND.n1768 185
R1354 VGND.n1771 VGND.n1716 185
R1355 VGND.n1774 VGND.n1773 185
R1356 VGND.n1775 VGND.n1715 185
R1357 VGND.n2207 VGND.n2206 185
R1358 VGND.n1743 VGND.n1723 185
R1359 VGND.n1745 VGND.n1744 185
R1360 VGND.n1747 VGND.n1722 185
R1361 VGND.n1750 VGND.n1749 185
R1362 VGND.n1751 VGND.n1721 185
R1363 VGND.n1753 VGND.n1752 185
R1364 VGND.n1755 VGND.n1720 185
R1365 VGND.n1758 VGND.n1757 185
R1366 VGND.n1759 VGND.n1719 185
R1367 VGND.n2241 VGND.n2240 185
R1368 VGND.n1728 VGND.n1703 185
R1369 VGND.n1730 VGND.n1729 185
R1370 VGND.n1732 VGND.n1726 185
R1371 VGND.n1734 VGND.n1733 185
R1372 VGND.n1735 VGND.n1725 185
R1373 VGND.n1737 VGND.n1736 185
R1374 VGND.n1739 VGND.n1724 185
R1375 VGND.n1742 VGND.n1741 185
R1376 VGND.n2239 VGND.n1702 185
R1377 VGND.n2237 VGND.n2236 185
R1378 VGND.n1706 VGND.n1705 185
R1379 VGND.n2227 VGND.n2226 185
R1380 VGND.n2224 VGND.n1709 185
R1381 VGND.n2222 VGND.n2221 185
R1382 VGND.n1711 VGND.n1710 185
R1383 VGND.n2212 VGND.n2211 185
R1384 VGND.n2209 VGND.n1714 185
R1385 VGND.n241 VGND.n240 185
R1386 VGND.n243 VGND.n242 185
R1387 VGND.n245 VGND.n244 185
R1388 VGND.n247 VGND.n246 185
R1389 VGND.n249 VGND.n248 185
R1390 VGND.n251 VGND.n250 185
R1391 VGND.n253 VGND.n252 185
R1392 VGND.n254 VGND.n175 185
R1393 VGND.n258 VGND.n257 185
R1394 VGND.n223 VGND.n222 185
R1395 VGND.n225 VGND.n224 185
R1396 VGND.n227 VGND.n226 185
R1397 VGND.n229 VGND.n228 185
R1398 VGND.n231 VGND.n230 185
R1399 VGND.n233 VGND.n232 185
R1400 VGND.n235 VGND.n234 185
R1401 VGND.n237 VGND.n236 185
R1402 VGND.n239 VGND.n238 185
R1403 VGND.n205 VGND.n204 185
R1404 VGND.n207 VGND.n206 185
R1405 VGND.n209 VGND.n208 185
R1406 VGND.n211 VGND.n210 185
R1407 VGND.n213 VGND.n212 185
R1408 VGND.n215 VGND.n214 185
R1409 VGND.n217 VGND.n216 185
R1410 VGND.n219 VGND.n218 185
R1411 VGND.n221 VGND.n220 185
R1412 VGND.n203 VGND.n202 185
R1413 VGND.n197 VGND.n196 185
R1414 VGND.n195 VGND.n194 185
R1415 VGND.n190 VGND.n189 185
R1416 VGND.n188 VGND.n187 185
R1417 VGND.n183 VGND.n182 185
R1418 VGND.n179 VGND.n158 185
R1419 VGND.n262 VGND.n261 185
R1420 VGND.n157 VGND.n155 185
R1421 VGND.n707 VGND.n672 180.118
R1422 VGND.n1045 VGND.n1044 175.546
R1423 VGND.n1047 VGND.n1045 175.546
R1424 VGND.n1051 VGND.n437 175.546
R1425 VGND.n1055 VGND.n1053 175.546
R1426 VGND.n1059 VGND.n435 175.546
R1427 VGND.n1062 VGND.n1061 175.546
R1428 VGND.n1038 VGND.n440 175.546
R1429 VGND.n1038 VGND.n442 175.546
R1430 VGND.n1034 VGND.n442 175.546
R1431 VGND.n1034 VGND.n445 175.546
R1432 VGND.n1030 VGND.n445 175.546
R1433 VGND.n1030 VGND.n447 175.546
R1434 VGND.n1026 VGND.n447 175.546
R1435 VGND.n1026 VGND.n449 175.546
R1436 VGND.n1022 VGND.n449 175.546
R1437 VGND.n1022 VGND.n1019 175.546
R1438 VGND.n1019 VGND.n1018 175.546
R1439 VGND.n984 VGND.n983 175.546
R1440 VGND.n989 VGND.n986 175.546
R1441 VGND.n992 VGND.n991 175.546
R1442 VGND.n996 VGND.n994 175.546
R1443 VGND.n1109 VGND.n357 175.546
R1444 VGND.n2048 VGND.n1980 175.546
R1445 VGND.n1985 VGND.n1984 175.546
R1446 VGND.n1990 VGND.n1987 175.546
R1447 VGND.n1993 VGND.n1992 175.546
R1448 VGND.n1997 VGND.n1995 175.546
R1449 VGND.n2110 VGND.n1900 175.546
R1450 VGND.n2114 VGND.n2112 175.546
R1451 VGND.n2125 VGND.n1895 175.546
R1452 VGND.n2129 VGND.n2127 175.546
R1453 VGND.n2140 VGND.n1888 175.546
R1454 VGND.n2077 VGND.n1968 175.546
R1455 VGND.n2081 VGND.n2079 175.546
R1456 VGND.n2085 VGND.n1966 175.546
R1457 VGND.n2089 VGND.n2087 175.546
R1458 VGND.n2093 VGND.n1964 175.546
R1459 VGND.n2094 VGND.n2093 175.546
R1460 VGND.n2069 VGND.n1970 175.546
R1461 VGND.n2065 VGND.n2064 175.546
R1462 VGND.n2062 VGND.n1973 175.546
R1463 VGND.n2058 VGND.n2057 175.546
R1464 VGND.n2055 VGND.n1976 175.546
R1465 VGND.n2046 VGND.n2017 175.546
R1466 VGND.n2015 VGND.n1982 175.546
R1467 VGND.n2011 VGND.n2009 175.546
R1468 VGND.n2007 VGND.n1989 175.546
R1469 VGND.n2003 VGND.n2001 175.546
R1470 VGND.n2041 VGND.n2019 175.546
R1471 VGND.n2037 VGND.n2036 175.546
R1472 VGND.n2034 VGND.n2022 175.546
R1473 VGND.n2030 VGND.n2029 175.546
R1474 VGND.n2027 VGND.n2025 175.546
R1475 VGND.n2159 VGND.n1821 175.546
R1476 VGND.n2163 VGND.n2161 175.546
R1477 VGND.n2174 VGND.n1816 175.546
R1478 VGND.n2178 VGND.n2176 175.546
R1479 VGND.n2189 VGND.n1809 175.546
R1480 VGND.n2296 VGND.n1676 175.546
R1481 VGND.n1793 VGND.n1786 175.546
R1482 VGND.n1797 VGND.n1795 175.546
R1483 VGND.n1805 VGND.n1781 175.546
R1484 VGND.n2195 VGND.n1807 175.546
R1485 VGND.n493 VGND.n484 175.546
R1486 VGND.n489 VGND.n484 175.546
R1487 VGND.n489 VGND.n486 175.546
R1488 VGND.n486 VGND.n27 175.546
R1489 VGND.n2336 VGND.n27 175.546
R1490 VGND.n2336 VGND.n25 175.546
R1491 VGND.n2340 VGND.n25 175.546
R1492 VGND.n2340 VGND.n23 175.546
R1493 VGND.n2344 VGND.n23 175.546
R1494 VGND.n2344 VGND.n19 175.546
R1495 VGND.n2349 VGND.n19 175.546
R1496 VGND.n517 VGND.n471 175.546
R1497 VGND.n513 VGND.n471 175.546
R1498 VGND.n513 VGND.n473 175.546
R1499 VGND.n509 VGND.n473 175.546
R1500 VGND.n509 VGND.n476 175.546
R1501 VGND.n505 VGND.n476 175.546
R1502 VGND.n505 VGND.n478 175.546
R1503 VGND.n501 VGND.n478 175.546
R1504 VGND.n501 VGND.n480 175.546
R1505 VGND.n497 VGND.n480 175.546
R1506 VGND.n497 VGND.n482 175.546
R1507 VGND.n559 VGND.n558 175.546
R1508 VGND.n555 VGND.n554 175.546
R1509 VGND.n552 VGND.n525 175.546
R1510 VGND.n548 VGND.n546 175.546
R1511 VGND.n544 VGND.n534 175.546
R1512 VGND.n1012 VGND.n1011 175.546
R1513 VGND.n1008 VGND.n1007 175.546
R1514 VGND.n1005 VGND.n988 175.546
R1515 VGND.n1001 VGND.n999 175.546
R1516 VGND.n1111 VGND.n355 175.546
R1517 VGND.n980 VGND.n979 175.546
R1518 VGND.n979 VGND.n454 175.546
R1519 VGND.n975 VGND.n454 175.546
R1520 VGND.n975 VGND.n457 175.546
R1521 VGND.n971 VGND.n457 175.546
R1522 VGND.n971 VGND.n460 175.546
R1523 VGND.n573 VGND.n460 175.546
R1524 VGND.n573 VGND.n463 175.546
R1525 VGND.n569 VGND.n463 175.546
R1526 VGND.n569 VGND.n466 175.546
R1527 VGND.n565 VGND.n466 175.546
R1528 VGND.n521 VGND.n520 175.546
R1529 VGND.n526 VGND.n523 175.546
R1530 VGND.n529 VGND.n528 175.546
R1531 VGND.n535 VGND.n531 175.546
R1532 VGND.n538 VGND.n537 175.546
R1533 VGND.n1119 VGND.n1118 175.546
R1534 VGND.n1128 VGND.n1127 175.546
R1535 VGND.n1131 VGND.n1130 175.546
R1536 VGND.n1142 VGND.n1141 175.546
R1537 VGND.n1154 VGND.n278 175.546
R1538 VGND.n1091 VGND.n1090 175.546
R1539 VGND.n1087 VGND.n1086 175.546
R1540 VGND.n1080 VGND.n1079 175.546
R1541 VGND.n1073 VGND.n1072 175.546
R1542 VGND.n1101 VGND.n1100 175.546
R1543 VGND.n1611 VGND.n1163 175.546
R1544 VGND.n1607 VGND.n1163 175.546
R1545 VGND.n1607 VGND.n1165 175.546
R1546 VGND.n1603 VGND.n1165 175.546
R1547 VGND.n1603 VGND.n1601 175.546
R1548 VGND.n1601 VGND.n1600 175.546
R1549 VGND.n1600 VGND.n1168 175.546
R1550 VGND.n1596 VGND.n1168 175.546
R1551 VGND.n1596 VGND.n1170 175.546
R1552 VGND.n1592 VGND.n1170 175.546
R1553 VGND.n1592 VGND.n1173 175.546
R1554 VGND.n1645 VGND.n120 175.546
R1555 VGND.n1649 VGND.n1647 175.546
R1556 VGND.n1659 VGND.n116 175.546
R1557 VGND.n1662 VGND.n1661 175.546
R1558 VGND.n1664 VGND.n114 175.546
R1559 VGND.n1632 VGND.n1631 175.546
R1560 VGND.n1628 VGND.n1627 175.546
R1561 VGND.n1624 VGND.n1623 175.546
R1562 VGND.n1620 VGND.n1619 175.546
R1563 VGND.n1616 VGND.n1615 175.546
R1564 VGND.n1643 VGND.n1641 175.546
R1565 VGND.n1651 VGND.n118 175.546
R1566 VGND.n1657 VGND.n1653 175.546
R1567 VGND.n1655 VGND.n1654 175.546
R1568 VGND.n1667 VGND.n1666 175.546
R1569 VGND.n2326 VGND.n2325 175.546
R1570 VGND.n2322 VGND.n2321 175.546
R1571 VGND.n2319 VGND.n86 175.546
R1572 VGND.n2315 VGND.n2313 175.546
R1573 VGND.n2311 VGND.n94 175.546
R1574 VGND.n125 VGND.n124 175.546
R1575 VGND.n129 VGND.n128 175.546
R1576 VGND.n133 VGND.n132 175.546
R1577 VGND.n137 VGND.n136 175.546
R1578 VGND.n141 VGND.n140 175.546
R1579 VGND.n82 VGND.n81 175.546
R1580 VGND.n87 VGND.n84 175.546
R1581 VGND.n90 VGND.n89 175.546
R1582 VGND.n95 VGND.n92 175.546
R1583 VGND.n98 VGND.n97 175.546
R1584 VGND.n1333 VGND.n1331 175.546
R1585 VGND.n1337 VGND.n1306 175.546
R1586 VGND.n1341 VGND.n1339 175.546
R1587 VGND.n1345 VGND.n1304 175.546
R1588 VGND.n1348 VGND.n1347 175.546
R1589 VGND.n1325 VGND.n1324 175.546
R1590 VGND.n1321 VGND.n1320 175.546
R1591 VGND.n1317 VGND.n1316 175.546
R1592 VGND.n1313 VGND.n1312 175.546
R1593 VGND.n1309 VGND.n72 175.546
R1594 VGND.n1555 VGND.n1482 175.546
R1595 VGND.n1559 VGND.n1557 175.546
R1596 VGND.n1570 VGND.n1476 175.546
R1597 VGND.n1574 VGND.n1572 175.546
R1598 VGND.n1585 VGND.n1469 175.546
R1599 VGND.n1293 VGND.n1181 175.546
R1600 VGND.n1286 VGND.n1285 175.546
R1601 VGND.n1211 VGND.n1210 175.546
R1602 VGND.n1216 VGND.n1215 175.546
R1603 VGND.n1224 VGND.n1223 175.546
R1604 VGND.n1353 VGND.n1300 175.546
R1605 VGND.n1457 VGND.n1456 175.546
R1606 VGND.n1383 VGND.n1382 175.546
R1607 VGND.n1388 VGND.n1387 175.546
R1608 VGND.n1396 VGND.n1395 175.546
R1609 VGND.n2270 VGND.n2269 175.546
R1610 VGND.n2269 VGND.n1688 175.546
R1611 VGND.n2265 VGND.n1688 175.546
R1612 VGND.n2265 VGND.n1691 175.546
R1613 VGND.n2261 VGND.n1691 175.546
R1614 VGND.n2261 VGND.n2260 175.546
R1615 VGND.n2260 VGND.n2259 175.546
R1616 VGND.n2259 VGND.n1694 175.546
R1617 VGND.n2255 VGND.n1694 175.546
R1618 VGND.n2255 VGND.n1697 175.546
R1619 VGND.n2250 VGND.n1697 175.546
R1620 VGND.n2214 VGND.n1713 175.546
R1621 VGND.n2218 VGND.n2216 175.546
R1622 VGND.n2229 VGND.n1708 175.546
R1623 VGND.n2233 VGND.n2231 175.546
R1624 VGND.n2244 VGND.n1701 175.546
R1625 VGND.n2294 VGND.n1678 175.546
R1626 VGND.n1791 VGND.n1789 175.546
R1627 VGND.n1799 VGND.n1783 175.546
R1628 VGND.n1803 VGND.n1801 175.546
R1629 VGND.n2197 VGND.n1779 175.546
R1630 VGND.n2289 VGND.n1679 175.546
R1631 VGND.n2285 VGND.n2284 175.546
R1632 VGND.n2282 VGND.n1682 175.546
R1633 VGND.n2278 VGND.n2277 175.546
R1634 VGND.n2275 VGND.n1685 175.546
R1635 VGND.n264 VGND.n148 175.546
R1636 VGND.n180 VGND.n154 175.546
R1637 VGND.n185 VGND.n184 175.546
R1638 VGND.n192 VGND.n191 175.546
R1639 VGND.n200 VGND.n199 175.546
R1640 VGND.t193 VGND.n50 172.876
R1641 VGND.t193 VGND.n52 172.876
R1642 VGND.t193 VGND.n39 172.876
R1643 VGND.t193 VGND.n51 172.615
R1644 VGND.t193 VGND.n53 172.615
R1645 VGND.t193 VGND.n37 172.615
R1646 VGND.n844 VGND.n843 167.743
R1647 VGND.t270 VGND.n672 167.251
R1648 VGND.n809 VGND.n808 166.63
R1649 VGND.n789 VGND.n788 166.63
R1650 VGND.n2136 VGND.n2135 163.333
R1651 VGND.n2185 VGND.n2184 163.333
R1652 VGND.n1149 VGND.n1148 163.333
R1653 VGND.n372 VGND.n362 163.333
R1654 VGND.n1581 VGND.n1580 163.333
R1655 VGND.n1228 VGND.n1227 163.333
R1656 VGND.n1400 VGND.n1399 163.333
R1657 VGND.n2240 VGND.n2239 163.333
R1658 VGND.n204 VGND.n203 163.333
R1659 VGND.n969 VGND.n576 157.601
R1660 VGND.t155 VGND.t69 154.649
R1661 VGND.n894 VGND.n890 153.601
R1662 VGND.t37 VGND.t41 152.681
R1663 VGND.t34 VGND.t37 152.681
R1664 VGND.t129 VGND.t153 152.681
R1665 VGND.t248 VGND.t129 152.681
R1666 VGND.t256 VGND.t248 152.681
R1667 VGND.t109 VGND.t298 152.681
R1668 VGND.t21 VGND.t109 152.681
R1669 VGND.t146 VGND.t141 152.681
R1670 VGND.t139 VGND.t146 152.681
R1671 VGND.t276 VGND.t139 152.681
R1672 VGND.t133 VGND.t144 152.681
R1673 VGND.t144 VGND.t245 152.681
R1674 VGND.t77 VGND.t107 152.681
R1675 VGND.t107 VGND.t79 152.681
R1676 VGND.t79 VGND.t5 152.681
R1677 VGND.t23 VGND.t96 152.681
R1678 VGND.t104 VGND.t23 152.681
R1679 VGND.t13 VGND.t278 152.681
R1680 VGND.t289 VGND.t13 152.681
R1681 VGND.t177 VGND.t289 152.681
R1682 VGND.t28 VGND.t120 152.681
R1683 VGND.t148 VGND.t28 152.681
R1684 VGND.t291 VGND.t254 152.681
R1685 VGND.t254 VGND.t266 152.681
R1686 VGND.t266 VGND.t121 152.681
R1687 VGND.t102 VGND.t281 152.681
R1688 VGND.t283 VGND.t100 152.681
R1689 VGND.t44 VGND.t283 152.681
R1690 VGND.t67 VGND.t44 152.681
R1691 VGND.t187 VGND.t85 152.681
R1692 VGND.t157 VGND.t187 152.681
R1693 VGND.t65 VGND.t157 152.681
R1694 VGND.t71 VGND.t25 152.681
R1695 VGND.t118 VGND.t71 152.681
R1696 VGND.t131 VGND.t118 152.681
R1697 VGND.t11 VGND.t35 152.681
R1698 VGND.t105 VGND.t190 152.681
R1699 VGND.t166 VGND.t105 152.681
R1700 VGND.t246 VGND.t166 152.681
R1701 VGND.n959 VGND.t58 150.249
R1702 VGND.n1944 VGND.n1942 150
R1703 VGND.n1940 VGND.n1908 150
R1704 VGND.n1936 VGND.n1934 150
R1705 VGND.n1932 VGND.n1910 150
R1706 VGND.n1928 VGND.n1926 150
R1707 VGND.n1924 VGND.n1912 150
R1708 VGND.n1920 VGND.n1919 150
R1709 VGND.n1917 VGND.n1915 150
R1710 VGND.n2107 VGND.n2105 150
R1711 VGND.n2118 VGND.n1897 150
R1712 VGND.n2122 VGND.n2120 150
R1713 VGND.n2133 VGND.n1892 150
R1714 VGND.n1952 VGND.n1950 150
R1715 VGND.n1956 VGND.n1904 150
R1716 VGND.n1960 VGND.n1958 150
R1717 VGND.n2103 VGND.n1902 150
R1718 VGND.n1865 VGND.n1863 150
R1719 VGND.n1861 VGND.n1829 150
R1720 VGND.n1857 VGND.n1855 150
R1721 VGND.n1853 VGND.n1831 150
R1722 VGND.n1849 VGND.n1847 150
R1723 VGND.n1845 VGND.n1833 150
R1724 VGND.n1841 VGND.n1840 150
R1725 VGND.n1838 VGND.n1836 150
R1726 VGND.n2156 VGND.n2154 150
R1727 VGND.n2167 VGND.n1818 150
R1728 VGND.n2171 VGND.n2169 150
R1729 VGND.n2182 VGND.n1813 150
R1730 VGND.n1873 VGND.n1871 150
R1731 VGND.n1877 VGND.n1825 150
R1732 VGND.n1881 VGND.n1879 150
R1733 VGND.n2152 VGND.n1823 150
R1734 VGND.n332 VGND.n295 150
R1735 VGND.n328 VGND.n326 150
R1736 VGND.n324 VGND.n297 150
R1737 VGND.n320 VGND.n318 150
R1738 VGND.n316 VGND.n299 150
R1739 VGND.n312 VGND.n311 150
R1740 VGND.n309 VGND.n302 150
R1741 VGND.n305 VGND.n304 150
R1742 VGND.n1124 VGND.n1122 150
R1743 VGND.n1134 VGND.n286 150
R1744 VGND.n1138 VGND.n1136 150
R1745 VGND.n1146 VGND.n282 150
R1746 VGND.n340 VGND.n293 150
R1747 VGND.n344 VGND.n342 150
R1748 VGND.n348 VGND.n291 150
R1749 VGND.n351 VGND.n350 150
R1750 VGND.n412 VGND.n411 150
R1751 VGND.n408 VGND.n407 150
R1752 VGND.n404 VGND.n403 150
R1753 VGND.n400 VGND.n399 150
R1754 VGND.n396 VGND.n395 150
R1755 VGND.n392 VGND.n391 150
R1756 VGND.n388 VGND.n387 150
R1757 VGND.n384 VGND.n383 150
R1758 VGND.n1094 VGND.n381 150
R1759 VGND.n1083 VGND.n1082 150
R1760 VGND.n1076 VGND.n1075 150
R1761 VGND.n1097 VGND.n361 150
R1762 VGND.n420 VGND.n419 150
R1763 VGND.n424 VGND.n423 150
R1764 VGND.n428 VGND.n427 150
R1765 VGND.n430 VGND.n380 150
R1766 VGND.n1526 VGND.n1524 150
R1767 VGND.n1522 VGND.n1490 150
R1768 VGND.n1518 VGND.n1516 150
R1769 VGND.n1514 VGND.n1492 150
R1770 VGND.n1510 VGND.n1508 150
R1771 VGND.n1506 VGND.n1494 150
R1772 VGND.n1502 VGND.n1501 150
R1773 VGND.n1499 VGND.n1497 150
R1774 VGND.n1552 VGND.n1550 150
R1775 VGND.n1563 VGND.n1478 150
R1776 VGND.n1567 VGND.n1565 150
R1777 VGND.n1578 VGND.n1473 150
R1778 VGND.n1534 VGND.n1532 150
R1779 VGND.n1538 VGND.n1486 150
R1780 VGND.n1542 VGND.n1540 150
R1781 VGND.n1548 VGND.n1484 150
R1782 VGND.n1260 VGND.n1259 150
R1783 VGND.n1256 VGND.n1255 150
R1784 VGND.n1252 VGND.n1251 150
R1785 VGND.n1248 VGND.n1247 150
R1786 VGND.n1244 VGND.n1243 150
R1787 VGND.n1240 VGND.n1239 150
R1788 VGND.n1236 VGND.n1235 150
R1789 VGND.n1232 VGND.n1231 150
R1790 VGND.n1290 VGND.n1289 150
R1791 VGND.n1282 VGND.n1189 150
R1792 VGND.n1213 VGND.n1190 150
R1793 VGND.n1220 VGND.n1219 150
R1794 VGND.n1279 VGND.n1206 150
R1795 VGND.n1275 VGND.n1274 150
R1796 VGND.n1271 VGND.n1270 150
R1797 VGND.n1267 VGND.n1266 150
R1798 VGND.n1432 VGND.n1431 150
R1799 VGND.n1428 VGND.n1427 150
R1800 VGND.n1424 VGND.n1423 150
R1801 VGND.n1420 VGND.n1419 150
R1802 VGND.n1416 VGND.n1415 150
R1803 VGND.n1412 VGND.n1411 150
R1804 VGND.n1408 VGND.n1407 150
R1805 VGND.n1404 VGND.n1403 150
R1806 VGND.n1461 VGND.n1460 150
R1807 VGND.n1453 VGND.n1359 150
R1808 VGND.n1385 VGND.n1360 150
R1809 VGND.n1392 VGND.n1391 150
R1810 VGND.n1450 VGND.n1376 150
R1811 VGND.n1446 VGND.n1445 150
R1812 VGND.n1442 VGND.n1441 150
R1813 VGND.n1438 VGND.n1437 150
R1814 VGND.n1757 VGND.n1755 150
R1815 VGND.n1753 VGND.n1721 150
R1816 VGND.n1749 VGND.n1747 150
R1817 VGND.n1745 VGND.n1723 150
R1818 VGND.n1741 VGND.n1739 150
R1819 VGND.n1737 VGND.n1725 150
R1820 VGND.n1733 VGND.n1732 150
R1821 VGND.n1730 VGND.n1728 150
R1822 VGND.n2211 VGND.n2209 150
R1823 VGND.n2222 VGND.n1710 150
R1824 VGND.n2226 VGND.n2224 150
R1825 VGND.n2237 VGND.n1705 150
R1826 VGND.n1765 VGND.n1763 150
R1827 VGND.n1769 VGND.n1717 150
R1828 VGND.n1773 VGND.n1771 150
R1829 VGND.n2207 VGND.n1715 150
R1830 VGND.n236 VGND.n235 150
R1831 VGND.n232 VGND.n231 150
R1832 VGND.n228 VGND.n227 150
R1833 VGND.n224 VGND.n223 150
R1834 VGND.n220 VGND.n219 150
R1835 VGND.n216 VGND.n215 150
R1836 VGND.n212 VGND.n211 150
R1837 VGND.n208 VGND.n207 150
R1838 VGND.n261 VGND.n157 150
R1839 VGND.n182 VGND.n158 150
R1840 VGND.n189 VGND.n188 150
R1841 VGND.n196 VGND.n195 150
R1842 VGND.n244 VGND.n243 150
R1843 VGND.n248 VGND.n247 150
R1844 VGND.n252 VGND.n251 150
R1845 VGND.n258 VGND.n175 150
R1846 VGND.n896 VGND.n895 146.25
R1847 VGND.n897 VGND.n896 146.25
R1848 VGND.n883 VGND.n882 146.25
R1849 VGND.n882 VGND.n881 146.25
R1850 VGND.n885 VGND.n884 144
R1851 VGND.n877 VGND.t170 134.954
R1852 VGND.n891 VGND.t188 134.651
R1853 VGND.n875 VGND.t189 134.651
R1854 VGND.n878 VGND.t57 134.651
R1855 VGND.n892 VGND.t103 134.62
R1856 VGND.n876 VGND.t251 134.62
R1857 VGND.n879 VGND.t47 134.62
R1858 VGND.n847 VGND.t226 134.501
R1859 VGND.n860 VGND.t210 134.501
R1860 VGND.n650 VGND.n649 134.268
R1861 VGND.n650 VGND.n643 134.268
R1862 VGND.n1350 VGND.n1349 132.721
R1863 VGND.n960 VGND.t73 131.468
R1864 VGND.n890 VGND.n874 131.201
R1865 VGND.n705 VGND.t50 130.713
R1866 VGND.n711 VGND.t117 130.001
R1867 VGND.n721 VGND.t99 130.001
R1868 VGND.n723 VGND.t184 130.001
R1869 VGND.n726 VGND.t52 130.001
R1870 VGND.n729 VGND.t20 130.001
R1871 VGND.n708 VGND.t115 130.001
R1872 VGND.n697 VGND.t54 130.001
R1873 VGND.n694 VGND.t288 130.001
R1874 VGND.n692 VGND.t64 130.001
R1875 VGND.n689 VGND.t56 130.001
R1876 VGND.n716 VGND.t275 130.001
R1877 VGND.n714 VGND.t297 130.001
R1878 VGND.n673 VGND.t271 130.001
R1879 VGND.t125 VGND.t237 129.706
R1880 VGND.t150 VGND.t175 129.706
R1881 VGND.t224 VGND.t39 129.706
R1882 VGND.n845 VGND.t205 125.066
R1883 VGND.n1107 VGND.n1106 124.832
R1884 VGND.n2143 VGND.n1886 124.832
R1885 VGND.n2145 VGND.n1885 124.832
R1886 VGND.n2193 VGND.n2192 124.832
R1887 VGND.n1159 VGND.n146 124.832
R1888 VGND.n1114 VGND.n1113 124.832
R1889 VGND.n540 VGND.n145 124.832
R1890 VGND.n2303 VGND.n106 124.832
R1891 VGND.n1669 VGND.n105 124.832
R1892 VGND.n2307 VGND.n2305 124.832
R1893 VGND.n104 VGND.n100 124.832
R1894 VGND.n2200 VGND.n2199 124.832
R1895 VGND.n773 VGND.t75 124.718
R1896 VGND.t209 VGND.t93 124.718
R1897 VGND.n869 VGND.n868 122.582
R1898 VGND.n731 VGND.t138 122.501
R1899 VGND.n734 VGND.t244 122.501
R1900 VGND.n736 VGND.t273 122.501
R1901 VGND.n680 VGND.t152 122.501
R1902 VGND.n677 VGND.t263 122.501
R1903 VGND.n683 VGND.t124 122.501
R1904 VGND.t15 VGND.n772 119.728
R1905 VGND.t264 VGND.n857 119.728
R1906 VGND.n654 VGND.n653 117.209
R1907 VGND.n653 VGND.t58 117.209
R1908 VGND.n661 VGND.n588 117.209
R1909 VGND.n819 VGND.t135 114.74
R1910 VGND.n961 VGND.t74 110.925
R1911 VGND.n16 VGND.t176 110.826
R1912 VGND.n962 VGND.t87 110.659
R1913 VGND.n965 VGND.t295 110.591
R1914 VGND.t197 VGND.t48 104.763
R1915 VGND.n844 VGND.n842 104.328
R1916 VGND.n1156 VGND.n54 103.144
R1917 VGND.n851 VGND.n850 102.136
R1918 VGND.n756 VGND.n755 102.136
R1919 VGND.n754 VGND.n753 102.136
R1920 VGND.n752 VGND.n751 102.136
R1921 VGND.n859 VGND.n744 102.136
R1922 VGND.n772 VGND.t285 99.7737
R1923 VGND.t193 VGND.n44 47.6748
R1924 VGND.n2334 VGND.n54 99.6276
R1925 VGND.n619 VGND.n609 93.7671
R1926 VGND.t193 VGND.n2334 91.423
R1927 VGND.n816 VGND.n811 91.3721
R1928 VGND.n824 VGND.n807 91.3721
R1929 VGND.n824 VGND.n823 91.3721
R1930 VGND.n792 VGND.n791 91.3721
R1931 VGND.n801 VGND.n787 91.3721
R1932 VGND.n801 VGND.n800 91.3721
R1933 VGND.n657 VGND.n594 91.069
R1934 VGND.n658 VGND.n657 91.069
R1935 VGND.n636 VGND.n635 91.069
R1936 VGND.n635 VGND.n591 91.069
R1937 VGND.n649 VGND.n648 91.069
R1938 VGND.n644 VGND.n643 91.069
R1939 VGND.n682 VGND.n681 90.9566
R1940 VGND.n839 VGND.n833 90.7567
R1941 VGND.n781 VGND.n764 90.7567
R1942 VGND.t73 VGND.t22 90.149
R1943 VGND.t22 VGND.t168 90.149
R1944 VGND.t168 VGND.t86 90.149
R1945 VGND.t164 VGND.t216 89.7964
R1946 VGND.n869 VGND.t9 84.8078
R1947 VGND.t75 VGND.t233 84.8078
R1948 VGND.t48 VGND.t81 84.8078
R1949 VGND.n798 VGND.n746 84.306
R1950 VGND.n797 VGND.n745 84.306
R1951 VGND.n818 VGND.n812 84.306
R1952 VGND.n821 VGND.n820 84.306
R1953 VGND.n774 VGND.n769 84.306
R1954 VGND.n775 VGND.n774 84.306
R1955 VGND.n841 VGND.n762 84.306
R1956 VGND.n854 VGND.n853 83.2005
R1957 VGND.n853 VGND.n750 83.2005
R1958 VGND.t205 VGND.n844 82.8853
R1959 VGND.t0 VGND.n584 82.0463
R1960 VGND.n1043 VGND.n1042 76.3222
R1961 VGND.n1047 VGND.n1046 76.3222
R1962 VGND.n1052 VGND.n1051 76.3222
R1963 VGND.n1055 VGND.n1054 76.3222
R1964 VGND.n1060 VGND.n1059 76.3222
R1965 VGND.n983 VGND.n982 76.3222
R1966 VGND.n986 VGND.n985 76.3222
R1967 VGND.n991 VGND.n990 76.3222
R1968 VGND.n994 VGND.n993 76.3222
R1969 VGND.n995 VGND.n357 76.3222
R1970 VGND.n1108 VGND.n1107 76.3222
R1971 VGND.n2049 VGND.n2048 76.3222
R1972 VGND.n1984 VGND.n1983 76.3222
R1973 VGND.n1987 VGND.n1986 76.3222
R1974 VGND.n1992 VGND.n1991 76.3222
R1975 VGND.n1995 VGND.n1994 76.3222
R1976 VGND.n1996 VGND.n1886 76.3222
R1977 VGND.n2098 VGND.n2097 76.3222
R1978 VGND.n2111 VGND.n2110 76.3222
R1979 VGND.n2114 VGND.n2113 76.3222
R1980 VGND.n2126 VGND.n2125 76.3222
R1981 VGND.n2129 VGND.n2128 76.3222
R1982 VGND.n2141 VGND.n2140 76.3222
R1983 VGND.n2073 VGND.n2072 76.3222
R1984 VGND.n2078 VGND.n2077 76.3222
R1985 VGND.n2081 VGND.n2080 76.3222
R1986 VGND.n2086 VGND.n2085 76.3222
R1987 VGND.n2089 VGND.n2088 76.3222
R1988 VGND.n2070 VGND.n2069 76.3222
R1989 VGND.n2065 VGND.n1972 76.3222
R1990 VGND.n2063 VGND.n2062 76.3222
R1991 VGND.n2058 VGND.n1975 76.3222
R1992 VGND.n2056 VGND.n2055 76.3222
R1993 VGND.n2051 VGND.n1978 76.3222
R1994 VGND.n2045 VGND.n2044 76.3222
R1995 VGND.n2017 VGND.n2016 76.3222
R1996 VGND.n2010 VGND.n1982 76.3222
R1997 VGND.n2009 VGND.n2008 76.3222
R1998 VGND.n2002 VGND.n1989 76.3222
R1999 VGND.n2001 VGND.n2000 76.3222
R2000 VGND.n2042 VGND.n2041 76.3222
R2001 VGND.n2037 VGND.n2021 76.3222
R2002 VGND.n2035 VGND.n2034 76.3222
R2003 VGND.n2030 VGND.n2024 76.3222
R2004 VGND.n2028 VGND.n2027 76.3222
R2005 VGND.n2299 VGND.n1675 76.3222
R2006 VGND.n2147 VGND.n2146 76.3222
R2007 VGND.n2160 VGND.n2159 76.3222
R2008 VGND.n2163 VGND.n2162 76.3222
R2009 VGND.n2175 VGND.n2174 76.3222
R2010 VGND.n2178 VGND.n2177 76.3222
R2011 VGND.n2190 VGND.n2189 76.3222
R2012 VGND.n2297 VGND.n2296 76.3222
R2013 VGND.n1786 VGND.n1785 76.3222
R2014 VGND.n1795 VGND.n1794 76.3222
R2015 VGND.n1796 VGND.n1781 76.3222
R2016 VGND.n1807 VGND.n1806 76.3222
R2017 VGND.n2194 VGND.n2193 76.3222
R2018 VGND.n561 VGND.n560 76.3222
R2019 VGND.n558 VGND.n518 76.3222
R2020 VGND.n554 VGND.n553 76.3222
R2021 VGND.n547 VGND.n525 76.3222
R2022 VGND.n546 VGND.n545 76.3222
R2023 VGND.n534 VGND.n533 76.3222
R2024 VGND.n1014 VGND.n1013 76.3222
R2025 VGND.n1011 VGND.n981 76.3222
R2026 VGND.n1007 VGND.n1006 76.3222
R2027 VGND.n1000 VGND.n988 76.3222
R2028 VGND.n999 VGND.n998 76.3222
R2029 VGND.n1112 VGND.n1111 76.3222
R2030 VGND.n520 VGND.n519 76.3222
R2031 VGND.n523 VGND.n522 76.3222
R2032 VGND.n528 VGND.n527 76.3222
R2033 VGND.n531 VGND.n530 76.3222
R2034 VGND.n537 VGND.n536 76.3222
R2035 VGND.n540 VGND.n539 76.3222
R2036 VGND.n1115 VGND.n272 76.3222
R2037 VGND.n1118 VGND.n273 76.3222
R2038 VGND.n1128 VGND.n274 76.3222
R2039 VGND.n1130 VGND.n275 76.3222
R2040 VGND.n1142 VGND.n276 76.3222
R2041 VGND.n1155 VGND.n1154 76.3222
R2042 VGND.n1065 VGND.n266 76.3222
R2043 VGND.n1091 VGND.n267 76.3222
R2044 VGND.n1086 VGND.n268 76.3222
R2045 VGND.n1079 VGND.n269 76.3222
R2046 VGND.n1072 VGND.n270 76.3222
R2047 VGND.n1101 VGND.n271 76.3222
R2048 VGND.n1637 VGND.n1636 76.3222
R2049 VGND.n1646 VGND.n1645 76.3222
R2050 VGND.n1649 VGND.n1648 76.3222
R2051 VGND.n1660 VGND.n1659 76.3222
R2052 VGND.n1663 VGND.n1662 76.3222
R2053 VGND.n114 VGND.n113 76.3222
R2054 VGND.n1632 VGND.n55 76.3222
R2055 VGND.n1628 VGND.n56 76.3222
R2056 VGND.n1624 VGND.n57 76.3222
R2057 VGND.n1620 VGND.n58 76.3222
R2058 VGND.n1616 VGND.n59 76.3222
R2059 VGND.n1612 VGND.n60 76.3222
R2060 VGND.n1641 VGND.n1640 76.3222
R2061 VGND.n1642 VGND.n118 76.3222
R2062 VGND.n1653 VGND.n1652 76.3222
R2063 VGND.n1656 VGND.n1655 76.3222
R2064 VGND.n1666 VGND.n111 76.3222
R2065 VGND.n1669 VGND.n1668 76.3222
R2066 VGND.n2328 VGND.n2327 76.3222
R2067 VGND.n2325 VGND.n79 76.3222
R2068 VGND.n2321 VGND.n2320 76.3222
R2069 VGND.n2314 VGND.n86 76.3222
R2070 VGND.n2313 VGND.n2312 76.3222
R2071 VGND.n2306 VGND.n94 76.3222
R2072 VGND.n124 VGND.n61 76.3222
R2073 VGND.n128 VGND.n62 76.3222
R2074 VGND.n132 VGND.n63 76.3222
R2075 VGND.n136 VGND.n64 76.3222
R2076 VGND.n140 VGND.n65 76.3222
R2077 VGND.n122 VGND.n66 76.3222
R2078 VGND.n81 VGND.n80 76.3222
R2079 VGND.n84 VGND.n83 76.3222
R2080 VGND.n89 VGND.n88 76.3222
R2081 VGND.n92 VGND.n91 76.3222
R2082 VGND.n97 VGND.n96 76.3222
R2083 VGND.n100 VGND.n99 76.3222
R2084 VGND.n1330 VGND.n1329 76.3222
R2085 VGND.n1333 VGND.n1332 76.3222
R2086 VGND.n1338 VGND.n1337 76.3222
R2087 VGND.n1341 VGND.n1340 76.3222
R2088 VGND.n1346 VGND.n1345 76.3222
R2089 VGND.n1349 VGND.n1348 76.3222
R2090 VGND.n1325 VGND.n67 76.3222
R2091 VGND.n1321 VGND.n68 76.3222
R2092 VGND.n1317 VGND.n69 76.3222
R2093 VGND.n1313 VGND.n70 76.3222
R2094 VGND.n1309 VGND.n71 76.3222
R2095 VGND.n2333 VGND.n2332 76.3222
R2096 VGND.n1481 VGND.n107 76.3222
R2097 VGND.n1556 VGND.n1555 76.3222
R2098 VGND.n1559 VGND.n1558 76.3222
R2099 VGND.n1571 VGND.n1570 76.3222
R2100 VGND.n1574 VGND.n1573 76.3222
R2101 VGND.n1586 VGND.n1585 76.3222
R2102 VGND.n1294 VGND.n102 76.3222
R2103 VGND.n1181 VGND.n1180 76.3222
R2104 VGND.n1285 VGND.n1179 76.3222
R2105 VGND.n1211 VGND.n1178 76.3222
R2106 VGND.n1215 VGND.n1177 76.3222
R2107 VGND.n1224 VGND.n1176 76.3222
R2108 VGND.n1467 VGND.n1466 76.3222
R2109 VGND.n1353 VGND.n1299 76.3222
R2110 VGND.n1456 VGND.n1298 76.3222
R2111 VGND.n1383 VGND.n1297 76.3222
R2112 VGND.n1387 VGND.n1296 76.3222
R2113 VGND.n1396 VGND.n1295 76.3222
R2114 VGND.n2202 VGND.n2201 76.3222
R2115 VGND.n2215 VGND.n2214 76.3222
R2116 VGND.n2218 VGND.n2217 76.3222
R2117 VGND.n2230 VGND.n2229 76.3222
R2118 VGND.n2233 VGND.n2232 76.3222
R2119 VGND.n2245 VGND.n2244 76.3222
R2120 VGND.n2293 VGND.n2292 76.3222
R2121 VGND.n1788 VGND.n1678 76.3222
R2122 VGND.n1791 VGND.n1790 76.3222
R2123 VGND.n1800 VGND.n1799 76.3222
R2124 VGND.n1803 VGND.n1802 76.3222
R2125 VGND.n2198 VGND.n2197 76.3222
R2126 VGND.n2290 VGND.n2289 76.3222
R2127 VGND.n2285 VGND.n1681 76.3222
R2128 VGND.n2283 VGND.n2282 76.3222
R2129 VGND.n2278 VGND.n1684 76.3222
R2130 VGND.n2276 VGND.n2275 76.3222
R2131 VGND.n2271 VGND.n1687 76.3222
R2132 VGND.n1687 VGND.n1685 76.3222
R2133 VGND.n2277 VGND.n2276 76.3222
R2134 VGND.n1684 VGND.n1682 76.3222
R2135 VGND.n2284 VGND.n2283 76.3222
R2136 VGND.n1681 VGND.n1679 76.3222
R2137 VGND.n2291 VGND.n2290 76.3222
R2138 VGND.n1467 VGND.n1300 76.3222
R2139 VGND.n1457 VGND.n1299 76.3222
R2140 VGND.n1382 VGND.n1298 76.3222
R2141 VGND.n1388 VGND.n1297 76.3222
R2142 VGND.n1395 VGND.n1296 76.3222
R2143 VGND.n1377 VGND.n1295 76.3222
R2144 VGND.n1294 VGND.n1293 76.3222
R2145 VGND.n1286 VGND.n1180 76.3222
R2146 VGND.n1210 VGND.n1179 76.3222
R2147 VGND.n1216 VGND.n1178 76.3222
R2148 VGND.n1223 VGND.n1177 76.3222
R2149 VGND.n1176 VGND.n1175 76.3222
R2150 VGND.n1482 VGND.n1481 76.3222
R2151 VGND.n1557 VGND.n1556 76.3222
R2152 VGND.n1558 VGND.n1476 76.3222
R2153 VGND.n1572 VGND.n1571 76.3222
R2154 VGND.n1573 VGND.n1469 76.3222
R2155 VGND.n1587 VGND.n1586 76.3222
R2156 VGND.n2333 VGND.n72 76.3222
R2157 VGND.n1312 VGND.n71 76.3222
R2158 VGND.n1316 VGND.n70 76.3222
R2159 VGND.n1320 VGND.n69 76.3222
R2160 VGND.n1324 VGND.n68 76.3222
R2161 VGND.n1308 VGND.n67 76.3222
R2162 VGND.n141 VGND.n66 76.3222
R2163 VGND.n137 VGND.n65 76.3222
R2164 VGND.n133 VGND.n64 76.3222
R2165 VGND.n129 VGND.n63 76.3222
R2166 VGND.n125 VGND.n62 76.3222
R2167 VGND.n78 VGND.n61 76.3222
R2168 VGND.n1615 VGND.n60 76.3222
R2169 VGND.n1619 VGND.n59 76.3222
R2170 VGND.n1623 VGND.n58 76.3222
R2171 VGND.n1627 VGND.n57 76.3222
R2172 VGND.n1631 VGND.n56 76.3222
R2173 VGND.n1635 VGND.n55 76.3222
R2174 VGND.n1090 VGND.n266 76.3222
R2175 VGND.n1087 VGND.n267 76.3222
R2176 VGND.n1080 VGND.n268 76.3222
R2177 VGND.n1073 VGND.n269 76.3222
R2178 VGND.n1100 VGND.n270 76.3222
R2179 VGND.n1105 VGND.n271 76.3222
R2180 VGND.n1119 VGND.n272 76.3222
R2181 VGND.n1127 VGND.n273 76.3222
R2182 VGND.n1131 VGND.n274 76.3222
R2183 VGND.n1141 VGND.n275 76.3222
R2184 VGND.n278 VGND.n276 76.3222
R2185 VGND.n1155 VGND.n277 76.3222
R2186 VGND.n1157 VGND.n148 76.3222
R2187 VGND.n265 VGND.n154 76.3222
R2188 VGND.n185 VGND.n153 76.3222
R2189 VGND.n192 VGND.n152 76.3222
R2190 VGND.n199 VGND.n151 76.3222
R2191 VGND.n150 VGND.n149 76.3222
R2192 VGND.n1158 VGND.n1157 76.3222
R2193 VGND.n265 VGND.n264 76.3222
R2194 VGND.n180 VGND.n153 76.3222
R2195 VGND.n184 VGND.n152 76.3222
R2196 VGND.n191 VGND.n151 76.3222
R2197 VGND.n200 VGND.n150 76.3222
R2198 VGND.n539 VGND.n538 76.3222
R2199 VGND.n536 VGND.n535 76.3222
R2200 VGND.n530 VGND.n529 76.3222
R2201 VGND.n527 VGND.n526 76.3222
R2202 VGND.n522 VGND.n521 76.3222
R2203 VGND.n519 VGND.n468 76.3222
R2204 VGND.n560 VGND.n559 76.3222
R2205 VGND.n555 VGND.n518 76.3222
R2206 VGND.n553 VGND.n552 76.3222
R2207 VGND.n548 VGND.n547 76.3222
R2208 VGND.n545 VGND.n544 76.3222
R2209 VGND.n533 VGND.n146 76.3222
R2210 VGND.n1668 VGND.n1667 76.3222
R2211 VGND.n1654 VGND.n111 76.3222
R2212 VGND.n1657 VGND.n1656 76.3222
R2213 VGND.n1652 VGND.n1651 76.3222
R2214 VGND.n1643 VGND.n1642 76.3222
R2215 VGND.n1640 VGND.n1639 76.3222
R2216 VGND.n1636 VGND.n120 76.3222
R2217 VGND.n1647 VGND.n1646 76.3222
R2218 VGND.n1648 VGND.n116 76.3222
R2219 VGND.n1661 VGND.n1660 76.3222
R2220 VGND.n1664 VGND.n1663 76.3222
R2221 VGND.n113 VGND.n106 76.3222
R2222 VGND.n2195 VGND.n2194 76.3222
R2223 VGND.n1806 VGND.n1805 76.3222
R2224 VGND.n1797 VGND.n1796 76.3222
R2225 VGND.n1794 VGND.n1793 76.3222
R2226 VGND.n1785 VGND.n1676 76.3222
R2227 VGND.n2298 VGND.n2297 76.3222
R2228 VGND.n2294 VGND.n2293 76.3222
R2229 VGND.n1789 VGND.n1788 76.3222
R2230 VGND.n1790 VGND.n1783 76.3222
R2231 VGND.n1801 VGND.n1800 76.3222
R2232 VGND.n1802 VGND.n1779 76.3222
R2233 VGND.n2199 VGND.n2198 76.3222
R2234 VGND.n2025 VGND.n1675 76.3222
R2235 VGND.n2029 VGND.n2028 76.3222
R2236 VGND.n2024 VGND.n2022 76.3222
R2237 VGND.n2036 VGND.n2035 76.3222
R2238 VGND.n2021 VGND.n2019 76.3222
R2239 VGND.n2043 VGND.n2042 76.3222
R2240 VGND.n1978 VGND.n1976 76.3222
R2241 VGND.n2057 VGND.n2056 76.3222
R2242 VGND.n1975 VGND.n1973 76.3222
R2243 VGND.n2064 VGND.n2063 76.3222
R2244 VGND.n1972 VGND.n1970 76.3222
R2245 VGND.n2071 VGND.n2070 76.3222
R2246 VGND.n1997 VGND.n1996 76.3222
R2247 VGND.n1994 VGND.n1993 76.3222
R2248 VGND.n1991 VGND.n1990 76.3222
R2249 VGND.n1986 VGND.n1985 76.3222
R2250 VGND.n1983 VGND.n1980 76.3222
R2251 VGND.n2050 VGND.n2049 76.3222
R2252 VGND.n2046 VGND.n2045 76.3222
R2253 VGND.n2016 VGND.n2015 76.3222
R2254 VGND.n2011 VGND.n2010 76.3222
R2255 VGND.n2008 VGND.n2007 76.3222
R2256 VGND.n2003 VGND.n2002 76.3222
R2257 VGND.n2000 VGND.n1885 76.3222
R2258 VGND.n99 VGND.n98 76.3222
R2259 VGND.n96 VGND.n95 76.3222
R2260 VGND.n91 VGND.n90 76.3222
R2261 VGND.n88 VGND.n87 76.3222
R2262 VGND.n83 VGND.n82 76.3222
R2263 VGND.n80 VGND.n73 76.3222
R2264 VGND.n2327 VGND.n2326 76.3222
R2265 VGND.n2322 VGND.n79 76.3222
R2266 VGND.n2320 VGND.n2319 76.3222
R2267 VGND.n2315 VGND.n2314 76.3222
R2268 VGND.n2312 VGND.n2311 76.3222
R2269 VGND.n2307 VGND.n2306 76.3222
R2270 VGND.n1109 VGND.n1108 76.3222
R2271 VGND.n996 VGND.n995 76.3222
R2272 VGND.n993 VGND.n992 76.3222
R2273 VGND.n990 VGND.n989 76.3222
R2274 VGND.n985 VGND.n984 76.3222
R2275 VGND.n982 VGND.n451 76.3222
R2276 VGND.n1013 VGND.n1012 76.3222
R2277 VGND.n1008 VGND.n981 76.3222
R2278 VGND.n1006 VGND.n1005 76.3222
R2279 VGND.n1001 VGND.n1000 76.3222
R2280 VGND.n998 VGND.n355 76.3222
R2281 VGND.n1113 VGND.n1112 76.3222
R2282 VGND.n2097 VGND.n1900 76.3222
R2283 VGND.n2112 VGND.n2111 76.3222
R2284 VGND.n2113 VGND.n1895 76.3222
R2285 VGND.n2127 VGND.n2126 76.3222
R2286 VGND.n2128 VGND.n1888 76.3222
R2287 VGND.n2142 VGND.n2141 76.3222
R2288 VGND.n2146 VGND.n1821 76.3222
R2289 VGND.n2161 VGND.n2160 76.3222
R2290 VGND.n2162 VGND.n1816 76.3222
R2291 VGND.n2176 VGND.n2175 76.3222
R2292 VGND.n2177 VGND.n1809 76.3222
R2293 VGND.n2191 VGND.n2190 76.3222
R2294 VGND.n2201 VGND.n1713 76.3222
R2295 VGND.n2216 VGND.n2215 76.3222
R2296 VGND.n2217 VGND.n1708 76.3222
R2297 VGND.n2231 VGND.n2230 76.3222
R2298 VGND.n2232 VGND.n1701 76.3222
R2299 VGND.n2246 VGND.n2245 76.3222
R2300 VGND.n2072 VGND.n1968 76.3222
R2301 VGND.n2079 VGND.n2078 76.3222
R2302 VGND.n2080 VGND.n1966 76.3222
R2303 VGND.n2087 VGND.n2086 76.3222
R2304 VGND.n2088 VGND.n1964 76.3222
R2305 VGND.n1331 VGND.n1330 76.3222
R2306 VGND.n1332 VGND.n1306 76.3222
R2307 VGND.n1339 VGND.n1338 76.3222
R2308 VGND.n1340 VGND.n1304 76.3222
R2309 VGND.n1347 VGND.n1346 76.3222
R2310 VGND.n1044 VGND.n1043 76.3222
R2311 VGND.n1046 VGND.n437 76.3222
R2312 VGND.n1053 VGND.n1052 76.3222
R2313 VGND.n1054 VGND.n435 76.3222
R2314 VGND.n1061 VGND.n1060 76.3222
R2315 VGND.t93 VGND.t7 74.8304
R2316 VGND.t173 VGND.t160 74.8304
R2317 VGND.t3 VGND.t212 74.8304
R2318 VGND.n1927 VGND.n1910 74.5978
R2319 VGND.n1928 VGND.n1927 74.5978
R2320 VGND.n1848 VGND.n1831 74.5978
R2321 VGND.n1849 VGND.n1848 74.5978
R2322 VGND.n318 VGND.n317 74.5978
R2323 VGND.n317 VGND.n316 74.5978
R2324 VGND.n399 VGND.n368 74.5978
R2325 VGND.n396 VGND.n368 74.5978
R2326 VGND.n1509 VGND.n1492 74.5978
R2327 VGND.n1510 VGND.n1509 74.5978
R2328 VGND.n1247 VGND.n1195 74.5978
R2329 VGND.n1244 VGND.n1195 74.5978
R2330 VGND.n1419 VGND.n1365 74.5978
R2331 VGND.n1416 VGND.n1365 74.5978
R2332 VGND.n1740 VGND.n1723 74.5978
R2333 VGND.n1741 VGND.n1740 74.5978
R2334 VGND.n223 VGND.n164 74.5978
R2335 VGND.n220 VGND.n164 74.5978
R2336 VGND.n711 VGND.n7 74.09
R2337 VGND.n721 VGND.n720 74.09
R2338 VGND.n723 VGND.n668 74.09
R2339 VGND.n727 VGND.n726 74.09
R2340 VGND.n729 VGND.n728 74.09
R2341 VGND.n708 VGND.n10 74.09
R2342 VGND.n698 VGND.n697 74.09
R2343 VGND.n694 VGND.n674 74.09
R2344 VGND.n692 VGND.n691 74.09
R2345 VGND.n690 VGND.n689 74.09
R2346 VGND.n736 VGND.n735 73.9572
R2347 VGND.n679 VGND.n677 73.8434
R2348 VGND.n731 VGND.n667 73.3478
R2349 VGND.n735 VGND.n734 73.3478
R2350 VGND.n680 VGND.n679 72.7809
R2351 VGND.n683 VGND.n675 72.7809
R2352 VGND.n662 VGND.n661 71.4976
R2353 VGND.t193 VGND.n46 70.6648
R2354 VGND.n688 VGND.n685 70.12
R2355 VGND.t201 VGND.t83 69.8418
R2356 VGND.n576 VGND.n461 69.4466
R2357 VGND.n2105 VGND.n2104 69.3109
R2358 VGND.n2104 VGND.n2103 69.3109
R2359 VGND.n2154 VGND.n2153 69.3109
R2360 VGND.n2153 VGND.n2152 69.3109
R2361 VGND.n1122 VGND.n289 69.3109
R2362 VGND.n351 VGND.n289 69.3109
R2363 VGND.n1095 VGND.n1094 69.3109
R2364 VGND.n1095 VGND.n380 69.3109
R2365 VGND.n1550 VGND.n1549 69.3109
R2366 VGND.n1549 VGND.n1548 69.3109
R2367 VGND.n1290 VGND.n1185 69.3109
R2368 VGND.n1266 VGND.n1185 69.3109
R2369 VGND.n1461 VGND.n1355 69.3109
R2370 VGND.n1437 VGND.n1355 69.3109
R2371 VGND.n2209 VGND.n2208 69.3109
R2372 VGND.n2208 VGND.n2207 69.3109
R2373 VGND.n259 VGND.n157 69.3109
R2374 VGND.n259 VGND.n258 69.3109
R2375 VGND.n717 VGND.n716 68.2005
R2376 VGND.n714 VGND.n671 68.2005
R2377 VGND.n701 VGND.n673 68.2005
R2378 VGND.n705 VGND.n704 68.2005
R2379 VGND.n947 VGND.n946 68.2005
R2380 VGND.n926 VGND.n925 68.2005
R2381 VGND.n864 VGND.n863 66.5605
R2382 VGND.n863 VGND.n743 66.5605
R2383 VGND.n1949 VGND.t194 65.8183
R2384 VGND.n1951 VGND.t194 65.8183
R2385 VGND.n1957 VGND.t194 65.8183
R2386 VGND.n1959 VGND.t194 65.8183
R2387 VGND.n1933 VGND.t194 65.8183
R2388 VGND.n1935 VGND.t194 65.8183
R2389 VGND.n1941 VGND.t194 65.8183
R2390 VGND.n1943 VGND.t194 65.8183
R2391 VGND.t194 VGND.n1891 65.8183
R2392 VGND.n1918 VGND.t194 65.8183
R2393 VGND.n1914 VGND.t194 65.8183
R2394 VGND.n1925 VGND.t194 65.8183
R2395 VGND.n2134 VGND.t194 65.8183
R2396 VGND.n2121 VGND.t194 65.8183
R2397 VGND.n2119 VGND.t194 65.8183
R2398 VGND.n2106 VGND.t194 65.8183
R2399 VGND.n1870 VGND.t235 65.8183
R2400 VGND.n1872 VGND.t235 65.8183
R2401 VGND.n1878 VGND.t235 65.8183
R2402 VGND.n1880 VGND.t235 65.8183
R2403 VGND.n1854 VGND.t235 65.8183
R2404 VGND.n1856 VGND.t235 65.8183
R2405 VGND.n1862 VGND.t235 65.8183
R2406 VGND.n1864 VGND.t235 65.8183
R2407 VGND.t235 VGND.n1812 65.8183
R2408 VGND.n1839 VGND.t235 65.8183
R2409 VGND.n1835 VGND.t235 65.8183
R2410 VGND.n1846 VGND.t235 65.8183
R2411 VGND.n2183 VGND.t235 65.8183
R2412 VGND.n2170 VGND.t235 65.8183
R2413 VGND.n2168 VGND.t235 65.8183
R2414 VGND.n2155 VGND.t235 65.8183
R2415 VGND.n335 VGND.t218 65.8183
R2416 VGND.n341 VGND.t218 65.8183
R2417 VGND.n343 VGND.t218 65.8183
R2418 VGND.n349 VGND.t218 65.8183
R2419 VGND.n319 VGND.t218 65.8183
R2420 VGND.n325 VGND.t218 65.8183
R2421 VGND.n327 VGND.t218 65.8183
R2422 VGND.n333 VGND.t218 65.8183
R2423 VGND.t218 VGND.n281 65.8183
R2424 VGND.n303 VGND.t218 65.8183
R2425 VGND.n310 VGND.t218 65.8183
R2426 VGND.n301 VGND.t218 65.8183
R2427 VGND.n1147 VGND.t218 65.8183
R2428 VGND.n1137 VGND.t218 65.8183
R2429 VGND.n1135 VGND.t218 65.8183
R2430 VGND.n1123 VGND.t218 65.8183
R2431 VGND.t199 VGND.n379 65.8183
R2432 VGND.t199 VGND.n378 65.8183
R2433 VGND.t199 VGND.n377 65.8183
R2434 VGND.t199 VGND.n376 65.8183
R2435 VGND.t199 VGND.n367 65.8183
R2436 VGND.t199 VGND.n374 65.8183
R2437 VGND.t199 VGND.n364 65.8183
R2438 VGND.t199 VGND.n375 65.8183
R2439 VGND.t199 VGND.n373 65.8183
R2440 VGND.t199 VGND.n371 65.8183
R2441 VGND.t199 VGND.n370 65.8183
R2442 VGND.t199 VGND.n369 65.8183
R2443 VGND.n1096 VGND.t199 65.8183
R2444 VGND.t199 VGND.n366 65.8183
R2445 VGND.t199 VGND.n365 65.8183
R2446 VGND.t199 VGND.n363 65.8183
R2447 VGND.n1531 VGND.t230 65.8183
R2448 VGND.n1533 VGND.t230 65.8183
R2449 VGND.n1539 VGND.t230 65.8183
R2450 VGND.n1541 VGND.t230 65.8183
R2451 VGND.n1515 VGND.t230 65.8183
R2452 VGND.n1517 VGND.t230 65.8183
R2453 VGND.n1523 VGND.t230 65.8183
R2454 VGND.n1525 VGND.t230 65.8183
R2455 VGND.t230 VGND.n1472 65.8183
R2456 VGND.n1500 VGND.t230 65.8183
R2457 VGND.n1496 VGND.t230 65.8183
R2458 VGND.n1507 VGND.t230 65.8183
R2459 VGND.n1579 VGND.t230 65.8183
R2460 VGND.n1566 VGND.t230 65.8183
R2461 VGND.n1564 VGND.t230 65.8183
R2462 VGND.n1551 VGND.t230 65.8183
R2463 VGND.t227 VGND.n1280 65.8183
R2464 VGND.t227 VGND.n1204 65.8183
R2465 VGND.t227 VGND.n1203 65.8183
R2466 VGND.t227 VGND.n1202 65.8183
R2467 VGND.t227 VGND.n1193 65.8183
R2468 VGND.t227 VGND.n1200 65.8183
R2469 VGND.t227 VGND.n1191 65.8183
R2470 VGND.t227 VGND.n1201 65.8183
R2471 VGND.t227 VGND.n1199 65.8183
R2472 VGND.t227 VGND.n1198 65.8183
R2473 VGND.t227 VGND.n1197 65.8183
R2474 VGND.t227 VGND.n1196 65.8183
R2475 VGND.t227 VGND.n1194 65.8183
R2476 VGND.t227 VGND.n1192 65.8183
R2477 VGND.n1281 VGND.t227 65.8183
R2478 VGND.t227 VGND.n1186 65.8183
R2479 VGND.t192 VGND.n1451 65.8183
R2480 VGND.t192 VGND.n1374 65.8183
R2481 VGND.t192 VGND.n1373 65.8183
R2482 VGND.t192 VGND.n1372 65.8183
R2483 VGND.t192 VGND.n1363 65.8183
R2484 VGND.t192 VGND.n1370 65.8183
R2485 VGND.t192 VGND.n1361 65.8183
R2486 VGND.t192 VGND.n1371 65.8183
R2487 VGND.t192 VGND.n1369 65.8183
R2488 VGND.t192 VGND.n1368 65.8183
R2489 VGND.t192 VGND.n1367 65.8183
R2490 VGND.t192 VGND.n1366 65.8183
R2491 VGND.t192 VGND.n1364 65.8183
R2492 VGND.t192 VGND.n1362 65.8183
R2493 VGND.n1452 VGND.t192 65.8183
R2494 VGND.t192 VGND.n1356 65.8183
R2495 VGND.n1762 VGND.t195 65.8183
R2496 VGND.n1764 VGND.t195 65.8183
R2497 VGND.n1770 VGND.t195 65.8183
R2498 VGND.n1772 VGND.t195 65.8183
R2499 VGND.n1746 VGND.t195 65.8183
R2500 VGND.n1748 VGND.t195 65.8183
R2501 VGND.n1754 VGND.t195 65.8183
R2502 VGND.n1756 VGND.t195 65.8183
R2503 VGND.t195 VGND.n1704 65.8183
R2504 VGND.n1731 VGND.t195 65.8183
R2505 VGND.n1727 VGND.t195 65.8183
R2506 VGND.n1738 VGND.t195 65.8183
R2507 VGND.n2238 VGND.t195 65.8183
R2508 VGND.n2225 VGND.t195 65.8183
R2509 VGND.n2223 VGND.t195 65.8183
R2510 VGND.n2210 VGND.t195 65.8183
R2511 VGND.t231 VGND.n174 65.8183
R2512 VGND.t231 VGND.n173 65.8183
R2513 VGND.t231 VGND.n172 65.8183
R2514 VGND.t231 VGND.n171 65.8183
R2515 VGND.t231 VGND.n162 65.8183
R2516 VGND.t231 VGND.n169 65.8183
R2517 VGND.t231 VGND.n159 65.8183
R2518 VGND.t231 VGND.n170 65.8183
R2519 VGND.t231 VGND.n168 65.8183
R2520 VGND.t231 VGND.n167 65.8183
R2521 VGND.t231 VGND.n166 65.8183
R2522 VGND.t231 VGND.n165 65.8183
R2523 VGND.t231 VGND.n163 65.8183
R2524 VGND.t231 VGND.n161 65.8183
R2525 VGND.t231 VGND.n160 65.8183
R2526 VGND.n260 VGND.t231 65.8183
R2527 VGND.t241 VGND.t201 64.8531
R2528 VGND.t258 VGND.t241 64.8531
R2529 VGND.t111 VGND.t258 64.8531
R2530 VGND.n1610 VGND.t27 63.9747
R2531 VGND.t193 VGND.n38 60.9488
R2532 VGND.t193 VGND.n42 60.9488
R2533 VGND.n748 VGND.t136 60.0005
R2534 VGND.n748 VGND.t174 60.0005
R2535 VGND.n747 VGND.t242 60.0005
R2536 VGND.n747 VGND.t112 60.0005
R2537 VGND.n749 VGND.t186 60.0005
R2538 VGND.n749 VGND.t213 60.0005
R2539 VGND.n741 VGND.t10 60.0005
R2540 VGND.n741 VGND.t76 60.0005
R2541 VGND.n740 VGND.t229 60.0005
R2542 VGND.n740 VGND.t163 60.0005
R2543 VGND.n742 VGND.t126 60.0005
R2544 VGND.n742 VGND.t238 60.0005
R2545 VGND.n843 VGND.n760 59.0609
R2546 VGND.n2104 VGND.t194 57.8461
R2547 VGND.n2153 VGND.t235 57.8461
R2548 VGND.n289 VGND.t218 57.8461
R2549 VGND.t199 VGND.n1095 57.8461
R2550 VGND.n1549 VGND.t230 57.8461
R2551 VGND.t227 VGND.n1185 57.8461
R2552 VGND.t192 VGND.n1355 57.8461
R2553 VGND.n2208 VGND.t195 57.8461
R2554 VGND.t231 VGND.n259 57.8461
R2555 VGND.t193 VGND.n43 57.0946
R2556 VGND.n1063 VGND.n1062 56.3995
R2557 VGND.n1064 VGND.n1063 56.3995
R2558 VGND.n2095 VGND.n2094 56.3995
R2559 VGND.n2349 VGND.n2348 56.3995
R2560 VGND.n1589 VGND.n1173 56.3995
R2561 VGND.n2251 VGND.n2250 56.3995
R2562 VGND.n2251 VGND.n2247 56.3995
R2563 VGND.n1589 VGND.n1588 56.3995
R2564 VGND.n2348 VGND.n20 56.3995
R2565 VGND.n2096 VGND.n2095 56.3995
R2566 VGND.n1350 VGND.n1301 56.3995
R2567 VGND.n853 VGND.n852 55.4005
R2568 VGND.n1927 VGND.t194 55.2026
R2569 VGND.n1848 VGND.t235 55.2026
R2570 VGND.n317 VGND.t218 55.2026
R2571 VGND.t199 VGND.n368 55.2026
R2572 VGND.n1509 VGND.t230 55.2026
R2573 VGND.t227 VGND.n1195 55.2026
R2574 VGND.t192 VGND.n1365 55.2026
R2575 VGND.n1740 VGND.t195 55.2026
R2576 VGND.t231 VGND.n164 55.2026
R2577 VGND.t7 VGND.t150 54.8758
R2578 VGND.t160 VGND.t185 54.8758
R2579 VGND.t185 VGND.t3 54.8758
R2580 VGND.n828 VGND.n827 53.5422
R2581 VGND.n826 VGND.n825 53.5422
R2582 VGND.n805 VGND.n804 53.5422
R2583 VGND.n803 VGND.n802 53.5422
R2584 VGND.n785 VGND.n784 53.5422
R2585 VGND.n783 VGND.n782 53.5422
R2586 VGND.n1943 VGND.n1906 53.3664
R2587 VGND.n1942 VGND.n1941 53.3664
R2588 VGND.n1935 VGND.n1908 53.3664
R2589 VGND.n1934 VGND.n1933 53.3664
R2590 VGND.n1925 VGND.n1924 53.3664
R2591 VGND.n1920 VGND.n1914 53.3664
R2592 VGND.n1918 VGND.n1917 53.3664
R2593 VGND.n2136 VGND.n1891 53.3664
R2594 VGND.n2107 VGND.n2106 53.3664
R2595 VGND.n2119 VGND.n2118 53.3664
R2596 VGND.n2122 VGND.n2121 53.3664
R2597 VGND.n2134 VGND.n2133 53.3664
R2598 VGND.n1950 VGND.n1949 53.3664
R2599 VGND.n1952 VGND.n1951 53.3664
R2600 VGND.n1957 VGND.n1956 53.3664
R2601 VGND.n1960 VGND.n1959 53.3664
R2602 VGND.n1949 VGND.n1948 53.3664
R2603 VGND.n1951 VGND.n1904 53.3664
R2604 VGND.n1958 VGND.n1957 53.3664
R2605 VGND.n1959 VGND.n1902 53.3664
R2606 VGND.n1933 VGND.n1932 53.3664
R2607 VGND.n1936 VGND.n1935 53.3664
R2608 VGND.n1941 VGND.n1940 53.3664
R2609 VGND.n1944 VGND.n1943 53.3664
R2610 VGND.n1915 VGND.n1891 53.3664
R2611 VGND.n1919 VGND.n1918 53.3664
R2612 VGND.n1914 VGND.n1912 53.3664
R2613 VGND.n1926 VGND.n1925 53.3664
R2614 VGND.n2135 VGND.n2134 53.3664
R2615 VGND.n2121 VGND.n1892 53.3664
R2616 VGND.n2120 VGND.n2119 53.3664
R2617 VGND.n2106 VGND.n1897 53.3664
R2618 VGND.n1864 VGND.n1827 53.3664
R2619 VGND.n1863 VGND.n1862 53.3664
R2620 VGND.n1856 VGND.n1829 53.3664
R2621 VGND.n1855 VGND.n1854 53.3664
R2622 VGND.n1846 VGND.n1845 53.3664
R2623 VGND.n1841 VGND.n1835 53.3664
R2624 VGND.n1839 VGND.n1838 53.3664
R2625 VGND.n2185 VGND.n1812 53.3664
R2626 VGND.n2156 VGND.n2155 53.3664
R2627 VGND.n2168 VGND.n2167 53.3664
R2628 VGND.n2171 VGND.n2170 53.3664
R2629 VGND.n2183 VGND.n2182 53.3664
R2630 VGND.n1871 VGND.n1870 53.3664
R2631 VGND.n1873 VGND.n1872 53.3664
R2632 VGND.n1878 VGND.n1877 53.3664
R2633 VGND.n1881 VGND.n1880 53.3664
R2634 VGND.n1870 VGND.n1869 53.3664
R2635 VGND.n1872 VGND.n1825 53.3664
R2636 VGND.n1879 VGND.n1878 53.3664
R2637 VGND.n1880 VGND.n1823 53.3664
R2638 VGND.n1854 VGND.n1853 53.3664
R2639 VGND.n1857 VGND.n1856 53.3664
R2640 VGND.n1862 VGND.n1861 53.3664
R2641 VGND.n1865 VGND.n1864 53.3664
R2642 VGND.n1836 VGND.n1812 53.3664
R2643 VGND.n1840 VGND.n1839 53.3664
R2644 VGND.n1835 VGND.n1833 53.3664
R2645 VGND.n1847 VGND.n1846 53.3664
R2646 VGND.n2184 VGND.n2183 53.3664
R2647 VGND.n2170 VGND.n1813 53.3664
R2648 VGND.n2169 VGND.n2168 53.3664
R2649 VGND.n2155 VGND.n1818 53.3664
R2650 VGND.n334 VGND.n333 53.3664
R2651 VGND.n327 VGND.n295 53.3664
R2652 VGND.n326 VGND.n325 53.3664
R2653 VGND.n319 VGND.n297 53.3664
R2654 VGND.n312 VGND.n301 53.3664
R2655 VGND.n310 VGND.n309 53.3664
R2656 VGND.n305 VGND.n303 53.3664
R2657 VGND.n1149 VGND.n281 53.3664
R2658 VGND.n1124 VGND.n1123 53.3664
R2659 VGND.n1135 VGND.n1134 53.3664
R2660 VGND.n1138 VGND.n1137 53.3664
R2661 VGND.n1147 VGND.n1146 53.3664
R2662 VGND.n335 VGND.n293 53.3664
R2663 VGND.n341 VGND.n340 53.3664
R2664 VGND.n344 VGND.n343 53.3664
R2665 VGND.n349 VGND.n348 53.3664
R2666 VGND.n336 VGND.n335 53.3664
R2667 VGND.n342 VGND.n341 53.3664
R2668 VGND.n343 VGND.n291 53.3664
R2669 VGND.n350 VGND.n349 53.3664
R2670 VGND.n320 VGND.n319 53.3664
R2671 VGND.n325 VGND.n324 53.3664
R2672 VGND.n328 VGND.n327 53.3664
R2673 VGND.n333 VGND.n332 53.3664
R2674 VGND.n304 VGND.n281 53.3664
R2675 VGND.n303 VGND.n302 53.3664
R2676 VGND.n311 VGND.n310 53.3664
R2677 VGND.n301 VGND.n299 53.3664
R2678 VGND.n1148 VGND.n1147 53.3664
R2679 VGND.n1137 VGND.n282 53.3664
R2680 VGND.n1136 VGND.n1135 53.3664
R2681 VGND.n1123 VGND.n286 53.3664
R2682 VGND.n415 VGND.n375 53.3664
R2683 VGND.n411 VGND.n364 53.3664
R2684 VGND.n407 VGND.n374 53.3664
R2685 VGND.n403 VGND.n367 53.3664
R2686 VGND.n392 VGND.n369 53.3664
R2687 VGND.n388 VGND.n370 53.3664
R2688 VGND.n384 VGND.n371 53.3664
R2689 VGND.n373 VGND.n372 53.3664
R2690 VGND.n381 VGND.n363 53.3664
R2691 VGND.n1083 VGND.n365 53.3664
R2692 VGND.n1076 VGND.n366 53.3664
R2693 VGND.n1097 VGND.n1096 53.3664
R2694 VGND.n419 VGND.n379 53.3664
R2695 VGND.n420 VGND.n378 53.3664
R2696 VGND.n424 VGND.n377 53.3664
R2697 VGND.n428 VGND.n376 53.3664
R2698 VGND.n416 VGND.n379 53.3664
R2699 VGND.n423 VGND.n378 53.3664
R2700 VGND.n427 VGND.n377 53.3664
R2701 VGND.n430 VGND.n376 53.3664
R2702 VGND.n400 VGND.n367 53.3664
R2703 VGND.n404 VGND.n374 53.3664
R2704 VGND.n408 VGND.n364 53.3664
R2705 VGND.n412 VGND.n375 53.3664
R2706 VGND.n383 VGND.n373 53.3664
R2707 VGND.n387 VGND.n371 53.3664
R2708 VGND.n391 VGND.n370 53.3664
R2709 VGND.n395 VGND.n369 53.3664
R2710 VGND.n1096 VGND.n362 53.3664
R2711 VGND.n366 VGND.n361 53.3664
R2712 VGND.n1075 VGND.n365 53.3664
R2713 VGND.n1082 VGND.n363 53.3664
R2714 VGND.n1525 VGND.n1488 53.3664
R2715 VGND.n1524 VGND.n1523 53.3664
R2716 VGND.n1517 VGND.n1490 53.3664
R2717 VGND.n1516 VGND.n1515 53.3664
R2718 VGND.n1507 VGND.n1506 53.3664
R2719 VGND.n1502 VGND.n1496 53.3664
R2720 VGND.n1500 VGND.n1499 53.3664
R2721 VGND.n1581 VGND.n1472 53.3664
R2722 VGND.n1552 VGND.n1551 53.3664
R2723 VGND.n1564 VGND.n1563 53.3664
R2724 VGND.n1567 VGND.n1566 53.3664
R2725 VGND.n1579 VGND.n1578 53.3664
R2726 VGND.n1532 VGND.n1531 53.3664
R2727 VGND.n1534 VGND.n1533 53.3664
R2728 VGND.n1539 VGND.n1538 53.3664
R2729 VGND.n1542 VGND.n1541 53.3664
R2730 VGND.n1531 VGND.n1530 53.3664
R2731 VGND.n1533 VGND.n1486 53.3664
R2732 VGND.n1540 VGND.n1539 53.3664
R2733 VGND.n1541 VGND.n1484 53.3664
R2734 VGND.n1515 VGND.n1514 53.3664
R2735 VGND.n1518 VGND.n1517 53.3664
R2736 VGND.n1523 VGND.n1522 53.3664
R2737 VGND.n1526 VGND.n1525 53.3664
R2738 VGND.n1497 VGND.n1472 53.3664
R2739 VGND.n1501 VGND.n1500 53.3664
R2740 VGND.n1496 VGND.n1494 53.3664
R2741 VGND.n1508 VGND.n1507 53.3664
R2742 VGND.n1580 VGND.n1579 53.3664
R2743 VGND.n1566 VGND.n1473 53.3664
R2744 VGND.n1565 VGND.n1564 53.3664
R2745 VGND.n1551 VGND.n1478 53.3664
R2746 VGND.n1262 VGND.n1201 53.3664
R2747 VGND.n1259 VGND.n1191 53.3664
R2748 VGND.n1255 VGND.n1200 53.3664
R2749 VGND.n1251 VGND.n1193 53.3664
R2750 VGND.n1240 VGND.n1196 53.3664
R2751 VGND.n1236 VGND.n1197 53.3664
R2752 VGND.n1232 VGND.n1198 53.3664
R2753 VGND.n1228 VGND.n1199 53.3664
R2754 VGND.n1289 VGND.n1186 53.3664
R2755 VGND.n1282 VGND.n1281 53.3664
R2756 VGND.n1213 VGND.n1192 53.3664
R2757 VGND.n1220 VGND.n1194 53.3664
R2758 VGND.n1280 VGND.n1279 53.3664
R2759 VGND.n1206 VGND.n1204 53.3664
R2760 VGND.n1274 VGND.n1203 53.3664
R2761 VGND.n1270 VGND.n1202 53.3664
R2762 VGND.n1280 VGND.n1205 53.3664
R2763 VGND.n1275 VGND.n1204 53.3664
R2764 VGND.n1271 VGND.n1203 53.3664
R2765 VGND.n1267 VGND.n1202 53.3664
R2766 VGND.n1248 VGND.n1193 53.3664
R2767 VGND.n1252 VGND.n1200 53.3664
R2768 VGND.n1256 VGND.n1191 53.3664
R2769 VGND.n1260 VGND.n1201 53.3664
R2770 VGND.n1231 VGND.n1199 53.3664
R2771 VGND.n1235 VGND.n1198 53.3664
R2772 VGND.n1239 VGND.n1197 53.3664
R2773 VGND.n1243 VGND.n1196 53.3664
R2774 VGND.n1227 VGND.n1194 53.3664
R2775 VGND.n1219 VGND.n1192 53.3664
R2776 VGND.n1281 VGND.n1190 53.3664
R2777 VGND.n1189 VGND.n1186 53.3664
R2778 VGND.n1434 VGND.n1371 53.3664
R2779 VGND.n1431 VGND.n1361 53.3664
R2780 VGND.n1427 VGND.n1370 53.3664
R2781 VGND.n1423 VGND.n1363 53.3664
R2782 VGND.n1412 VGND.n1366 53.3664
R2783 VGND.n1408 VGND.n1367 53.3664
R2784 VGND.n1404 VGND.n1368 53.3664
R2785 VGND.n1400 VGND.n1369 53.3664
R2786 VGND.n1460 VGND.n1356 53.3664
R2787 VGND.n1453 VGND.n1452 53.3664
R2788 VGND.n1385 VGND.n1362 53.3664
R2789 VGND.n1392 VGND.n1364 53.3664
R2790 VGND.n1451 VGND.n1450 53.3664
R2791 VGND.n1376 VGND.n1374 53.3664
R2792 VGND.n1445 VGND.n1373 53.3664
R2793 VGND.n1441 VGND.n1372 53.3664
R2794 VGND.n1451 VGND.n1375 53.3664
R2795 VGND.n1446 VGND.n1374 53.3664
R2796 VGND.n1442 VGND.n1373 53.3664
R2797 VGND.n1438 VGND.n1372 53.3664
R2798 VGND.n1420 VGND.n1363 53.3664
R2799 VGND.n1424 VGND.n1370 53.3664
R2800 VGND.n1428 VGND.n1361 53.3664
R2801 VGND.n1432 VGND.n1371 53.3664
R2802 VGND.n1403 VGND.n1369 53.3664
R2803 VGND.n1407 VGND.n1368 53.3664
R2804 VGND.n1411 VGND.n1367 53.3664
R2805 VGND.n1415 VGND.n1366 53.3664
R2806 VGND.n1399 VGND.n1364 53.3664
R2807 VGND.n1391 VGND.n1362 53.3664
R2808 VGND.n1452 VGND.n1360 53.3664
R2809 VGND.n1359 VGND.n1356 53.3664
R2810 VGND.n1756 VGND.n1719 53.3664
R2811 VGND.n1755 VGND.n1754 53.3664
R2812 VGND.n1748 VGND.n1721 53.3664
R2813 VGND.n1747 VGND.n1746 53.3664
R2814 VGND.n1738 VGND.n1737 53.3664
R2815 VGND.n1733 VGND.n1727 53.3664
R2816 VGND.n1731 VGND.n1730 53.3664
R2817 VGND.n2240 VGND.n1704 53.3664
R2818 VGND.n2211 VGND.n2210 53.3664
R2819 VGND.n2223 VGND.n2222 53.3664
R2820 VGND.n2226 VGND.n2225 53.3664
R2821 VGND.n2238 VGND.n2237 53.3664
R2822 VGND.n1763 VGND.n1762 53.3664
R2823 VGND.n1765 VGND.n1764 53.3664
R2824 VGND.n1770 VGND.n1769 53.3664
R2825 VGND.n1773 VGND.n1772 53.3664
R2826 VGND.n1762 VGND.n1761 53.3664
R2827 VGND.n1764 VGND.n1717 53.3664
R2828 VGND.n1771 VGND.n1770 53.3664
R2829 VGND.n1772 VGND.n1715 53.3664
R2830 VGND.n1746 VGND.n1745 53.3664
R2831 VGND.n1749 VGND.n1748 53.3664
R2832 VGND.n1754 VGND.n1753 53.3664
R2833 VGND.n1757 VGND.n1756 53.3664
R2834 VGND.n1728 VGND.n1704 53.3664
R2835 VGND.n1732 VGND.n1731 53.3664
R2836 VGND.n1727 VGND.n1725 53.3664
R2837 VGND.n1739 VGND.n1738 53.3664
R2838 VGND.n2239 VGND.n2238 53.3664
R2839 VGND.n2225 VGND.n1705 53.3664
R2840 VGND.n2224 VGND.n2223 53.3664
R2841 VGND.n2210 VGND.n1710 53.3664
R2842 VGND.n239 VGND.n170 53.3664
R2843 VGND.n235 VGND.n159 53.3664
R2844 VGND.n231 VGND.n169 53.3664
R2845 VGND.n227 VGND.n162 53.3664
R2846 VGND.n216 VGND.n165 53.3664
R2847 VGND.n212 VGND.n166 53.3664
R2848 VGND.n208 VGND.n167 53.3664
R2849 VGND.n204 VGND.n168 53.3664
R2850 VGND.n261 VGND.n260 53.3664
R2851 VGND.n182 VGND.n160 53.3664
R2852 VGND.n189 VGND.n161 53.3664
R2853 VGND.n196 VGND.n163 53.3664
R2854 VGND.n243 VGND.n174 53.3664
R2855 VGND.n244 VGND.n173 53.3664
R2856 VGND.n248 VGND.n172 53.3664
R2857 VGND.n252 VGND.n171 53.3664
R2858 VGND.n240 VGND.n174 53.3664
R2859 VGND.n247 VGND.n173 53.3664
R2860 VGND.n251 VGND.n172 53.3664
R2861 VGND.n175 VGND.n171 53.3664
R2862 VGND.n224 VGND.n162 53.3664
R2863 VGND.n228 VGND.n169 53.3664
R2864 VGND.n232 VGND.n159 53.3664
R2865 VGND.n236 VGND.n170 53.3664
R2866 VGND.n207 VGND.n168 53.3664
R2867 VGND.n211 VGND.n167 53.3664
R2868 VGND.n215 VGND.n166 53.3664
R2869 VGND.n219 VGND.n165 53.3664
R2870 VGND.n203 VGND.n163 53.3664
R2871 VGND.n195 VGND.n161 53.3664
R2872 VGND.n188 VGND.n160 53.3664
R2873 VGND.n260 VGND.n158 53.3664
R2874 VGND.n863 VGND.n862 53.3255
R2875 VGND.t69 VGND.t264 49.8871
R2876 VGND.n846 VGND.n759 49.8871
R2877 VGND.t46 VGND.n880 49.3595
R2878 VGND.n3 VGND.t167 48.0005
R2879 VGND.n3 VGND.t247 48.0005
R2880 VGND.n933 VGND.t191 48.0005
R2881 VGND.n933 VGND.t106 48.0005
R2882 VGND.n936 VGND.t119 48.0005
R2883 VGND.n936 VGND.t132 48.0005
R2884 VGND.n938 VGND.t26 48.0005
R2885 VGND.n938 VGND.t72 48.0005
R2886 VGND.n940 VGND.t158 48.0005
R2887 VGND.n940 VGND.t66 48.0005
R2888 VGND.n942 VGND.t45 48.0005
R2889 VGND.n942 VGND.t68 48.0005
R2890 VGND.n944 VGND.t101 48.0005
R2891 VGND.n944 VGND.t284 48.0005
R2892 VGND.n929 VGND.t267 48.0005
R2893 VGND.n929 VGND.t122 48.0005
R2894 VGND.n927 VGND.t292 48.0005
R2895 VGND.n927 VGND.t255 48.0005
R2896 VGND.n663 VGND.t290 48.0005
R2897 VGND.n663 VGND.t178 48.0005
R2898 VGND.n918 VGND.t279 48.0005
R2899 VGND.n918 VGND.t14 48.0005
R2900 VGND.n920 VGND.t97 48.0005
R2901 VGND.n920 VGND.t24 48.0005
R2902 VGND.n916 VGND.t80 48.0005
R2903 VGND.n916 VGND.t6 48.0005
R2904 VGND.n914 VGND.t78 48.0005
R2905 VGND.n914 VGND.t108 48.0005
R2906 VGND.n912 VGND.t134 48.0005
R2907 VGND.n912 VGND.t145 48.0005
R2908 VGND.n665 VGND.t140 48.0005
R2909 VGND.n665 VGND.t277 48.0005
R2910 VGND.n904 VGND.t142 48.0005
R2911 VGND.n904 VGND.t147 48.0005
R2912 VGND.n906 VGND.t299 48.0005
R2913 VGND.n906 VGND.t110 48.0005
R2914 VGND.n902 VGND.t249 48.0005
R2915 VGND.n902 VGND.t257 48.0005
R2916 VGND.n900 VGND.t154 48.0005
R2917 VGND.n900 VGND.t130 48.0005
R2918 VGND.n899 VGND.t42 48.0005
R2919 VGND.n899 VGND.t38 48.0005
R2920 VGND.t193 VGND.n45 46.4131
R2921 VGND.t233 VGND.t125 44.8985
R2922 VGND.t237 VGND.t15 44.8985
R2923 VGND.n846 VGND.n845 39.9098
R2924 VGND.n492 VGND.n491 37.6324
R2925 VGND.n491 VGND.n490 37.6324
R2926 VGND.n490 VGND.n485 37.6324
R2927 VGND.n485 VGND.n28 37.6324
R2928 VGND.n2335 VGND.n28 37.6324
R2929 VGND.n2341 VGND.n24 37.6324
R2930 VGND.n2342 VGND.n2341 37.6324
R2931 VGND.n2343 VGND.n2342 37.6324
R2932 VGND.n2343 VGND.n17 37.6324
R2933 VGND.n2350 VGND.n18 37.6324
R2934 VGND.n1610 VGND.n1609 37.6324
R2935 VGND.n1609 VGND.n1608 37.6324
R2936 VGND.n1608 VGND.n1164 37.6324
R2937 VGND.n1602 VGND.n1164 37.6324
R2938 VGND.n1602 VGND.n49 37.6324
R2939 VGND.n1171 VGND.n48 37.6324
R2940 VGND.n1595 VGND.n1171 37.6324
R2941 VGND.n1595 VGND.n1594 37.6324
R2942 VGND.n1594 VGND.n1593 37.6324
R2943 VGND.n1593 VGND.n1172 37.6324
R2944 VGND.n1172 VGND.n45 37.6324
R2945 VGND.n2268 VGND.n46 37.6324
R2946 VGND.n2268 VGND.n2267 37.6324
R2947 VGND.n2267 VGND.n2266 37.6324
R2948 VGND.n2266 VGND.n1690 37.6324
R2949 VGND.n1690 VGND.n40 37.6324
R2950 VGND.n2258 VGND.n41 37.6324
R2951 VGND.n2258 VGND.n2257 37.6324
R2952 VGND.n2257 VGND.n2256 37.6324
R2953 VGND.n2256 VGND.n1696 37.6324
R2954 VGND.n2249 VGND.n1696 37.6324
R2955 VGND.n2249 VGND.n2248 37.6324
R2956 VGND.t216 VGND.t173 34.9211
R2957 VGND.t86 VGND.n959 33.8062
R2958 VGND.n656 VGND.n634 33.0531
R2959 VGND.n2351 VGND.n2350 33.0329
R2960 VGND.t193 VGND.n47 32.9056
R2961 VGND.t143 VGND.t95 32.6148
R2962 VGND.n641 VGND.n580 32.3969
R2963 VGND.t193 VGND.n36 31.5314
R2964 VGND.n566 VGND.n467 31.5314
R2965 VGND.t193 VGND.n35 30.857
R2966 VGND.n516 VGND.n467 30.857
R2967 VGND.n858 VGND.t285 29.9325
R2968 VGND.t81 VGND.t252 29.9325
R2969 VGND.n857 VGND.t83 29.9325
R2970 VGND.n1947 VGND.n1946 27.5561
R2971 VGND.n1868 VGND.n1867 27.5561
R2972 VGND.n337 VGND.n294 27.5561
R2973 VGND.n417 VGND.n414 27.5561
R2974 VGND.n1529 VGND.n1528 27.5561
R2975 VGND.n1264 VGND.n1263 27.5561
R2976 VGND.n1436 VGND.n1435 27.5561
R2977 VGND.n1760 VGND.n1759 27.5561
R2978 VGND.n241 VGND.n238 27.5561
R2979 VGND.n771 VGND.n770 27.2005
R2980 VGND.n866 VGND.n865 27.2005
R2981 VGND.n1156 VGND.n38 26.9584
R2982 VGND.n1700 VGND.n42 26.9584
R2983 VGND.n1930 VGND.n1929 26.6672
R2984 VGND.n1851 VGND.n1850 26.6672
R2985 VGND.n315 VGND.n298 26.6672
R2986 VGND.n398 VGND.n397 26.6672
R2987 VGND.n1512 VGND.n1511 26.6672
R2988 VGND.n1246 VGND.n1245 26.6672
R2989 VGND.n1418 VGND.n1417 26.6672
R2990 VGND.n1743 VGND.n1742 26.6672
R2991 VGND.n222 VGND.n221 26.6672
R2992 VGND.n758 VGND.n757 25.6005
R2993 VGND.n856 VGND.n855 25.6005
R2994 VGND.n2335 VGND.t193 25.5065
R2995 VGND.t193 VGND.n49 25.5065
R2996 VGND.t193 VGND.n40 25.5065
R2997 VGND.n651 VGND.n650 25.3679
R2998 VGND.n848 VGND.n847 24.8279
R2999 VGND.n861 VGND.n860 24.8279
R3000 VGND.n850 VGND.t161 24.0005
R3001 VGND.n850 VGND.t225 24.0005
R3002 VGND.n755 VGND.t259 24.0005
R3003 VGND.n755 VGND.t165 24.0005
R3004 VGND.n753 VGND.t70 24.0005
R3005 VGND.n753 VGND.t84 24.0005
R3006 VGND.n751 VGND.t18 24.0005
R3007 VGND.n751 VGND.t82 24.0005
R3008 VGND.t210 VGND.n859 24.0005
R3009 VGND.n859 VGND.t8 24.0005
R3010 VGND.n885 VGND.n874 22.4005
R3011 VGND.t39 VGND.n759 19.9551
R3012 VGND.n2357 VGND.n2356 18.8382
R3013 VGND.n1613 VGND.n1162 17.5843
R3014 VGND.n2272 VGND.n1686 17.5843
R3015 VGND.n495 VGND.n494 17.5843
R3016 VGND.n968 VGND.n459 16.9605
R3017 VGND.n2074 VGND.n1969 16.9379
R3018 VGND.n1041 VGND.n1040 16.9379
R3019 VGND.n1328 VGND.n1327 16.9379
R3020 VGND.n1161 VGND.n1160 16.7709
R3021 VGND.n2302 VGND.n2301 16.7709
R3022 VGND.n1977 VGND.n103 16.7709
R3023 VGND.n2330 VGND.n76 16.7709
R3024 VGND.n1947 VGND.n1905 16.0005
R3025 VGND.n1953 VGND.n1905 16.0005
R3026 VGND.n1954 VGND.n1953 16.0005
R3027 VGND.n1955 VGND.n1954 16.0005
R3028 VGND.n1955 VGND.n1903 16.0005
R3029 VGND.n1961 VGND.n1903 16.0005
R3030 VGND.n1962 VGND.n1961 16.0005
R3031 VGND.n2102 VGND.n1962 16.0005
R3032 VGND.n1946 VGND.n1945 16.0005
R3033 VGND.n1945 VGND.n1907 16.0005
R3034 VGND.n1939 VGND.n1907 16.0005
R3035 VGND.n1939 VGND.n1938 16.0005
R3036 VGND.n1938 VGND.n1937 16.0005
R3037 VGND.n1937 VGND.n1909 16.0005
R3038 VGND.n1931 VGND.n1909 16.0005
R3039 VGND.n1931 VGND.n1930 16.0005
R3040 VGND.n1929 VGND.n1911 16.0005
R3041 VGND.n1923 VGND.n1911 16.0005
R3042 VGND.n1923 VGND.n1922 16.0005
R3043 VGND.n1922 VGND.n1921 16.0005
R3044 VGND.n1921 VGND.n1913 16.0005
R3045 VGND.n1916 VGND.n1913 16.0005
R3046 VGND.n1916 VGND.n1890 16.0005
R3047 VGND.n2137 VGND.n1890 16.0005
R3048 VGND.n1868 VGND.n1826 16.0005
R3049 VGND.n1874 VGND.n1826 16.0005
R3050 VGND.n1875 VGND.n1874 16.0005
R3051 VGND.n1876 VGND.n1875 16.0005
R3052 VGND.n1876 VGND.n1824 16.0005
R3053 VGND.n1882 VGND.n1824 16.0005
R3054 VGND.n1883 VGND.n1882 16.0005
R3055 VGND.n2151 VGND.n1883 16.0005
R3056 VGND.n1867 VGND.n1866 16.0005
R3057 VGND.n1866 VGND.n1828 16.0005
R3058 VGND.n1860 VGND.n1828 16.0005
R3059 VGND.n1860 VGND.n1859 16.0005
R3060 VGND.n1859 VGND.n1858 16.0005
R3061 VGND.n1858 VGND.n1830 16.0005
R3062 VGND.n1852 VGND.n1830 16.0005
R3063 VGND.n1852 VGND.n1851 16.0005
R3064 VGND.n1850 VGND.n1832 16.0005
R3065 VGND.n1844 VGND.n1832 16.0005
R3066 VGND.n1844 VGND.n1843 16.0005
R3067 VGND.n1843 VGND.n1842 16.0005
R3068 VGND.n1842 VGND.n1834 16.0005
R3069 VGND.n1837 VGND.n1834 16.0005
R3070 VGND.n1837 VGND.n1811 16.0005
R3071 VGND.n2186 VGND.n1811 16.0005
R3072 VGND.n338 VGND.n337 16.0005
R3073 VGND.n339 VGND.n338 16.0005
R3074 VGND.n339 VGND.n292 16.0005
R3075 VGND.n345 VGND.n292 16.0005
R3076 VGND.n346 VGND.n345 16.0005
R3077 VGND.n347 VGND.n346 16.0005
R3078 VGND.n347 VGND.n290 16.0005
R3079 VGND.n352 VGND.n290 16.0005
R3080 VGND.n331 VGND.n294 16.0005
R3081 VGND.n331 VGND.n330 16.0005
R3082 VGND.n330 VGND.n329 16.0005
R3083 VGND.n329 VGND.n296 16.0005
R3084 VGND.n323 VGND.n296 16.0005
R3085 VGND.n323 VGND.n322 16.0005
R3086 VGND.n322 VGND.n321 16.0005
R3087 VGND.n321 VGND.n298 16.0005
R3088 VGND.n315 VGND.n314 16.0005
R3089 VGND.n314 VGND.n313 16.0005
R3090 VGND.n313 VGND.n300 16.0005
R3091 VGND.n308 VGND.n300 16.0005
R3092 VGND.n308 VGND.n307 16.0005
R3093 VGND.n307 VGND.n306 16.0005
R3094 VGND.n306 VGND.n280 16.0005
R3095 VGND.n1150 VGND.n280 16.0005
R3096 VGND.n418 VGND.n417 16.0005
R3097 VGND.n421 VGND.n418 16.0005
R3098 VGND.n422 VGND.n421 16.0005
R3099 VGND.n425 VGND.n422 16.0005
R3100 VGND.n426 VGND.n425 16.0005
R3101 VGND.n429 VGND.n426 16.0005
R3102 VGND.n431 VGND.n429 16.0005
R3103 VGND.n432 VGND.n431 16.0005
R3104 VGND.n414 VGND.n413 16.0005
R3105 VGND.n413 VGND.n410 16.0005
R3106 VGND.n410 VGND.n409 16.0005
R3107 VGND.n409 VGND.n406 16.0005
R3108 VGND.n406 VGND.n405 16.0005
R3109 VGND.n405 VGND.n402 16.0005
R3110 VGND.n402 VGND.n401 16.0005
R3111 VGND.n401 VGND.n398 16.0005
R3112 VGND.n397 VGND.n394 16.0005
R3113 VGND.n394 VGND.n393 16.0005
R3114 VGND.n393 VGND.n390 16.0005
R3115 VGND.n390 VGND.n389 16.0005
R3116 VGND.n389 VGND.n386 16.0005
R3117 VGND.n386 VGND.n385 16.0005
R3118 VGND.n385 VGND.n382 16.0005
R3119 VGND.n382 VGND.n358 16.0005
R3120 VGND.n1529 VGND.n1487 16.0005
R3121 VGND.n1535 VGND.n1487 16.0005
R3122 VGND.n1536 VGND.n1535 16.0005
R3123 VGND.n1537 VGND.n1536 16.0005
R3124 VGND.n1537 VGND.n1485 16.0005
R3125 VGND.n1543 VGND.n1485 16.0005
R3126 VGND.n1544 VGND.n1543 16.0005
R3127 VGND.n1547 VGND.n1544 16.0005
R3128 VGND.n1528 VGND.n1527 16.0005
R3129 VGND.n1527 VGND.n1489 16.0005
R3130 VGND.n1521 VGND.n1489 16.0005
R3131 VGND.n1521 VGND.n1520 16.0005
R3132 VGND.n1520 VGND.n1519 16.0005
R3133 VGND.n1519 VGND.n1491 16.0005
R3134 VGND.n1513 VGND.n1491 16.0005
R3135 VGND.n1513 VGND.n1512 16.0005
R3136 VGND.n1511 VGND.n1493 16.0005
R3137 VGND.n1505 VGND.n1493 16.0005
R3138 VGND.n1505 VGND.n1504 16.0005
R3139 VGND.n1504 VGND.n1503 16.0005
R3140 VGND.n1503 VGND.n1495 16.0005
R3141 VGND.n1498 VGND.n1495 16.0005
R3142 VGND.n1498 VGND.n1471 16.0005
R3143 VGND.n1582 VGND.n1471 16.0005
R3144 VGND.n1278 VGND.n1264 16.0005
R3145 VGND.n1278 VGND.n1277 16.0005
R3146 VGND.n1277 VGND.n1276 16.0005
R3147 VGND.n1276 VGND.n1273 16.0005
R3148 VGND.n1273 VGND.n1272 16.0005
R3149 VGND.n1272 VGND.n1269 16.0005
R3150 VGND.n1269 VGND.n1268 16.0005
R3151 VGND.n1268 VGND.n1265 16.0005
R3152 VGND.n1263 VGND.n1261 16.0005
R3153 VGND.n1261 VGND.n1258 16.0005
R3154 VGND.n1258 VGND.n1257 16.0005
R3155 VGND.n1257 VGND.n1254 16.0005
R3156 VGND.n1254 VGND.n1253 16.0005
R3157 VGND.n1253 VGND.n1250 16.0005
R3158 VGND.n1250 VGND.n1249 16.0005
R3159 VGND.n1249 VGND.n1246 16.0005
R3160 VGND.n1245 VGND.n1242 16.0005
R3161 VGND.n1242 VGND.n1241 16.0005
R3162 VGND.n1241 VGND.n1238 16.0005
R3163 VGND.n1238 VGND.n1237 16.0005
R3164 VGND.n1237 VGND.n1234 16.0005
R3165 VGND.n1234 VGND.n1233 16.0005
R3166 VGND.n1233 VGND.n1230 16.0005
R3167 VGND.n1230 VGND.n1229 16.0005
R3168 VGND.n1449 VGND.n1436 16.0005
R3169 VGND.n1449 VGND.n1448 16.0005
R3170 VGND.n1448 VGND.n1447 16.0005
R3171 VGND.n1447 VGND.n1444 16.0005
R3172 VGND.n1444 VGND.n1443 16.0005
R3173 VGND.n1443 VGND.n1440 16.0005
R3174 VGND.n1440 VGND.n1439 16.0005
R3175 VGND.n1439 VGND.n1352 16.0005
R3176 VGND.n1435 VGND.n1433 16.0005
R3177 VGND.n1433 VGND.n1430 16.0005
R3178 VGND.n1430 VGND.n1429 16.0005
R3179 VGND.n1429 VGND.n1426 16.0005
R3180 VGND.n1426 VGND.n1425 16.0005
R3181 VGND.n1425 VGND.n1422 16.0005
R3182 VGND.n1422 VGND.n1421 16.0005
R3183 VGND.n1421 VGND.n1418 16.0005
R3184 VGND.n1417 VGND.n1414 16.0005
R3185 VGND.n1414 VGND.n1413 16.0005
R3186 VGND.n1413 VGND.n1410 16.0005
R3187 VGND.n1410 VGND.n1409 16.0005
R3188 VGND.n1409 VGND.n1406 16.0005
R3189 VGND.n1406 VGND.n1405 16.0005
R3190 VGND.n1405 VGND.n1402 16.0005
R3191 VGND.n1402 VGND.n1401 16.0005
R3192 VGND.n1760 VGND.n1718 16.0005
R3193 VGND.n1766 VGND.n1718 16.0005
R3194 VGND.n1767 VGND.n1766 16.0005
R3195 VGND.n1768 VGND.n1767 16.0005
R3196 VGND.n1768 VGND.n1716 16.0005
R3197 VGND.n1774 VGND.n1716 16.0005
R3198 VGND.n1775 VGND.n1774 16.0005
R3199 VGND.n2206 VGND.n1775 16.0005
R3200 VGND.n1759 VGND.n1758 16.0005
R3201 VGND.n1758 VGND.n1720 16.0005
R3202 VGND.n1752 VGND.n1720 16.0005
R3203 VGND.n1752 VGND.n1751 16.0005
R3204 VGND.n1751 VGND.n1750 16.0005
R3205 VGND.n1750 VGND.n1722 16.0005
R3206 VGND.n1744 VGND.n1722 16.0005
R3207 VGND.n1744 VGND.n1743 16.0005
R3208 VGND.n1742 VGND.n1724 16.0005
R3209 VGND.n1736 VGND.n1724 16.0005
R3210 VGND.n1736 VGND.n1735 16.0005
R3211 VGND.n1735 VGND.n1734 16.0005
R3212 VGND.n1734 VGND.n1726 16.0005
R3213 VGND.n1729 VGND.n1726 16.0005
R3214 VGND.n1729 VGND.n1703 16.0005
R3215 VGND.n2241 VGND.n1703 16.0005
R3216 VGND.n242 VGND.n241 16.0005
R3217 VGND.n245 VGND.n242 16.0005
R3218 VGND.n246 VGND.n245 16.0005
R3219 VGND.n249 VGND.n246 16.0005
R3220 VGND.n250 VGND.n249 16.0005
R3221 VGND.n253 VGND.n250 16.0005
R3222 VGND.n254 VGND.n253 16.0005
R3223 VGND.n257 VGND.n254 16.0005
R3224 VGND.n238 VGND.n237 16.0005
R3225 VGND.n237 VGND.n234 16.0005
R3226 VGND.n234 VGND.n233 16.0005
R3227 VGND.n233 VGND.n230 16.0005
R3228 VGND.n230 VGND.n229 16.0005
R3229 VGND.n229 VGND.n226 16.0005
R3230 VGND.n226 VGND.n225 16.0005
R3231 VGND.n225 VGND.n222 16.0005
R3232 VGND.n221 VGND.n218 16.0005
R3233 VGND.n218 VGND.n217 16.0005
R3234 VGND.n217 VGND.n214 16.0005
R3235 VGND.n214 VGND.n213 16.0005
R3236 VGND.n213 VGND.n210 16.0005
R3237 VGND.n210 VGND.n209 16.0005
R3238 VGND.n209 VGND.n206 16.0005
R3239 VGND.n206 VGND.n205 16.0005
R3240 VGND.n1037 VGND.n443 15.1758
R3241 VGND.n1037 VGND.n1036 15.1758
R3242 VGND.n1036 VGND.n1035 15.1758
R3243 VGND.n1035 VGND.n444 15.1758
R3244 VGND.n1029 VGND.n444 15.1758
R3245 VGND.n1028 VGND.n1027 15.1758
R3246 VGND.n1027 VGND.n448 15.1758
R3247 VGND.n1021 VGND.n448 15.1758
R3248 VGND.n1021 VGND.n1020 15.1758
R3249 VGND.n1020 VGND.n36 15.1758
R3250 VGND.n978 VGND.n35 15.1758
R3251 VGND.n978 VGND.n977 15.1758
R3252 VGND.n977 VGND.n976 15.1758
R3253 VGND.n976 VGND.n456 15.1758
R3254 VGND.n970 VGND.n456 15.1758
R3255 VGND.n575 VGND.n574 15.1758
R3256 VGND.n574 VGND.n462 15.1758
R3257 VGND.n568 VGND.n462 15.1758
R3258 VGND.n568 VGND.n567 15.1758
R3259 VGND.n567 VGND.n566 15.1758
R3260 VGND.n516 VGND.n515 15.1758
R3261 VGND.n515 VGND.n514 15.1758
R3262 VGND.n514 VGND.n472 15.1758
R3263 VGND.n508 VGND.n472 15.1758
R3264 VGND.n508 VGND.n507 15.1758
R3265 VGND.n506 VGND.n477 15.1758
R3266 VGND.n500 VGND.n477 15.1758
R3267 VGND.n500 VGND.n499 15.1758
R3268 VGND.n499 VGND.n498 15.1758
R3269 VGND.n498 VGND.n481 15.1758
R3270 VGND.n839 VGND.t207 15.0005
R3271 VGND.n827 VGND.t40 15.0005
R3272 VGND.n827 VGND.t206 15.0005
R3273 VGND.n825 VGND.t217 15.0005
R3274 VGND.n825 VGND.t4 15.0005
R3275 VGND.n804 VGND.t265 15.0005
R3276 VGND.n804 VGND.t202 15.0005
R3277 VGND.n802 VGND.t198 15.0005
R3278 VGND.n802 VGND.t253 15.0005
R3279 VGND.n784 VGND.t286 15.0005
R3280 VGND.n784 VGND.t221 15.0005
R3281 VGND.n782 VGND.t234 15.0005
R3282 VGND.n782 VGND.t16 15.0005
R3283 VGND.t234 VGND.n781 15.0005
R3284 VGND.t217 VGND.n824 15.0005
R3285 VGND.n816 VGND.t203 15.0005
R3286 VGND.t198 VGND.n801 15.0005
R3287 VGND.n792 VGND.t222 15.0005
R3288 VGND.t175 VGND.t17 14.9665
R3289 VGND.t252 VGND.t155 14.9665
R3290 VGND.n819 VGND.t111 14.9665
R3291 VGND.t212 VGND.t224 14.9665
R3292 VGND.n1468 VGND.n47 14.555
R3293 VGND.n770 VGND.n743 14.0805
R3294 VGND.n865 VGND.n864 14.0805
R3295 VGND.n849 VGND.n848 14.0349
R3296 VGND.n862 VGND.n861 14.0349
R3297 VGND.n617 VGND.n616 12.8005
R3298 VGND.n616 VGND.n613 12.8005
R3299 VGND.n757 VGND.n750 12.8005
R3300 VGND.n855 VGND.n854 12.8005
R3301 VGND.n621 VGND.n605 12.8005
R3302 VGND.n606 VGND.n605 12.8005
R3303 VGND.n963 VGND.n577 12.8005
R3304 VGND.n968 VGND.n577 12.8005
R3305 VGND.t193 VGND.n24 12.1263
R3306 VGND.t193 VGND.n48 12.1263
R3307 VGND.t193 VGND.n41 12.1263
R3308 VGND.n2356 VGND.t300 12.051
R3309 VGND.n662 VGND.t58 12.0198
R3310 VGND.n609 VGND.t0 11.7213
R3311 VGND.n2075 VGND.n2074 11.6369
R3312 VGND.n2076 VGND.n2075 11.6369
R3313 VGND.n2076 VGND.n1967 11.6369
R3314 VGND.n2082 VGND.n1967 11.6369
R3315 VGND.n2083 VGND.n2082 11.6369
R3316 VGND.n2084 VGND.n2083 11.6369
R3317 VGND.n2084 VGND.n1965 11.6369
R3318 VGND.n2090 VGND.n1965 11.6369
R3319 VGND.n2091 VGND.n2090 11.6369
R3320 VGND.n2092 VGND.n2091 11.6369
R3321 VGND.n1040 VGND.n1039 11.6369
R3322 VGND.n1039 VGND.n441 11.6369
R3323 VGND.n1033 VGND.n441 11.6369
R3324 VGND.n1033 VGND.n1032 11.6369
R3325 VGND.n1032 VGND.n1031 11.6369
R3326 VGND.n1031 VGND.n446 11.6369
R3327 VGND.n1025 VGND.n446 11.6369
R3328 VGND.n1025 VGND.n1024 11.6369
R3329 VGND.n1024 VGND.n1023 11.6369
R3330 VGND.n1023 VGND.n450 11.6369
R3331 VGND.n1017 VGND.n450 11.6369
R3332 VGND.n1041 VGND.n439 11.6369
R3333 VGND.n439 VGND.n438 11.6369
R3334 VGND.n1048 VGND.n438 11.6369
R3335 VGND.n1049 VGND.n1048 11.6369
R3336 VGND.n1050 VGND.n1049 11.6369
R3337 VGND.n1050 VGND.n436 11.6369
R3338 VGND.n1056 VGND.n436 11.6369
R3339 VGND.n1057 VGND.n1056 11.6369
R3340 VGND.n1058 VGND.n1057 11.6369
R3341 VGND.n1058 VGND.n434 11.6369
R3342 VGND.n123 VGND.n75 11.6369
R3343 VGND.n126 VGND.n123 11.6369
R3344 VGND.n127 VGND.n126 11.6369
R3345 VGND.n130 VGND.n127 11.6369
R3346 VGND.n131 VGND.n130 11.6369
R3347 VGND.n134 VGND.n131 11.6369
R3348 VGND.n135 VGND.n134 11.6369
R3349 VGND.n138 VGND.n135 11.6369
R3350 VGND.n139 VGND.n138 11.6369
R3351 VGND.n142 VGND.n139 11.6369
R3352 VGND.n143 VGND.n142 11.6369
R3353 VGND.n1634 VGND.n1633 11.6369
R3354 VGND.n1633 VGND.n1630 11.6369
R3355 VGND.n1630 VGND.n1629 11.6369
R3356 VGND.n1629 VGND.n1626 11.6369
R3357 VGND.n1626 VGND.n1625 11.6369
R3358 VGND.n1625 VGND.n1622 11.6369
R3359 VGND.n1622 VGND.n1621 11.6369
R3360 VGND.n1621 VGND.n1618 11.6369
R3361 VGND.n1618 VGND.n1617 11.6369
R3362 VGND.n1617 VGND.n1614 11.6369
R3363 VGND.n1614 VGND.n1613 11.6369
R3364 VGND.n1166 VGND.n1162 11.6369
R3365 VGND.n1606 VGND.n1166 11.6369
R3366 VGND.n1606 VGND.n1605 11.6369
R3367 VGND.n1605 VGND.n1604 11.6369
R3368 VGND.n1604 VGND.n1167 11.6369
R3369 VGND.n1599 VGND.n1167 11.6369
R3370 VGND.n1599 VGND.n1598 11.6369
R3371 VGND.n1598 VGND.n1597 11.6369
R3372 VGND.n1597 VGND.n1169 11.6369
R3373 VGND.n1591 VGND.n1169 11.6369
R3374 VGND.n1327 VGND.n1326 11.6369
R3375 VGND.n1326 VGND.n1323 11.6369
R3376 VGND.n1323 VGND.n1322 11.6369
R3377 VGND.n1322 VGND.n1319 11.6369
R3378 VGND.n1319 VGND.n1318 11.6369
R3379 VGND.n1318 VGND.n1315 11.6369
R3380 VGND.n1315 VGND.n1314 11.6369
R3381 VGND.n1314 VGND.n1311 11.6369
R3382 VGND.n1311 VGND.n1310 11.6369
R3383 VGND.n1310 VGND.n74 11.6369
R3384 VGND.n2331 VGND.n74 11.6369
R3385 VGND.n1328 VGND.n1307 11.6369
R3386 VGND.n1334 VGND.n1307 11.6369
R3387 VGND.n1335 VGND.n1334 11.6369
R3388 VGND.n1336 VGND.n1335 11.6369
R3389 VGND.n1336 VGND.n1305 11.6369
R3390 VGND.n1342 VGND.n1305 11.6369
R3391 VGND.n1343 VGND.n1342 11.6369
R3392 VGND.n1344 VGND.n1343 11.6369
R3393 VGND.n1344 VGND.n1303 11.6369
R3394 VGND.n1303 VGND.n1302 11.6369
R3395 VGND.n1689 VGND.n1686 11.6369
R3396 VGND.n1692 VGND.n1689 11.6369
R3397 VGND.n2264 VGND.n1692 11.6369
R3398 VGND.n2264 VGND.n2263 11.6369
R3399 VGND.n2263 VGND.n2262 11.6369
R3400 VGND.n2262 VGND.n1693 11.6369
R3401 VGND.n1695 VGND.n1693 11.6369
R3402 VGND.n1698 VGND.n1695 11.6369
R3403 VGND.n2254 VGND.n1698 11.6369
R3404 VGND.n2254 VGND.n2253 11.6369
R3405 VGND.n2288 VGND.n1672 11.6369
R3406 VGND.n2288 VGND.n2287 11.6369
R3407 VGND.n2287 VGND.n2286 11.6369
R3408 VGND.n2286 VGND.n1680 11.6369
R3409 VGND.n2281 VGND.n1680 11.6369
R3410 VGND.n2281 VGND.n2280 11.6369
R3411 VGND.n2280 VGND.n2279 11.6369
R3412 VGND.n2279 VGND.n1683 11.6369
R3413 VGND.n2274 VGND.n1683 11.6369
R3414 VGND.n2274 VGND.n2273 11.6369
R3415 VGND.n2273 VGND.n2272 11.6369
R3416 VGND.n494 VGND.n483 11.6369
R3417 VGND.n488 VGND.n483 11.6369
R3418 VGND.n488 VGND.n487 11.6369
R3419 VGND.n487 VGND.n26 11.6369
R3420 VGND.n2337 VGND.n26 11.6369
R3421 VGND.n2338 VGND.n2337 11.6369
R3422 VGND.n2339 VGND.n2338 11.6369
R3423 VGND.n2339 VGND.n22 11.6369
R3424 VGND.n2345 VGND.n22 11.6369
R3425 VGND.n2346 VGND.n2345 11.6369
R3426 VGND.n474 VGND.n469 11.6369
R3427 VGND.n512 VGND.n474 11.6369
R3428 VGND.n512 VGND.n511 11.6369
R3429 VGND.n511 VGND.n510 11.6369
R3430 VGND.n510 VGND.n475 11.6369
R3431 VGND.n504 VGND.n475 11.6369
R3432 VGND.n504 VGND.n503 11.6369
R3433 VGND.n503 VGND.n502 11.6369
R3434 VGND.n502 VGND.n479 11.6369
R3435 VGND.n496 VGND.n479 11.6369
R3436 VGND.n496 VGND.n495 11.6369
R3437 VGND.n455 VGND.n452 11.6369
R3438 VGND.n458 VGND.n455 11.6369
R3439 VGND.n974 VGND.n458 11.6369
R3440 VGND.n974 VGND.n973 11.6369
R3441 VGND.n973 VGND.n972 11.6369
R3442 VGND.n572 VGND.n464 11.6369
R3443 VGND.n572 VGND.n571 11.6369
R3444 VGND.n571 VGND.n570 11.6369
R3445 VGND.n570 VGND.n465 11.6369
R3446 VGND.n564 VGND.n465 11.6369
R3447 VGND.n2040 VGND.n2018 11.6369
R3448 VGND.n2040 VGND.n2039 11.6369
R3449 VGND.n2039 VGND.n2038 11.6369
R3450 VGND.n2038 VGND.n2020 11.6369
R3451 VGND.n2033 VGND.n2020 11.6369
R3452 VGND.n2033 VGND.n2032 11.6369
R3453 VGND.n2032 VGND.n2031 11.6369
R3454 VGND.n2031 VGND.n2023 11.6369
R3455 VGND.n2026 VGND.n2023 11.6369
R3456 VGND.n2026 VGND.n1674 11.6369
R3457 VGND.n2300 VGND.n1674 11.6369
R3458 VGND.n2068 VGND.n1969 11.6369
R3459 VGND.n2068 VGND.n2067 11.6369
R3460 VGND.n2067 VGND.n2066 11.6369
R3461 VGND.n2066 VGND.n1971 11.6369
R3462 VGND.n2061 VGND.n1971 11.6369
R3463 VGND.n2061 VGND.n2060 11.6369
R3464 VGND.n2060 VGND.n2059 11.6369
R3465 VGND.n2059 VGND.n1974 11.6369
R3466 VGND.n2054 VGND.n1974 11.6369
R3467 VGND.n2054 VGND.n2053 11.6369
R3468 VGND.n2053 VGND.n2052 11.6369
R3469 VGND.n2356 VGND.t303 11.4829
R3470 VGND.t17 VGND.t197 9.97782
R3471 VGND.n635 VGND.t62 9.6005
R3472 VGND.n657 VGND.t61 9.6005
R3473 VGND.n643 VGND.t59 9.6005
R3474 VGND.n649 VGND.t60 9.6005
R3475 VGND.n617 VGND.n611 9.36264
R3476 VGND.n606 VGND.n603 9.36264
R3477 VGND.n964 VGND.n963 9.36264
R3478 VGND.n956 VGND.n955 9.32966
R3479 VGND.n616 VGND.n615 9.3005
R3480 VGND.n614 VGND.n613 9.3005
R3481 VGND.n835 VGND.n832 9.3005
R3482 VGND.n840 VGND.n831 9.3005
R3483 VGND.n778 VGND.n766 9.3005
R3484 VGND.n780 VGND.n779 9.3005
R3485 VGND.n605 VGND.n604 9.3005
R3486 VGND.n622 VGND.n621 9.3005
R3487 VGND.n578 VGND.n577 9.3005
R3488 VGND.n968 VGND.n967 9.3005
R3489 VGND.n886 VGND.n885 9.3005
R3490 VGND.n890 VGND.n889 9.3005
R3491 VGND.n894 VGND.n893 9.3005
R3492 VGND.n884 VGND.n877 9.3005
R3493 VGND.n54 VGND.t143 8.78127
R3494 VGND.n2304 VGND.n47 8.60107
R3495 VGND.n1029 VGND.t193 7.92539
R3496 VGND.n970 VGND.t193 7.92539
R3497 VGND.n507 VGND.t193 7.92539
R3498 VGND.t193 VGND.n1028 7.25093
R3499 VGND.t193 VGND.n575 7.25093
R3500 VGND.t193 VGND.n506 7.25093
R3501 VGND.n840 VGND.n832 7.11161
R3502 VGND.n780 VGND.n766 7.11161
R3503 VGND.n2382 VGND.n0 7.09427
R3504 VGND.n1017 VGND.n1016 6.72373
R3505 VGND.n1161 VGND.n143 6.72373
R3506 VGND.n2331 VGND.n2330 6.72373
R3507 VGND.n564 VGND.n563 6.72373
R3508 VGND.n2301 VGND.n2300 6.72373
R3509 VGND.n2052 VGND.n1977 6.72373
R3510 VGND.t27 VGND.n54 6.69061
R3511 VGND.n2330 VGND.n75 6.20656
R3512 VGND.n1634 VGND.n1161 6.20656
R3513 VGND.n2301 VGND.n1672 6.20656
R3514 VGND.n563 VGND.n469 6.20656
R3515 VGND.n1016 VGND.n452 6.20656
R3516 VGND.n2018 VGND.n1977 6.20656
R3517 VGND.n972 VGND.n459 6.07727
R3518 VGND.n887 VGND.n877 5.84425
R3519 VGND.n651 VGND.n641 5.81868
R3520 VGND.n651 VGND.n642 5.81868
R3521 VGND.n716 VGND.n715 5.68939
R3522 VGND.n715 VGND.n714 5.68939
R3523 VGND.n706 VGND.n673 5.68939
R3524 VGND.n464 VGND.n459 5.5601
R3525 VGND.n2138 VGND.n2137 5.51161
R3526 VGND.n2187 VGND.n2186 5.51161
R3527 VGND.n1152 VGND.n1150 5.51161
R3528 VGND.n1103 VGND.n358 5.51161
R3529 VGND.n1583 VGND.n1582 5.51161
R3530 VGND.n1229 VGND.n1207 5.51161
R3531 VGND.n1401 VGND.n1379 5.51161
R3532 VGND.n2242 VGND.n2241 5.51161
R3533 VGND.n205 VGND.n176 5.51161
R3534 VGND.t58 VGND.n43 5.25917
R3535 VGND.n1590 VGND.n1174 5.1717
R3536 VGND.n2252 VGND.n1699 5.1717
R3537 VGND.n2347 VGND.n21 5.1717
R3538 VGND.n893 VGND.n0 5.07862
R3539 VGND.n889 VGND.n888 5.07862
R3540 VGND.n887 VGND.n886 5.07862
R3541 VGND.t95 VGND.n18 5.01808
R3542 VGND.n773 VGND.t9 4.98916
R3543 VGND.t220 VGND.t91 4.98916
R3544 VGND.t91 VGND.t209 4.98916
R3545 VGND.t135 VGND.t164 4.98916
R3546 VGND.n783 VGND.n763 4.98488
R3547 VGND.n706 VGND.n705 4.97828
R3548 VGND.n2099 VGND.n1963 4.9157
R3549 VGND.n1066 VGND.n433 4.9157
R3550 VGND.n1465 VGND.n1351 4.9157
R3551 VGND.n815 VGND.n806 4.78398
R3552 VGND.n794 VGND.n786 4.78398
R3553 VGND.n830 VGND.n829 4.64112
R3554 VGND.n2351 VGND.n17 4.59995
R3555 VGND.n597 VGND.n596 4.5005
R3556 VGND.n624 VGND.n599 4.5005
R3557 VGND.n626 VGND.n625 4.5005
R3558 VGND.n625 VGND.n624 4.5005
R3559 VGND.n614 VGND.n601 4.5005
R3560 VGND.n623 VGND.n622 4.5005
R3561 VGND.n967 VGND.n966 4.5005
R3562 VGND.n562 VGND.n470 4.26717
R3563 VGND.n557 VGND.n470 4.26717
R3564 VGND.n557 VGND.n556 4.26717
R3565 VGND.n556 VGND.n524 4.26717
R3566 VGND.n551 VGND.n524 4.26717
R3567 VGND.n551 VGND.n550 4.26717
R3568 VGND.n550 VGND.n549 4.26717
R3569 VGND.n549 VGND.n532 4.26717
R3570 VGND.n543 VGND.n532 4.26717
R3571 VGND.n543 VGND.n542 4.26717
R3572 VGND.n542 VGND.n541 4.26717
R3573 VGND.n1638 VGND.n121 4.26717
R3574 VGND.n1644 VGND.n121 4.26717
R3575 VGND.n1644 VGND.n119 4.26717
R3576 VGND.n1650 VGND.n119 4.26717
R3577 VGND.n1650 VGND.n117 4.26717
R3578 VGND.n1658 VGND.n117 4.26717
R3579 VGND.n1658 VGND.n115 4.26717
R3580 VGND.n115 VGND.n112 4.26717
R3581 VGND.n1665 VGND.n112 4.26717
R3582 VGND.n1665 VGND.n110 4.26717
R3583 VGND.n1670 VGND.n110 4.26717
R3584 VGND.n2295 VGND.n1673 4.26717
R3585 VGND.n2295 VGND.n1677 4.26717
R3586 VGND.n1787 VGND.n1677 4.26717
R3587 VGND.n1792 VGND.n1787 4.26717
R3588 VGND.n1792 VGND.n1784 4.26717
R3589 VGND.n1798 VGND.n1784 4.26717
R3590 VGND.n1798 VGND.n1782 4.26717
R3591 VGND.n1804 VGND.n1782 4.26717
R3592 VGND.n1804 VGND.n1780 4.26717
R3593 VGND.n2196 VGND.n1780 4.26717
R3594 VGND.n2196 VGND.n1778 4.26717
R3595 VGND.n2047 VGND.n1979 4.26717
R3596 VGND.n2047 VGND.n1981 4.26717
R3597 VGND.n2014 VGND.n1981 4.26717
R3598 VGND.n2014 VGND.n2013 4.26717
R3599 VGND.n2013 VGND.n2012 4.26717
R3600 VGND.n2012 VGND.n1988 4.26717
R3601 VGND.n2006 VGND.n1988 4.26717
R3602 VGND.n2006 VGND.n2005 4.26717
R3603 VGND.n2005 VGND.n2004 4.26717
R3604 VGND.n2004 VGND.n1999 4.26717
R3605 VGND.n1999 VGND.n1998 4.26717
R3606 VGND.n2329 VGND.n77 4.26717
R3607 VGND.n2324 VGND.n77 4.26717
R3608 VGND.n2324 VGND.n2323 4.26717
R3609 VGND.n2323 VGND.n85 4.26717
R3610 VGND.n2318 VGND.n85 4.26717
R3611 VGND.n2318 VGND.n2317 4.26717
R3612 VGND.n2317 VGND.n2316 4.26717
R3613 VGND.n2316 VGND.n93 4.26717
R3614 VGND.n2310 VGND.n93 4.26717
R3615 VGND.n2310 VGND.n2309 4.26717
R3616 VGND.n2309 VGND.n2308 4.26717
R3617 VGND.n1015 VGND.n453 4.26717
R3618 VGND.n1010 VGND.n453 4.26717
R3619 VGND.n1010 VGND.n1009 4.26717
R3620 VGND.n1009 VGND.n987 4.26717
R3621 VGND.n1004 VGND.n987 4.26717
R3622 VGND.n1004 VGND.n1003 4.26717
R3623 VGND.n1003 VGND.n1002 4.26717
R3624 VGND.n1002 VGND.n997 4.26717
R3625 VGND.n997 VGND.n356 4.26717
R3626 VGND.n1110 VGND.n356 4.26717
R3627 VGND.n1110 VGND.n354 4.26717
R3628 VGND.n2376 VGND.n7 4.17862
R3629 VGND.n2372 VGND.n10 4.17862
R3630 VGND.n2380 VGND.n4 4.01225
R3631 VGND.n563 VGND.n562 3.93531
R3632 VGND.n1638 VGND.n1161 3.93531
R3633 VGND.n2301 VGND.n1673 3.93531
R3634 VGND.n1979 VGND.n1977 3.93531
R3635 VGND.n2330 VGND.n2329 3.93531
R3636 VGND.n1016 VGND.n1015 3.93531
R3637 VGND.n2100 VGND.n1901 3.7893
R3638 VGND.n2109 VGND.n2108 3.7893
R3639 VGND.n1899 VGND.n1898 3.7893
R3640 VGND.n2117 VGND.n2115 3.7893
R3641 VGND.n2116 VGND.n1896 3.7893
R3642 VGND.n2124 VGND.n2123 3.7893
R3643 VGND.n1894 VGND.n1893 3.7893
R3644 VGND.n2132 VGND.n2130 3.7893
R3645 VGND.n2131 VGND.n1889 3.7893
R3646 VGND.n2149 VGND.n1822 3.7893
R3647 VGND.n2158 VGND.n2157 3.7893
R3648 VGND.n1820 VGND.n1819 3.7893
R3649 VGND.n2166 VGND.n2164 3.7893
R3650 VGND.n2165 VGND.n1817 3.7893
R3651 VGND.n2173 VGND.n2172 3.7893
R3652 VGND.n1815 VGND.n1814 3.7893
R3653 VGND.n2181 VGND.n2179 3.7893
R3654 VGND.n2180 VGND.n1810 3.7893
R3655 VGND.n1121 VGND.n1120 3.7893
R3656 VGND.n1125 VGND.n288 3.7893
R3657 VGND.n1126 VGND.n287 3.7893
R3658 VGND.n1133 VGND.n1129 3.7893
R3659 VGND.n1132 VGND.n285 3.7893
R3660 VGND.n1139 VGND.n284 3.7893
R3661 VGND.n1140 VGND.n283 3.7893
R3662 VGND.n1145 VGND.n1143 3.7893
R3663 VGND.n1144 VGND.n279 3.7893
R3664 VGND.n1093 VGND.n1068 3.7893
R3665 VGND.n1092 VGND.n1089 3.7893
R3666 VGND.n1088 VGND.n1069 3.7893
R3667 VGND.n1085 VGND.n1084 3.7893
R3668 VGND.n1081 VGND.n1070 3.7893
R3669 VGND.n1078 VGND.n1077 3.7893
R3670 VGND.n1074 VGND.n1071 3.7893
R3671 VGND.n1098 VGND.n360 3.7893
R3672 VGND.n1099 VGND.n359 3.7893
R3673 VGND.n1545 VGND.n1483 3.7893
R3674 VGND.n1554 VGND.n1553 3.7893
R3675 VGND.n1480 VGND.n1479 3.7893
R3676 VGND.n1562 VGND.n1560 3.7893
R3677 VGND.n1561 VGND.n1477 3.7893
R3678 VGND.n1569 VGND.n1568 3.7893
R3679 VGND.n1475 VGND.n1474 3.7893
R3680 VGND.n1577 VGND.n1575 3.7893
R3681 VGND.n1576 VGND.n1470 3.7893
R3682 VGND.n1292 VGND.n1291 3.7893
R3683 VGND.n1288 VGND.n1184 3.7893
R3684 VGND.n1287 VGND.n1187 3.7893
R3685 VGND.n1284 VGND.n1283 3.7893
R3686 VGND.n1209 VGND.n1188 3.7893
R3687 VGND.n1214 VGND.n1212 3.7893
R3688 VGND.n1218 VGND.n1217 3.7893
R3689 VGND.n1221 VGND.n1208 3.7893
R3690 VGND.n1226 VGND.n1222 3.7893
R3691 VGND.n1463 VGND.n1462 3.7893
R3692 VGND.n1459 VGND.n1354 3.7893
R3693 VGND.n1458 VGND.n1357 3.7893
R3694 VGND.n1455 VGND.n1454 3.7893
R3695 VGND.n1381 VGND.n1358 3.7893
R3696 VGND.n1386 VGND.n1384 3.7893
R3697 VGND.n1390 VGND.n1389 3.7893
R3698 VGND.n1393 VGND.n1380 3.7893
R3699 VGND.n1398 VGND.n1394 3.7893
R3700 VGND.n2204 VGND.n1714 3.7893
R3701 VGND.n2213 VGND.n2212 3.7893
R3702 VGND.n1712 VGND.n1711 3.7893
R3703 VGND.n2221 VGND.n2219 3.7893
R3704 VGND.n2220 VGND.n1709 3.7893
R3705 VGND.n2228 VGND.n2227 3.7893
R3706 VGND.n1707 VGND.n1706 3.7893
R3707 VGND.n2236 VGND.n2234 3.7893
R3708 VGND.n2235 VGND.n1702 3.7893
R3709 VGND.n255 VGND.n155 3.7893
R3710 VGND.n263 VGND.n262 3.7893
R3711 VGND.n179 VGND.n156 3.7893
R3712 VGND.n183 VGND.n181 3.7893
R3713 VGND.n187 VGND.n186 3.7893
R3714 VGND.n190 VGND.n178 3.7893
R3715 VGND.n194 VGND.n193 3.7893
R3716 VGND.n197 VGND.n177 3.7893
R3717 VGND.n202 VGND.n198 3.7893
R3718 VGND.n849 VGND.n581 3.63619
R3719 VGND.n836 VGND.n835 3.55702
R3720 VGND.n778 VGND.n777 3.55702
R3721 VGND.n833 VGND.n832 3.48951
R3722 VGND.n834 VGND.n833 3.48951
R3723 VGND.n766 VGND.n764 3.48951
R3724 VGND.n776 VGND.n764 3.48951
R3725 VGND.n2380 VGND.n2378 3.4105
R3726 VGND.n2381 VGND.n2380 3.4105
R3727 VGND.n2376 VGND.n2374 3.4105
R3728 VGND.n2377 VGND.n2376 3.4105
R3729 VGND.n2372 VGND.n2370 3.4105
R3730 VGND.n2373 VGND.n2372 3.4105
R3731 VGND.n2368 VGND.n2366 3.4105
R3732 VGND.n2369 VGND.n2368 3.4105
R3733 VGND.n2364 VGND.n2362 3.4105
R3734 VGND.n2365 VGND.n2364 3.4105
R3735 VGND.n2359 VGND.n2357 3.4105
R3736 VGND.n2361 VGND.n2360 3.4105
R3737 VGND.n2359 VGND.n2358 3.4105
R3738 VGND.n2360 VGND.n2359 3.4105
R3739 VGND.n829 VGND.n13 3.16181
R3740 VGND.n810 VGND.n809 3.14514
R3741 VGND.n790 VGND.n789 3.14514
R3742 VGND.n822 VGND.n810 3.1005
R3743 VGND.n814 VGND.n813 3.1005
R3744 VGND.n817 VGND.n815 3.1005
R3745 VGND.n799 VGND.n790 3.1005
R3746 VGND.n796 VGND.n795 3.1005
R3747 VGND.n794 VGND.n793 3.1005
R3748 VGND.n2368 VGND.n13 3.08096
R3749 VGND.n637 VGND.n636 2.86505
R3750 VGND.n637 VGND.n594 2.86505
R3751 VGND.n659 VGND.n591 2.86505
R3752 VGND.n659 VGND.n658 2.86505
R3753 VGND.n594 VGND.n593 2.86505
R3754 VGND.n658 VGND.n592 2.86505
R3755 VGND.n656 VGND.n636 2.86505
R3756 VGND.n593 VGND.n591 2.86505
R3757 VGND.n645 VGND.n644 2.86505
R3758 VGND.n648 VGND.n645 2.86505
R3759 VGND.n648 VGND.n647 2.86505
R3760 VGND.n644 VGND.n642 2.86505
R3761 VGND.n2101 VGND.n2099 2.6629
R3762 VGND.n1887 VGND.n1884 2.6629
R3763 VGND.n2150 VGND.n2148 2.6629
R3764 VGND.n1808 VGND.n1776 2.6629
R3765 VGND.n1117 VGND.n1116 2.6629
R3766 VGND.n1151 VGND.n144 2.6629
R3767 VGND.n1067 VGND.n1066 2.6629
R3768 VGND.n1104 VGND.n353 2.6629
R3769 VGND.n1546 VGND.n108 2.6629
R3770 VGND.n1183 VGND.n1182 2.6629
R3771 VGND.n1671 VGND.n109 2.6629
R3772 VGND.n1465 VGND.n1464 2.6629
R3773 VGND.n1378 VGND.n101 2.6629
R3774 VGND.n2205 VGND.n2203 2.6629
R3775 VGND.n256 VGND.n147 2.6629
R3776 VGND.n838 VGND.n836 2.60059
R3777 VGND.n777 VGND.n765 2.60059
R3778 VGND.n2364 VGND.n2352 2.59541
R3779 VGND.n836 VGND.n834 2.55763
R3780 VGND.n777 VGND.n776 2.55763
R3781 VGND.n2138 VGND.n1887 2.4581
R3782 VGND.n2148 VGND.n1884 2.4581
R3783 VGND.n2187 VGND.n1808 2.4581
R3784 VGND.n1116 VGND.n353 2.4581
R3785 VGND.n1152 VGND.n1151 2.4581
R3786 VGND.n1104 VGND.n1103 2.4581
R3787 VGND.n1671 VGND.n108 2.4581
R3788 VGND.n1583 VGND.n1174 2.4581
R3789 VGND.n1182 VGND.n101 2.4581
R3790 VGND.n1207 VGND.n109 2.4581
R3791 VGND.n1379 VGND.n1378 2.4581
R3792 VGND.n2203 VGND.n1776 2.4581
R3793 VGND.n2242 VGND.n1699 2.4581
R3794 VGND.n147 VGND.n144 2.4581
R3795 VGND.n176 VGND.n21 2.4581
R3796 VGND.n957 VGND.n956 2.44675
R3797 VGND.n956 VGND.n579 2.44675
R3798 VGND.n955 VGND.n580 2.36678
R3799 VGND.n633 VGND.n632 2.26187
R3800 VGND.n813 VGND.n807 2.25882
R3801 VGND.n813 VGND.n811 2.25882
R3802 VGND.n823 VGND.n809 2.25882
R3803 VGND.n822 VGND.n811 2.25882
R3804 VGND.n817 VGND.n807 2.25882
R3805 VGND.n823 VGND.n822 2.25882
R3806 VGND.n796 VGND.n787 2.25882
R3807 VGND.n796 VGND.n791 2.25882
R3808 VGND.n800 VGND.n789 2.25882
R3809 VGND.n799 VGND.n791 2.25882
R3810 VGND.n793 VGND.n787 2.25882
R3811 VGND.n800 VGND.n799 2.25882
R3812 VGND.n631 VGND.n630 2.24063
R3813 VGND.n629 VGND.n595 2.24063
R3814 VGND.n627 VGND.n626 2.24063
R3815 VGND.n602 VGND.n600 2.24063
R3816 VGND.n634 VGND.n633 2.24063
R3817 VGND.n628 VGND.n598 2.24063
R3818 VGND.n611 VGND.n601 2.22018
R3819 VGND.n623 VGND.n603 2.22018
R3820 VGND.n966 VGND.n964 2.22018
R3821 VGND.n541 VGND.n144 2.18124
R3822 VGND.n1671 VGND.n1670 2.18124
R3823 VGND.n1778 VGND.n1776 2.18124
R3824 VGND.n1998 VGND.n1884 2.18124
R3825 VGND.n2308 VGND.n101 2.18124
R3826 VGND.n354 VGND.n353 2.18124
R3827 VGND.n2139 VGND.n2138 2.1509
R3828 VGND.n2188 VGND.n2187 2.1509
R3829 VGND.n1153 VGND.n1152 2.1509
R3830 VGND.n1103 VGND.n1102 2.1509
R3831 VGND.n1584 VGND.n1583 2.1509
R3832 VGND.n1225 VGND.n1207 2.1509
R3833 VGND.n1397 VGND.n1379 2.1509
R3834 VGND.n2243 VGND.n2242 2.1509
R3835 VGND.n201 VGND.n176 2.1509
R3836 VGND.n2102 VGND.n2101 2.13383
R3837 VGND.n2151 VGND.n2150 2.13383
R3838 VGND.n1117 VGND.n352 2.13383
R3839 VGND.n1067 VGND.n432 2.13383
R3840 VGND.n1547 VGND.n1546 2.13383
R3841 VGND.n1265 VGND.n1183 2.13383
R3842 VGND.n1464 VGND.n1352 2.13383
R3843 VGND.n2206 VGND.n2205 2.13383
R3844 VGND.n257 VGND.n256 2.13383
R3845 VGND.n1160 VGND.n144 2.08643
R3846 VGND.n2302 VGND.n1671 2.08643
R3847 VGND.n1777 VGND.n1776 2.08643
R3848 VGND.n2144 VGND.n1884 2.08643
R3849 VGND.n103 VGND.n101 2.08643
R3850 VGND.n353 VGND.n76 2.08643
R3851 VGND.n2101 VGND.n2100 1.9461
R3852 VGND.n2150 VGND.n2149 1.9461
R3853 VGND.n1120 VGND.n1117 1.9461
R3854 VGND.n1068 VGND.n1067 1.9461
R3855 VGND.n1546 VGND.n1545 1.9461
R3856 VGND.n1292 VGND.n1183 1.9461
R3857 VGND.n1464 VGND.n1463 1.9461
R3858 VGND.n2205 VGND.n2204 1.9461
R3859 VGND.n256 VGND.n255 1.9461
R3860 VGND.n2374 VGND.n6 1.70675
R3861 VGND.n2370 VGND.n9 1.70675
R3862 VGND.n2366 VGND.n12 1.70675
R3863 VGND.n2362 VGND.n15 1.70675
R3864 VGND.n2378 VGND.n2 1.70675
R3865 VGND.n2381 VGND.n2 1.706
R3866 VGND.n2377 VGND.n6 1.706
R3867 VGND.n2373 VGND.n9 1.706
R3868 VGND.n2369 VGND.n12 1.706
R3869 VGND.n2365 VGND.n15 1.706
R3870 VGND.n2379 VGND.n1 1.70307
R3871 VGND.n2375 VGND.n5 1.70307
R3872 VGND.n2371 VGND.n8 1.70307
R3873 VGND.n2367 VGND.n11 1.70307
R3874 VGND.n2363 VGND.n14 1.70307
R3875 VGND.n2355 VGND.n2353 1.70248
R3876 VGND.n2361 VGND.n2354 1.70149
R3877 VGND.n2092 VGND.n1963 1.47392
R3878 VGND.n434 VGND.n433 1.47392
R3879 VGND.n1591 VGND.n1590 1.47392
R3880 VGND.n1351 VGND.n1302 1.47392
R3881 VGND.n2253 VGND.n2252 1.47392
R3882 VGND.n2347 VGND.n2346 1.47392
R3883 VGND.n966 VGND.n965 1.20883
R3884 VGND.n2366 VGND.n2365 1.20488
R3885 VGND.n966 VGND.n962 1.14633
R3886 VGND.n943 VGND.n941 1.063
R3887 VGND.n926 VGND.n664 1.03175
R3888 VGND.n921 VGND.n919 0.891125
R3889 VGND.n907 VGND.n905 0.859875
R3890 VGND.n915 VGND.n913 0.859875
R3891 VGND.n892 VGND.n891 0.819774
R3892 VGND.n876 VGND.n875 0.819774
R3893 VGND.n879 VGND.n878 0.819774
R3894 VGND.n2109 VGND.n1901 0.8197
R3895 VGND.n2108 VGND.n1899 0.8197
R3896 VGND.n2115 VGND.n1898 0.8197
R3897 VGND.n2117 VGND.n2116 0.8197
R3898 VGND.n2124 VGND.n1896 0.8197
R3899 VGND.n2123 VGND.n1894 0.8197
R3900 VGND.n2130 VGND.n1893 0.8197
R3901 VGND.n2132 VGND.n2131 0.8197
R3902 VGND.n2139 VGND.n1889 0.8197
R3903 VGND.n2158 VGND.n1822 0.8197
R3904 VGND.n2157 VGND.n1820 0.8197
R3905 VGND.n2164 VGND.n1819 0.8197
R3906 VGND.n2166 VGND.n2165 0.8197
R3907 VGND.n2173 VGND.n1817 0.8197
R3908 VGND.n2172 VGND.n1815 0.8197
R3909 VGND.n2179 VGND.n1814 0.8197
R3910 VGND.n2181 VGND.n2180 0.8197
R3911 VGND.n2188 VGND.n1810 0.8197
R3912 VGND.n1121 VGND.n288 0.8197
R3913 VGND.n1126 VGND.n1125 0.8197
R3914 VGND.n1129 VGND.n287 0.8197
R3915 VGND.n1133 VGND.n1132 0.8197
R3916 VGND.n285 VGND.n284 0.8197
R3917 VGND.n1140 VGND.n1139 0.8197
R3918 VGND.n1143 VGND.n283 0.8197
R3919 VGND.n1145 VGND.n1144 0.8197
R3920 VGND.n1153 VGND.n279 0.8197
R3921 VGND.n1093 VGND.n1092 0.8197
R3922 VGND.n1089 VGND.n1088 0.8197
R3923 VGND.n1085 VGND.n1069 0.8197
R3924 VGND.n1084 VGND.n1081 0.8197
R3925 VGND.n1078 VGND.n1070 0.8197
R3926 VGND.n1077 VGND.n1074 0.8197
R3927 VGND.n1071 VGND.n360 0.8197
R3928 VGND.n1099 VGND.n1098 0.8197
R3929 VGND.n1102 VGND.n359 0.8197
R3930 VGND.n1554 VGND.n1483 0.8197
R3931 VGND.n1553 VGND.n1480 0.8197
R3932 VGND.n1560 VGND.n1479 0.8197
R3933 VGND.n1562 VGND.n1561 0.8197
R3934 VGND.n1569 VGND.n1477 0.8197
R3935 VGND.n1568 VGND.n1475 0.8197
R3936 VGND.n1575 VGND.n1474 0.8197
R3937 VGND.n1577 VGND.n1576 0.8197
R3938 VGND.n1584 VGND.n1470 0.8197
R3939 VGND.n1291 VGND.n1184 0.8197
R3940 VGND.n1288 VGND.n1287 0.8197
R3941 VGND.n1284 VGND.n1187 0.8197
R3942 VGND.n1283 VGND.n1188 0.8197
R3943 VGND.n1212 VGND.n1209 0.8197
R3944 VGND.n1217 VGND.n1214 0.8197
R3945 VGND.n1218 VGND.n1208 0.8197
R3946 VGND.n1222 VGND.n1221 0.8197
R3947 VGND.n1226 VGND.n1225 0.8197
R3948 VGND.n1462 VGND.n1354 0.8197
R3949 VGND.n1459 VGND.n1458 0.8197
R3950 VGND.n1455 VGND.n1357 0.8197
R3951 VGND.n1454 VGND.n1358 0.8197
R3952 VGND.n1384 VGND.n1381 0.8197
R3953 VGND.n1389 VGND.n1386 0.8197
R3954 VGND.n1390 VGND.n1380 0.8197
R3955 VGND.n1394 VGND.n1393 0.8197
R3956 VGND.n1398 VGND.n1397 0.8197
R3957 VGND.n2213 VGND.n1714 0.8197
R3958 VGND.n2212 VGND.n1712 0.8197
R3959 VGND.n2219 VGND.n1711 0.8197
R3960 VGND.n2221 VGND.n2220 0.8197
R3961 VGND.n2228 VGND.n1709 0.8197
R3962 VGND.n2227 VGND.n1707 0.8197
R3963 VGND.n2234 VGND.n1706 0.8197
R3964 VGND.n2236 VGND.n2235 0.8197
R3965 VGND.n2243 VGND.n1702 0.8197
R3966 VGND.n263 VGND.n155 0.8197
R3967 VGND.n262 VGND.n156 0.8197
R3968 VGND.n181 VGND.n179 0.8197
R3969 VGND.n186 VGND.n183 0.8197
R3970 VGND.n187 VGND.n178 0.8197
R3971 VGND.n193 VGND.n190 0.8197
R3972 VGND.n194 VGND.n177 0.8197
R3973 VGND.n198 VGND.n197 0.8197
R3974 VGND.n202 VGND.n201 0.8197
R3975 VGND.n679 VGND.n678 0.813
R3976 VGND.n888 VGND.n887 0.813
R3977 VGND.n888 VGND.n0 0.813
R3978 VGND.n946 VGND.n945 0.734875
R3979 VGND.n935 VGND.n934 0.734875
R3980 VGND.n946 VGND.n932 0.71925
R3981 VGND.n727 VGND.n668 0.688
R3982 VGND.n690 VGND.n675 0.688
R3983 VGND.n785 VGND.n783 0.688
R3984 VGND.n805 VGND.n803 0.688
R3985 VGND.n828 VGND.n826 0.688
R3986 VGND.n941 VGND.n939 0.688
R3987 VGND.n728 VGND.n667 0.672375
R3988 VGND.n631 VGND.n580 0.65675
R3989 VGND.n698 VGND.n674 0.6255
R3990 VGND.n752 VGND.n744 0.6255
R3991 VGND.n754 VGND.n752 0.6255
R3992 VGND.n756 VGND.n754 0.6255
R3993 VGND.n735 VGND.n667 0.609875
R3994 VGND.n932 VGND.n931 0.547375
R3995 VGND.n629 VGND.n628 0.542167
R3996 VGND.n937 VGND.n935 0.53175
R3997 VGND.n728 VGND.n727 0.516125
R3998 VGND.n691 VGND.n690 0.516125
R3999 VGND.n691 VGND.n674 0.516125
R4000 VGND.n928 VGND.n926 0.516125
R4001 VGND.n786 VGND.n785 0.5005
R4002 VGND.n803 VGND.n786 0.5005
R4003 VGND.n806 VGND.n805 0.5005
R4004 VGND.n826 VGND.n806 0.5005
R4005 VGND.n954 VGND.n581 0.472458
R4006 VGND.n720 VGND.n668 0.46925
R4007 VGND.n719 VGND.n718 0.46925
R4008 VGND.n670 VGND.n669 0.46925
R4009 VGND.n700 VGND.n699 0.46925
R4010 VGND.n703 VGND.n702 0.46925
R4011 VGND.n908 VGND.n907 0.438
R4012 VGND.n913 VGND.n911 0.438
R4013 VGND.n678 VGND.n675 0.40675
R4014 VGND.n922 VGND.n921 0.40675
R4015 VGND.n908 VGND.n903 0.391125
R4016 VGND.n911 VGND.n666 0.391125
R4017 VGND.n922 VGND.n917 0.391125
R4018 VGND.n931 VGND.n930 0.391125
R4019 VGND.n852 VGND.n851 0.3755
R4020 VGND.n704 VGND.n703 0.359875
R4021 VGND.n720 VGND.n719 0.34425
R4022 VGND.n718 VGND.n717 0.34425
R4023 VGND.n671 VGND.n670 0.34425
R4024 VGND.n669 VGND.n7 0.34425
R4025 VGND.n699 VGND.n698 0.34425
R4026 VGND.n701 VGND.n700 0.34425
R4027 VGND.n702 VGND.n10 0.34425
R4028 VGND.n829 VGND.n828 0.34425
R4029 VGND.n903 VGND.n901 0.34425
R4030 VGND.n905 VGND.n666 0.34425
R4031 VGND.n917 VGND.n915 0.34425
R4032 VGND.n919 VGND.n664 0.34425
R4033 VGND.n930 VGND.n928 0.34425
R4034 VGND.n945 VGND.n943 0.34425
R4035 VGND.n939 VGND.n937 0.34425
R4036 VGND.n934 VGND.n4 0.34425
R4037 VGND.n862 VGND.n744 0.313
R4038 VGND.n851 VGND.n849 0.313
R4039 VGND.n2378 VGND.n2377 0.29425
R4040 VGND.n2352 VGND.n16 0.28175
R4041 VGND.n893 VGND.n892 0.279967
R4042 VGND.n889 VGND.n876 0.279967
R4043 VGND.n886 VGND.n879 0.279967
R4044 VGND.n2374 VGND.n2373 0.26605
R4045 VGND.n717 VGND.n671 0.2505
R4046 VGND.n852 VGND.n756 0.2505
R4047 VGND.n704 VGND.n701 0.234875
R4048 VGND.n867 VGND.n581 0.233542
R4049 VGND.n965 VGND.n16 0.224458
R4050 VGND.n831 VGND.n830 0.188
R4051 VGND.n779 VGND.n763 0.188
R4052 VGND.n624 VGND.n623 0.188
R4053 VGND.n626 VGND.n601 0.188
R4054 VGND.n962 VGND.n961 0.188
R4055 VGND.n867 VGND.n13 0.159125
R4056 VGND.n835 VGND.n831 0.15675
R4057 VGND.n779 VGND.n778 0.15675
R4058 VGND.n2382 VGND.n2381 0.13993
R4059 VGND.n955 VGND.n954 0.13302
R4060 VGND.n615 VGND.n614 0.1255
R4061 VGND.n622 VGND.n604 0.1255
R4062 VGND.n967 VGND.n578 0.1255
R4063 VGND.n2362 VGND.n2361 0.06865
R4064 VGND.n615 VGND.n611 0.0626438
R4065 VGND.n604 VGND.n603 0.0626438
R4066 VGND.n964 VGND.n578 0.0626438
R4067 VGND VGND.n2382 0.0600243
R4068 VGND.n815 VGND.n814 0.0451429
R4069 VGND.n814 VGND.n810 0.0451429
R4070 VGND.n795 VGND.n794 0.0451429
R4071 VGND.n795 VGND.n790 0.0451429
R4072 VGND.n626 VGND.n600 0.0421667
R4073 VGND.n2370 VGND.n2369 0.029875
R4074 VGND.n2375 VGND.n6 0.0256998
R4075 VGND.n2371 VGND.n9 0.0256998
R4076 VGND.n2367 VGND.n12 0.0256998
R4077 VGND.n2363 VGND.n15 0.0256998
R4078 VGND.n2379 VGND.n2 0.0256998
R4079 VGND.n634 VGND.n595 0.0217373
R4080 VGND.n630 VGND.n596 0.0217373
R4081 VGND.n628 VGND.n627 0.0217373
R4082 VGND.n625 VGND.n602 0.0217373
R4083 VGND.n597 VGND.n595 0.0217373
R4084 VGND.n630 VGND.n629 0.0217373
R4085 VGND.n627 VGND.n599 0.0217373
R4086 VGND.n602 VGND.n599 0.0217373
R4087 VGND.n632 VGND.n597 0.0217373
R4088 VGND.n633 VGND.n596 0.0217373
R4089 VGND.n632 VGND.n631 0.0217373
R4090 VGND.n624 VGND.n598 0.0217373
R4091 VGND.n600 VGND.n598 0.0217373
R4092 VGND.n2376 VGND.n2375 0.0200833
R4093 VGND.n2372 VGND.n2371 0.0200833
R4094 VGND.n2368 VGND.n2367 0.0200833
R4095 VGND.n2364 VGND.n2363 0.0200833
R4096 VGND.n2380 VGND.n2379 0.0200833
R4097 VGND.n2358 VGND.n2355 0.0185769
R4098 VGND.n2360 VGND.n2355 0.0185769
R4099 VGND.n2358 VGND.n2354 0.0100146
R4100 VGND.n2357 VGND.n2354 0.0100146
R4101 VGND.n2361 VGND.n2353 0.00803545
R4102 VGND.n2359 VGND.n2353 0.00803545
R4103 VGND.n2365 VGND.n14 0.0068649
R4104 VGND.n2369 VGND.n11 0.0068649
R4105 VGND.n2373 VGND.n8 0.0068649
R4106 VGND.n2377 VGND.n5 0.0068649
R4107 VGND.n2381 VGND.n1 0.0068649
R4108 VGND.n2378 VGND.n1 0.0068649
R4109 VGND.n2374 VGND.n5 0.0068649
R4110 VGND.n2370 VGND.n8 0.0068649
R4111 VGND.n2366 VGND.n11 0.0068649
R4112 VGND.n2362 VGND.n14 0.0068649
R4113 V_CONT.n25 V_CONT.t14 404.683
R4114 V_CONT.n25 V_CONT.t9 403.755
R4115 V_CONT.n26 V_CONT.t12 403.755
R4116 V_CONT.n27 V_CONT.t10 396.866
R4117 V_CONT.n12 V_CONT.t13 377.567
R4118 V_CONT.n11 V_CONT.t8 297.233
R4119 V_CONT.n13 V_CONT.n11 232.001
R4120 V_CONT.n13 V_CONT.n12 228.2
R4121 V_CONT.n12 V_CONT.t11 216.9
R4122 V_CONT.n7 V_CONT.t4 163.706
R4123 V_CONT.n22 V_CONT.n21 158.589
R4124 V_CONT.n22 V_CONT.n20 148.901
R4125 V_CONT.n11 V_CONT.t15 136.567
R4126 V_CONT.n23 V_CONT.n19 49.3391
R4127 V_CONT.n20 V_CONT.t1 24.6255
R4128 V_CONT.n20 V_CONT.t2 24.6255
R4129 V_CONT.n21 V_CONT.t3 24.6255
R4130 V_CONT.n21 V_CONT.t6 24.6255
R4131 V_CONT.n14 V_CONT.n13 16.3148
R4132 V_CONT.n19 V_CONT.t0 15.0005
R4133 V_CONT.n19 V_CONT.t7 15.0005
R4134 V_CONT.n24 V_CONT.n23 11.461
R4135 V_CONT.n7 V_CONT.t5 6.75823
R4136 V_CONT.n17 V_CONT.n16 4.5005
R4137 V_CONT.n9 V_CONT.n5 4.5005
R4138 V_CONT.n17 V_CONT.n5 4.5005
R4139 V_CONT.n18 V_CONT.n1 4.5005
R4140 V_CONT.n18 V_CONT.n3 4.5005
R4141 V_CONT.n18 V_CONT.n17 4.5005
R4142 V_CONT.n16 V_CONT.n7 3.3845
R4143 V_CONT V_CONT.n27 2.68208
R4144 V_CONT.n15 V_CONT.n14 2.2458
R4145 V_CONT.n6 V_CONT.n0 2.2458
R4146 V_CONT.n18 V_CONT.n2 2.24063
R4147 V_CONT.n16 V_CONT.n10 2.24063
R4148 V_CONT.n16 V_CONT.n8 2.24063
R4149 V_CONT.n5 V_CONT.n4 2.24063
R4150 V_CONT V_CONT.n24 1.13071
R4151 V_CONT.n27 V_CONT.n26 1.01121
R4152 V_CONT.n26 V_CONT.n25 0.929071
R4153 V_CONT.n23 V_CONT.n22 0.438
R4154 V_CONT.n24 V_CONT.n18 0.336438
R4155 V_CONT.n17 V_CONT.n6 0.0421667
R4156 V_CONT.n14 V_CONT.n2 0.0217373
R4157 V_CONT.n9 V_CONT.n2 0.0217373
R4158 V_CONT.n8 V_CONT.n6 0.0217373
R4159 V_CONT.n4 V_CONT.n1 0.0217373
R4160 V_CONT.n10 V_CONT.n1 0.0217373
R4161 V_CONT.n10 V_CONT.n9 0.0217373
R4162 V_CONT.n8 V_CONT.n3 0.0217373
R4163 V_CONT.n4 V_CONT.n3 0.0217373
R4164 V_CONT.n15 V_CONT.n5 0.0113926
R4165 V_CONT.n16 V_CONT.n15 0.0113926
R4166 V_CONT.n18 V_CONT.n0 0.0113926
R4167 V_CONT.n5 V_CONT.n0 0.0113926
R4168 a_11860_6640.t5 a_11860_6640.t6 835.467
R4169 a_11860_6640.n2 a_11860_6640.t5 560.011
R4170 a_11860_6640.n0 a_11860_6640.t8 517.347
R4171 a_11860_6640.n1 a_11860_6640.t4 514.134
R4172 a_11860_6640.n2 a_11860_6640.n1 491.791
R4173 a_11860_6640.n3 a_11860_6640.n0 363.2
R4174 a_11860_6640.n1 a_11860_6640.t3 273.134
R4175 a_11860_6640.n5 a_11860_6640.n4 244.716
R4176 a_11860_6640.n0 a_11860_6640.t7 228.148
R4177 a_11860_6640.t1 a_11860_6640.n5 221.411
R4178 a_11860_6640.n5 a_11860_6640.n3 54.3734
R4179 a_11860_6640.n3 a_11860_6640.n2 37.6567
R4180 a_11860_6640.n4 a_11860_6640.t0 24.0005
R4181 a_11860_6640.n4 a_11860_6640.t2 24.0005
R4182 a_14930_6670.t0 a_14930_6670.n1 203.528
R4183 a_14930_6670.n0 a_14930_6670.t2 203.528
R4184 a_14930_6670.n0 a_14930_6670.t1 183.935
R4185 a_14930_6670.n1 a_14930_6670.t3 183.935
R4186 a_14930_6670.n1 a_14930_6670.n0 83.2005
R4187 a_17714_9374.n0 a_17714_9374.t8 486.438
R4188 a_17714_9374.n8 a_17714_9374.t10 377.567
R4189 a_17714_9374.n1 a_17714_9374.t11 377.567
R4190 a_17714_9374.n9 a_17714_9374.n8 257.067
R4191 a_17714_9374.n7 a_17714_9374.n6 257.067
R4192 a_17714_9374.n2 a_17714_9374.n1 257.067
R4193 a_17714_9374.n5 a_17714_9374.n4 161.3
R4194 a_17714_9374.n11 a_17714_9374.n10 161.3
R4195 a_17714_9374.n8 a_17714_9374.t9 120.501
R4196 a_17714_9374.n9 a_17714_9374.t6 120.501
R4197 a_17714_9374.n7 a_17714_9374.t0 120.501
R4198 a_17714_9374.n6 a_17714_9374.t4 120.501
R4199 a_17714_9374.n1 a_17714_9374.t12 120.501
R4200 a_17714_9374.n2 a_17714_9374.t2 120.501
R4201 a_17714_9374.n4 a_17714_9374.n3 119.237
R4202 a_17714_9374.n12 a_17714_9374.n11 119.237
R4203 a_17714_9374.n10 a_17714_9374.n9 85.6894
R4204 a_17714_9374.n10 a_17714_9374.n7 85.6894
R4205 a_17714_9374.n6 a_17714_9374.n5 85.6894
R4206 a_17714_9374.n5 a_17714_9374.n2 85.6894
R4207 a_17714_9374.n3 a_17714_9374.t3 19.7005
R4208 a_17714_9374.n3 a_17714_9374.t5 19.7005
R4209 a_17714_9374.t1 a_17714_9374.n12 19.7005
R4210 a_17714_9374.n12 a_17714_9374.t7 19.7005
R4211 a_17714_9374.n4 a_17714_9374.n0 5.1255
R4212 a_17714_9374.n11 a_17714_9374.n0 4.5005
R4213 a_18160_10940.n11 a_18160_10940.t3 384.967
R4214 a_18160_10940.n3 a_18160_10940.t1 384.967
R4215 a_18160_10940.t5 a_18160_10940.n11 378.358
R4216 a_18160_10940.n3 a_18160_10940.t2 375.896
R4217 a_18160_10940.n10 a_18160_10940.n0 313.846
R4218 a_18160_10940.n9 a_18160_10940.n1 313.846
R4219 a_18160_10940.n4 a_18160_10940.n2 313
R4220 a_18160_10940.n7 a_18160_10940.n6 130.143
R4221 a_18160_10940.n7 a_18160_10940.n5 119.267
R4222 a_18160_10940.n10 a_18160_10940.n9 83.2005
R4223 a_18160_10940.t2 a_18160_10940.n2 49.2505
R4224 a_18160_10940.n2 a_18160_10940.t10 49.2505
R4225 a_18160_10940.n0 a_18160_10940.t11 49.2505
R4226 a_18160_10940.n0 a_18160_10940.t4 49.2505
R4227 a_18160_10940.n1 a_18160_10940.t0 49.2505
R4228 a_18160_10940.n1 a_18160_10940.t12 49.2505
R4229 a_18160_10940.n8 a_18160_10940.n4 49.0672
R4230 a_18160_10940.n5 a_18160_10940.t6 19.7005
R4231 a_18160_10940.n5 a_18160_10940.t7 19.7005
R4232 a_18160_10940.n6 a_18160_10940.t8 19.7005
R4233 a_18160_10940.n6 a_18160_10940.t9 19.7005
R4234 a_18160_10940.n9 a_18160_10940.n8 17.0672
R4235 a_18160_10940.n4 a_18160_10940.n3 16.0005
R4236 a_18160_10940.n11 a_18160_10940.n10 16.0005
R4237 a_18160_10940.n8 a_18160_10940.n7 9.69113
R4238 VDPWR.n150 VDPWR.n149 6615
R4239 VDPWR.n178 VDPWR.n149 6495
R4240 VDPWR.n178 VDPWR.n148 4995
R4241 VDPWR.n175 VDPWR.n148 2985
R4242 VDPWR.t74 VDPWR.t125 2804.76
R4243 VDPWR.t153 VDPWR.t89 2533.33
R4244 VDPWR.t161 VDPWR.t384 2307.14
R4245 VDPWR.t242 VDPWR.t399 2216.67
R4246 VDPWR.t214 VDPWR.t337 2216.67
R4247 VDPWR.t371 VDPWR.t167 2216.67
R4248 VDPWR.t351 VDPWR.t395 2126.19
R4249 VDPWR.t61 VDPWR.t407 1538.1
R4250 VDPWR.t169 VDPWR.t36 1492.86
R4251 VDPWR.t14 VDPWR.t71 1492.86
R4252 VDPWR.n45 VDPWR.t367 1289.29
R4253 VDPWR.n46 VDPWR.t369 1289.29
R4254 VDPWR.t0 VDPWR.t113 1130.95
R4255 VDPWR.t201 VDPWR.t322 1130.95
R4256 VDPWR.t65 VDPWR.t157 1130.95
R4257 VDPWR.t72 VDPWR.t209 1130.95
R4258 VDPWR.t409 VDPWR.t182 1130.95
R4259 VDPWR.n13 VDPWR.t380 927.381
R4260 VDPWR.n14 VDPWR.t80 927.381
R4261 VDPWR.n25 VDPWR.t63 927.381
R4262 VDPWR.n26 VDPWR.t216 927.381
R4263 VDPWR.n204 VDPWR.n195 831.25
R4264 VDPWR.n198 VDPWR.n197 831.25
R4265 VDPWR.n378 VDPWR.n192 831.25
R4266 VDPWR.n373 VDPWR.n372 831.25
R4267 VDPWR.n34 VDPWR.t410 740.534
R4268 VDPWR.n33 VDPWR.t396 740.534
R4269 VDPWR.t321 VDPWR.n503 708.125
R4270 VDPWR.n526 VDPWR.t321 708.125
R4271 VDPWR.n523 VDPWR.t277 708.125
R4272 VDPWR.t277 VDPWR.n504 708.125
R4273 VDPWR.t253 VDPWR.n483 708.125
R4274 VDPWR.n536 VDPWR.t253 708.125
R4275 VDPWR.n533 VDPWR.t262 708.125
R4276 VDPWR.t262 VDPWR.n484 708.125
R4277 VDPWR.t298 VDPWR.n606 708.125
R4278 VDPWR.n613 VDPWR.t298 708.125
R4279 VDPWR.t295 VDPWR.n633 708.125
R4280 VDPWR.n649 VDPWR.t295 708.125
R4281 VDPWR.t288 VDPWR.n620 708.125
R4282 VDPWR.n659 VDPWR.t288 708.125
R4283 VDPWR.n151 VDPWR.n147 705.601
R4284 VDPWR.n610 VDPWR.t256 694.444
R4285 VDPWR.t256 VDPWR.n607 694.444
R4286 VDPWR.n179 VDPWR.n147 692.801
R4287 VDPWR.n12 VDPWR.t400 663.801
R4288 VDPWR.n47 VDPWR.t245 663.801
R4289 VDPWR.n44 VDPWR.t126 663.801
R4290 VDPWR.n27 VDPWR.t162 663.801
R4291 VDPWR.n24 VDPWR.t168 663.801
R4292 VDPWR.n15 VDPWR.t215 663.801
R4293 VDPWR.n8 VDPWR.n6 662.297
R4294 VDPWR.n1 VDPWR.n0 661.734
R4295 VDPWR.n40 VDPWR.n39 661.734
R4296 VDPWR.n38 VDPWR.n37 661.734
R4297 VDPWR.n36 VDPWR.n35 661.734
R4298 VDPWR.n32 VDPWR.n31 661.734
R4299 VDPWR.n30 VDPWR.n29 661.734
R4300 VDPWR.n3 VDPWR.n2 661.734
R4301 VDPWR.n22 VDPWR.n21 661.734
R4302 VDPWR.n20 VDPWR.n19 661.734
R4303 VDPWR.n18 VDPWR.n17 661.734
R4304 VDPWR.n5 VDPWR.n4 661.734
R4305 VDPWR.n10 VDPWR.n9 661.734
R4306 VDPWR.n8 VDPWR.n7 661.734
R4307 VDPWR.n42 VDPWR.n41 660.514
R4308 VDPWR.n525 VDPWR.t320 657.76
R4309 VDPWR.n535 VDPWR.t252 657.76
R4310 VDPWR.n612 VDPWR.t297 640.794
R4311 VDPWR.n648 VDPWR.t294 640.794
R4312 VDPWR.n658 VDPWR.t287 640.794
R4313 VDPWR.t399 VDPWR.n13 610.715
R4314 VDPWR.n14 VDPWR.t214 610.715
R4315 VDPWR.t167 VDPWR.n25 610.715
R4316 VDPWR.n26 VDPWR.t161 610.715
R4317 VDPWR.t125 VDPWR.n45 610.715
R4318 VDPWR.n46 VDPWR.t244 610.715
R4319 VDPWR.n559 VDPWR.n557 587.407
R4320 VDPWR.n563 VDPWR.n560 587.407
R4321 VDPWR.n589 VDPWR.n588 587.407
R4322 VDPWR.n584 VDPWR.n550 587.407
R4323 VDPWR.n473 VDPWR.n472 585
R4324 VDPWR.n452 VDPWR.n417 585
R4325 VDPWR.n588 VDPWR.n587 585
R4326 VDPWR.n586 VDPWR.n584 585
R4327 VDPWR.n570 VDPWR.n559 585
R4328 VDPWR.n567 VDPWR.n560 585
R4329 VDPWR.n193 VDPWR.n192 585
R4330 VDPWR.n375 VDPWR.n373 585
R4331 VDPWR.n196 VDPWR.n195 585
R4332 VDPWR.n201 VDPWR.n198 585
R4333 VDPWR.n291 VDPWR.n227 585
R4334 VDPWR.n286 VDPWR.n227 585
R4335 VDPWR.n235 VDPWR.n228 585
R4336 VDPWR.n230 VDPWR.n228 585
R4337 VDPWR.n282 VDPWR.n237 585
R4338 VDPWR.n275 VDPWR.n237 585
R4339 VDPWR.n272 VDPWR.n244 585
R4340 VDPWR.n267 VDPWR.n244 585
R4341 VDPWR.n252 VDPWR.n245 585
R4342 VDPWR.n247 VDPWR.n245 585
R4343 VDPWR.n264 VDPWR.n253 585
R4344 VDPWR.n260 VDPWR.n253 585
R4345 VDPWR.n104 VDPWR.n53 585
R4346 VDPWR.n108 VDPWR.n53 585
R4347 VDPWR.n97 VDPWR.n59 585
R4348 VDPWR.n88 VDPWR.n59 585
R4349 VDPWR.n77 VDPWR.n76 585
R4350 VDPWR.n77 VDPWR.n64 585
R4351 VDPWR.t255 VDPWR.n611 557.783
R4352 VDPWR.t276 VDPWR.n524 540.818
R4353 VDPWR.t261 VDPWR.n534 540.818
R4354 VDPWR.t300 VDPWR.n647 523.855
R4355 VDPWR.t317 VDPWR.n657 523.855
R4356 VDPWR.t113 VDPWR.t176 497.62
R4357 VDPWR.t380 VDPWR.t0 497.62
R4358 VDPWR.t322 VDPWR.t242 497.62
R4359 VDPWR.t80 VDPWR.t201 497.62
R4360 VDPWR.t337 VDPWR.t65 497.62
R4361 VDPWR.t157 VDPWR.t63 497.62
R4362 VDPWR.t209 VDPWR.t371 497.62
R4363 VDPWR.t216 VDPWR.t72 497.62
R4364 VDPWR.t384 VDPWR.t169 497.62
R4365 VDPWR.t36 VDPWR.t351 497.62
R4366 VDPWR.t395 VDPWR.t409 497.62
R4367 VDPWR.t182 VDPWR.t61 497.62
R4368 VDPWR.t407 VDPWR.t367 497.62
R4369 VDPWR.t149 VDPWR.t74 497.62
R4370 VDPWR.t71 VDPWR.t149 497.62
R4371 VDPWR.t89 VDPWR.t14 497.62
R4372 VDPWR.t369 VDPWR.t153 497.62
R4373 VDPWR.n203 VDPWR.t378 465.079
R4374 VDPWR.t378 VDPWR.n202 465.079
R4375 VDPWR.n377 VDPWR.t411 465.079
R4376 VDPWR.t411 VDPWR.n376 465.079
R4377 VDPWR.n338 VDPWR.t130 464.281
R4378 VDPWR.t130 VDPWR.n337 464.281
R4379 VDPWR.t140 VDPWR.n186 464.281
R4380 VDPWR.n382 VDPWR.t140 464.281
R4381 VDPWR.n392 VDPWR.t70 464.281
R4382 VDPWR.t70 VDPWR.n391 464.281
R4383 VDPWR.t35 VDPWR.n208 464.281
R4384 VDPWR.n352 VDPWR.t35 464.281
R4385 VDPWR.n362 VDPWR.t394 464.281
R4386 VDPWR.t394 VDPWR.n361 464.281
R4387 VDPWR.n347 VDPWR.t335 464.281
R4388 VDPWR.t335 VDPWR.n346 464.281
R4389 VDPWR.t25 VDPWR.n319 464.281
R4390 VDPWR.n322 VDPWR.t25 464.281
R4391 VDPWR.n314 VDPWR.t116 464.281
R4392 VDPWR.t116 VDPWR.n217 464.281
R4393 VDPWR.n307 VDPWR.t247 464.281
R4394 VDPWR.t247 VDPWR.n306 464.281
R4395 VDPWR.n297 VDPWR.t389 464.281
R4396 VDPWR.t389 VDPWR.n221 464.281
R4397 VDPWR.n127 VDPWR.t199 461.389
R4398 VDPWR.t199 VDPWR.n126 461.389
R4399 VDPWR.n121 VDPWR.t331 461.389
R4400 VDPWR.t331 VDPWR.n120 461.389
R4401 VDPWR.n143 VDPWR.t235 461.389
R4402 VDPWR.t235 VDPWR.n142 461.389
R4403 VDPWR.n137 VDPWR.t329 461.389
R4404 VDPWR.t329 VDPWR.n136 461.389
R4405 VDPWR.n168 VDPWR.t250 461.389
R4406 VDPWR.t250 VDPWR.n167 461.389
R4407 VDPWR.n162 VDPWR.t327 461.389
R4408 VDPWR.t327 VDPWR.n161 461.389
R4409 VDPWR.n615 VDPWR.t296 422.384
R4410 VDPWR.n608 VDPWR.t254 422.384
R4411 VDPWR.n117 VDPWR.t426 420.111
R4412 VDPWR.n133 VDPWR.t427 420.111
R4413 VDPWR.n158 VDPWR.t428 420.111
R4414 VDPWR.n651 VDPWR.t293 418.368
R4415 VDPWR.n644 VDPWR.t299 418.368
R4416 VDPWR.n661 VDPWR.t286 418.368
R4417 VDPWR.n654 VDPWR.t316 418.368
R4418 VDPWR.n236 VDPWR.t430 411.101
R4419 VDPWR.t320 VDPWR.t345 407.144
R4420 VDPWR.t345 VDPWR.t196 407.144
R4421 VDPWR.t196 VDPWR.t20 407.144
R4422 VDPWR.t20 VDPWR.t403 407.144
R4423 VDPWR.t403 VDPWR.t192 407.144
R4424 VDPWR.t192 VDPWR.t10 407.144
R4425 VDPWR.t10 VDPWR.t325 407.144
R4426 VDPWR.t325 VDPWR.t357 407.144
R4427 VDPWR.t357 VDPWR.t76 407.144
R4428 VDPWR.t76 VDPWR.t178 407.144
R4429 VDPWR.t178 VDPWR.t147 407.144
R4430 VDPWR.t147 VDPWR.t343 407.144
R4431 VDPWR.t343 VDPWR.t220 407.144
R4432 VDPWR.t220 VDPWR.t12 407.144
R4433 VDPWR.t12 VDPWR.t205 407.144
R4434 VDPWR.t205 VDPWR.t127 407.144
R4435 VDPWR.t127 VDPWR.t59 407.144
R4436 VDPWR.t59 VDPWR.t180 407.144
R4437 VDPWR.t180 VDPWR.t276 407.144
R4438 VDPWR.t252 VDPWR.t8 407.144
R4439 VDPWR.t8 VDPWR.t401 407.144
R4440 VDPWR.t401 VDPWR.t203 407.144
R4441 VDPWR.t203 VDPWR.t412 407.144
R4442 VDPWR.t412 VDPWR.t194 407.144
R4443 VDPWR.t194 VDPWR.t186 407.144
R4444 VDPWR.t186 VDPWR.t42 407.144
R4445 VDPWR.t42 VDPWR.t188 407.144
R4446 VDPWR.t188 VDPWR.t18 407.144
R4447 VDPWR.t18 VDPWR.t111 407.144
R4448 VDPWR.t111 VDPWR.t375 407.144
R4449 VDPWR.t375 VDPWR.t184 407.144
R4450 VDPWR.t184 VDPWR.t84 407.144
R4451 VDPWR.t84 VDPWR.t3 407.144
R4452 VDPWR.t3 VDPWR.t145 407.144
R4453 VDPWR.t145 VDPWR.t236 407.144
R4454 VDPWR.t236 VDPWR.t57 407.144
R4455 VDPWR.t57 VDPWR.t421 407.144
R4456 VDPWR.t421 VDPWR.t261 407.144
R4457 VDPWR.n457 VDPWR.t266 384.967
R4458 VDPWR.n461 VDPWR.t306 384.967
R4459 VDPWR.n424 VDPWR.t272 384.967
R4460 VDPWR.n428 VDPWR.t282 384.967
R4461 VDPWR.n47 VDPWR.n46 382.8
R4462 VDPWR.n45 VDPWR.n44 382.8
R4463 VDPWR.n27 VDPWR.n26 382.8
R4464 VDPWR.n25 VDPWR.n24 382.8
R4465 VDPWR.n15 VDPWR.n14 382.8
R4466 VDPWR.n13 VDPWR.n12 382.8
R4467 VDPWR.t297 VDPWR.t398 373.214
R4468 VDPWR.t398 VDPWR.t397 373.214
R4469 VDPWR.t397 VDPWR.t255 373.214
R4470 VDPWR.t294 VDPWR.t51 373.214
R4471 VDPWR.t51 VDPWR.t365 373.214
R4472 VDPWR.t365 VDPWR.t224 373.214
R4473 VDPWR.t224 VDPWR.t163 373.214
R4474 VDPWR.t163 VDPWR.t171 373.214
R4475 VDPWR.t171 VDPWR.t38 373.214
R4476 VDPWR.t38 VDPWR.t134 373.214
R4477 VDPWR.t134 VDPWR.t222 373.214
R4478 VDPWR.t222 VDPWR.t141 373.214
R4479 VDPWR.t141 VDPWR.t419 373.214
R4480 VDPWR.t419 VDPWR.t300 373.214
R4481 VDPWR.t287 VDPWR.t53 373.214
R4482 VDPWR.t53 VDPWR.t143 373.214
R4483 VDPWR.t143 VDPWR.t353 373.214
R4484 VDPWR.t353 VDPWR.t363 373.214
R4485 VDPWR.t363 VDPWR.t173 373.214
R4486 VDPWR.t173 VDPWR.t40 373.214
R4487 VDPWR.t40 VDPWR.t136 373.214
R4488 VDPWR.t136 VDPWR.t417 373.214
R4489 VDPWR.t417 VDPWR.t165 373.214
R4490 VDPWR.t165 VDPWR.t355 373.214
R4491 VDPWR.t355 VDPWR.t317 373.214
R4492 VDPWR.n528 VDPWR.t319 370.168
R4493 VDPWR.n521 VDPWR.t275 370.168
R4494 VDPWR.n538 VDPWR.t251 370.168
R4495 VDPWR.n531 VDPWR.t260 370.168
R4496 VDPWR.n442 VDPWR.t257 362.134
R4497 VDPWR.n541 VDPWR.t269 360.868
R4498 VDPWR.n595 VDPWR.t263 360.868
R4499 VDPWR.t314 VDPWR.t117 360.346
R4500 VDPWR.t117 VDPWR.t138 360.346
R4501 VDPWR.t138 VDPWR.t155 360.346
R4502 VDPWR.t155 VDPWR.t361 360.346
R4503 VDPWR.t361 VDPWR.t279 360.346
R4504 VDPWR.t382 VDPWR.t311 360.346
R4505 VDPWR.t339 VDPWR.t382 360.346
R4506 VDPWR.t341 VDPWR.t339 360.346
R4507 VDPWR.t123 VDPWR.t341 360.346
R4508 VDPWR.t290 VDPWR.t123 360.346
R4509 VDPWR.n478 VDPWR.t302 352.834
R4510 VDPWR.n635 VDPWR.t301 351.793
R4511 VDPWR.n622 VDPWR.t318 351.793
R4512 VDPWR.n180 VDPWR.n179 344
R4513 VDPWR.n74 VDPWR.t314 343.966
R4514 VDPWR.n99 VDPWR.t279 343.966
R4515 VDPWR.t311 VDPWR.n99 343.966
R4516 VDPWR.n106 VDPWR.t290 343.966
R4517 VDPWR.n462 VDPWR.t309 341.752
R4518 VDPWR.n456 VDPWR.t268 341.752
R4519 VDPWR.n427 VDPWR.t285 341.752
R4520 VDPWR.n423 VDPWR.t274 341.752
R4521 VDPWR.n57 VDPWR.t310 336.329
R4522 VDPWR.n57 VDPWR.t278 336.329
R4523 VDPWR.n62 VDPWR.t313 330
R4524 VDPWR.n110 VDPWR.t289 330
R4525 VDPWR.n430 VDPWR.n421 315.647
R4526 VDPWR.n429 VDPWR.n426 315.647
R4527 VDPWR.n425 VDPWR.n422 315.647
R4528 VDPWR.t2 VDPWR.t175 314.113
R4529 VDPWR.t55 VDPWR.t379 314.113
R4530 VDPWR.n459 VDPWR.n411 313.846
R4531 VDPWR.n460 VDPWR.n409 313.846
R4532 VDPWR.n458 VDPWR.n412 313.846
R4533 VDPWR.n214 VDPWR.t406 308.849
R4534 VDPWR.n423 VDPWR.t273 304.659
R4535 VDPWR.n643 VDPWR.n642 301.933
R4536 VDPWR.n641 VDPWR.n640 301.933
R4537 VDPWR.n639 VDPWR.n638 301.933
R4538 VDPWR.n637 VDPWR.n636 301.933
R4539 VDPWR.n632 VDPWR.n631 301.933
R4540 VDPWR.n630 VDPWR.n629 301.933
R4541 VDPWR.n628 VDPWR.n627 301.933
R4542 VDPWR.n626 VDPWR.n625 301.933
R4543 VDPWR.n624 VDPWR.n623 301.933
R4544 VDPWR.n619 VDPWR.n618 301.933
R4545 VDPWR.n520 VDPWR.n519 299.231
R4546 VDPWR.n518 VDPWR.n517 299.231
R4547 VDPWR.n516 VDPWR.n515 299.231
R4548 VDPWR.n514 VDPWR.n513 299.231
R4549 VDPWR.n512 VDPWR.n511 299.231
R4550 VDPWR.n510 VDPWR.n509 299.231
R4551 VDPWR.n508 VDPWR.n507 299.231
R4552 VDPWR.n506 VDPWR.n505 299.231
R4553 VDPWR.n502 VDPWR.n501 299.231
R4554 VDPWR.n500 VDPWR.n499 299.231
R4555 VDPWR.n498 VDPWR.n497 299.231
R4556 VDPWR.n496 VDPWR.n495 299.231
R4557 VDPWR.n494 VDPWR.n493 299.231
R4558 VDPWR.n492 VDPWR.n491 299.231
R4559 VDPWR.n490 VDPWR.n489 299.231
R4560 VDPWR.n488 VDPWR.n487 299.231
R4561 VDPWR.n486 VDPWR.n485 299.231
R4562 VDPWR.n482 VDPWR.n481 299.231
R4563 VDPWR.n84 VDPWR.n59 291.363
R4564 VDPWR.n96 VDPWR.n95 291.363
R4565 VDPWR.n95 VDPWR.n61 291.363
R4566 VDPWR.n472 VDPWR.n471 290.733
R4567 VDPWR.n472 VDPWR.n407 290.733
R4568 VDPWR.n420 VDPWR.n417 290.733
R4569 VDPWR.n445 VDPWR.n417 290.733
R4570 VDPWR.n289 VDPWR.n227 290.733
R4571 VDPWR.n229 VDPWR.n228 290.733
R4572 VDPWR.n276 VDPWR.n237 290.733
R4573 VDPWR.n270 VDPWR.n244 290.733
R4574 VDPWR.n246 VDPWR.n245 290.733
R4575 VDPWR.n258 VDPWR.n253 290.733
R4576 VDPWR.n101 VDPWR.n53 290.733
R4577 VDPWR.n77 VDPWR.n63 290.733
R4578 VDPWR.t249 VDPWR.t22 267.027
R4579 VDPWR.t347 VDPWR.t270 251.471
R4580 VDPWR.t131 VDPWR.t347 251.471
R4581 VDPWR.t28 VDPWR.t131 251.471
R4582 VDPWR.t32 VDPWR.t28 251.471
R4583 VDPWR.t415 VDPWR.t32 251.471
R4584 VDPWR.t239 VDPWR.t415 251.471
R4585 VDPWR.t26 VDPWR.t239 251.471
R4586 VDPWR.t30 VDPWR.t26 251.471
R4587 VDPWR.t228 VDPWR.t30 251.471
R4588 VDPWR.t121 VDPWR.t228 251.471
R4589 VDPWR.t349 VDPWR.t121 251.471
R4590 VDPWR.t86 VDPWR.t349 251.471
R4591 VDPWR.t226 VDPWR.t86 251.471
R4592 VDPWR.t119 VDPWR.t226 251.471
R4593 VDPWR.t44 VDPWR.t119 251.471
R4594 VDPWR.t212 VDPWR.t44 251.471
R4595 VDPWR.t264 VDPWR.t212 251.471
R4596 VDPWR.n393 VDPWR.n392 243.698
R4597 VDPWR.n363 VDPWR.n362 243.698
R4598 VDPWR.n339 VDPWR.n338 243.698
R4599 VDPWR.n315 VDPWR.n314 243.698
R4600 VDPWR.n298 VDPWR.n297 243.698
R4601 VDPWR.n386 VDPWR.n382 243.698
R4602 VDPWR.n356 VDPWR.n352 243.698
R4603 VDPWR.n346 VDPWR.n341 243.698
R4604 VDPWR.n322 VDPWR.n321 243.698
R4605 VDPWR.n306 VDPWR.n219 243.698
R4606 VDPWR.n524 VDPWR.n523 238.367
R4607 VDPWR.n524 VDPWR.n504 238.367
R4608 VDPWR.n534 VDPWR.n533 238.367
R4609 VDPWR.n534 VDPWR.n484 238.367
R4610 VDPWR.n591 VDPWR.n590 238.367
R4611 VDPWR.n611 VDPWR.n610 238.367
R4612 VDPWR.n611 VDPWR.n607 238.367
R4613 VDPWR.n647 VDPWR.n646 238.367
R4614 VDPWR.n647 VDPWR.n634 238.367
R4615 VDPWR.n657 VDPWR.n656 238.367
R4616 VDPWR.n657 VDPWR.n621 238.367
R4617 VDPWR.n381 VDPWR.n185 238.367
R4618 VDPWR.n379 VDPWR.n378 238.367
R4619 VDPWR.n372 VDPWR.n188 238.367
R4620 VDPWR.n351 VDPWR.n207 238.367
R4621 VDPWR.n334 VDPWR.n211 238.367
R4622 VDPWR.n318 VDPWR.n317 238.367
R4623 VDPWR.n301 VDPWR.n300 238.367
R4624 VDPWR.n396 VDPWR.n395 238.367
R4625 VDPWR.n204 VDPWR.n190 238.367
R4626 VDPWR.n366 VDPWR.n365 238.367
R4627 VDPWR.n349 VDPWR.n348 238.367
R4628 VDPWR.n327 VDPWR.n326 238.367
R4629 VDPWR.n309 VDPWR.n308 238.367
R4630 VDPWR.n197 VDPWR.n189 238.367
R4631 VDPWR.t270 VDPWR.n575 237.5
R4632 VDPWR.n592 VDPWR.t264 237.5
R4633 VDPWR.n172 VDPWR.t23 236.043
R4634 VDPWR.n474 VDPWR.n473 230.308
R4635 VDPWR.n477 VDPWR.n476 230.308
R4636 VDPWR.n444 VDPWR.n415 230.308
R4637 VDPWR.n292 VDPWR.n291 230.308
R4638 VDPWR.n286 VDPWR.n223 230.308
R4639 VDPWR.n273 VDPWR.n272 230.308
R4640 VDPWR.n267 VDPWR.n240 230.308
R4641 VDPWR.n235 VDPWR.n225 230.308
R4642 VDPWR.n282 VDPWR.n281 230.308
R4643 VDPWR.n279 VDPWR.n275 230.308
R4644 VDPWR.n252 VDPWR.n242 230.308
R4645 VDPWR.n247 VDPWR.n241 230.308
R4646 VDPWR.n230 VDPWR.n224 230.308
R4647 VDPWR.n105 VDPWR.n104 230.308
R4648 VDPWR.n108 VDPWR.n107 230.308
R4649 VDPWR.n98 VDPWR.n97 230.308
R4650 VDPWR.n88 VDPWR.n55 230.308
R4651 VDPWR.t200 VDPWR.t16 222.178
R4652 VDPWR.n174 VDPWR.n151 221.601
R4653 VDPWR.n299 VDPWR.n293 199.195
R4654 VDPWR.t198 VDPWR.t328 197.703
R4655 VDPWR.n427 VDPWR.n413 185.001
R4656 VDPWR.n456 VDPWR.n455 185.001
R4657 VDPWR.n463 VDPWR.n462 185.001
R4658 VDPWR.n467 VDPWR.n465 185
R4659 VDPWR.n470 VDPWR.n464 185
R4660 VDPWR.n475 VDPWR.n464 185
R4661 VDPWR.n469 VDPWR.n408 185
R4662 VDPWR.n453 VDPWR.n452 185
R4663 VDPWR.n454 VDPWR.n453 185
R4664 VDPWR.n418 VDPWR.n416 185
R4665 VDPWR.n449 VDPWR.n448 185
R4666 VDPWR.n447 VDPWR.n446 185
R4667 VDPWR.n580 VDPWR.n578 185
R4668 VDPWR.n587 VDPWR.n577 185
R4669 VDPWR.n592 VDPWR.n577 185
R4670 VDPWR.n586 VDPWR.n585 185
R4671 VDPWR.n583 VDPWR.n552 185
R4672 VDPWR.n594 VDPWR.n593 185
R4673 VDPWR.n593 VDPWR.n592 185
R4674 VDPWR.n574 VDPWR.n573 185
R4675 VDPWR.n575 VDPWR.n574 185
R4676 VDPWR.n571 VDPWR.n556 185
R4677 VDPWR.n570 VDPWR.n569 185
R4678 VDPWR.n568 VDPWR.n567 185
R4679 VDPWR.n562 VDPWR.n561 185
R4680 VDPWR.n564 VDPWR.n555 185
R4681 VDPWR.n575 VDPWR.n555 185
R4682 VDPWR.n251 VDPWR.n250 185
R4683 VDPWR.n249 VDPWR.n248 185
R4684 VDPWR.n239 VDPWR.n238 185
R4685 VDPWR.n278 VDPWR.n277 185
R4686 VDPWR.n234 VDPWR.n233 185
R4687 VDPWR.n232 VDPWR.n231 185
R4688 VDPWR.n303 VDPWR.n220 185
R4689 VDPWR.n305 VDPWR.n304 185
R4690 VDPWR.n325 VDPWR.n324 185
R4691 VDPWR.n323 VDPWR.n320 185
R4692 VDPWR.n343 VDPWR.n342 185
R4693 VDPWR.n345 VDPWR.n344 185
R4694 VDPWR.n353 VDPWR.n209 185
R4695 VDPWR.n355 VDPWR.n354 185
R4696 VDPWR.n199 VDPWR.n196 185
R4697 VDPWR.n201 VDPWR.n200 185
R4698 VDPWR.n383 VDPWR.n187 185
R4699 VDPWR.n385 VDPWR.n384 185
R4700 VDPWR.n271 VDPWR.n243 185
R4701 VDPWR.n269 VDPWR.n268 185
R4702 VDPWR.n290 VDPWR.n226 185
R4703 VDPWR.n288 VDPWR.n287 185
R4704 VDPWR.n296 VDPWR.n294 185
R4705 VDPWR.n295 VDPWR.n222 185
R4706 VDPWR.n313 VDPWR.n311 185
R4707 VDPWR.n312 VDPWR.n218 185
R4708 VDPWR.n213 VDPWR.n212 185
R4709 VDPWR.n336 VDPWR.n335 185
R4710 VDPWR.n358 VDPWR.n357 185
R4711 VDPWR.n360 VDPWR.n359 185
R4712 VDPWR.n193 VDPWR.n191 185
R4713 VDPWR.n375 VDPWR.n374 185
R4714 VDPWR.n388 VDPWR.n387 185
R4715 VDPWR.n390 VDPWR.n389 185
R4716 VDPWR.n264 VDPWR.n263 185
R4717 VDPWR.n263 VDPWR.n262 185
R4718 VDPWR.n255 VDPWR.n254 185
R4719 VDPWR.n259 VDPWR.n257 185
R4720 VDPWR.n261 VDPWR.n260 185
R4721 VDPWR.n262 VDPWR.n261 185
R4722 VDPWR.n175 VDPWR.n174 185
R4723 VDPWR.n60 VDPWR.n56 185
R4724 VDPWR.n86 VDPWR.n85 185
R4725 VDPWR.n102 VDPWR.n100 185
R4726 VDPWR.n54 VDPWR.n52 185
R4727 VDPWR.n76 VDPWR.n75 185
R4728 VDPWR.n75 VDPWR.n74 185
R4729 VDPWR.n67 VDPWR.n66 185
R4730 VDPWR.n72 VDPWR.n71 185
R4731 VDPWR.n73 VDPWR.n64 185
R4732 VDPWR.n74 VDPWR.n73 185
R4733 VDPWR.n262 VDPWR.t200 172.38
R4734 VDPWR.t190 VDPWR.n274 172.38
R4735 VDPWR.n280 VDPWR.t109 172.38
R4736 VDPWR.n97 VDPWR.n57 166.63
R4737 VDPWR.n176 VDPWR.n175 163.435
R4738 VDPWR.n173 VDPWR.n153 153.601
R4739 VDPWR.n180 VDPWR.n146 153.601
R4740 VDPWR.n50 VDPWR.n49 153.573
R4741 VDPWR.n92 VDPWR.n91 153.573
R4742 VDPWR.n94 VDPWR.n93 153.573
R4743 VDPWR.n83 VDPWR.n82 153.573
R4744 VDPWR.n81 VDPWR.n80 153.573
R4745 VDPWR.n79 VDPWR.n78 153.573
R4746 VDPWR.n578 VDPWR.n577 150
R4747 VDPWR.n585 VDPWR.n577 150
R4748 VDPWR.n593 VDPWR.n552 150
R4749 VDPWR.n574 VDPWR.n556 150
R4750 VDPWR.n569 VDPWR.n568 150
R4751 VDPWR.n561 VDPWR.n555 150
R4752 VDPWR.n389 VDPWR.n387 150
R4753 VDPWR.n374 VDPWR.n191 150
R4754 VDPWR.n359 VDPWR.n357 150
R4755 VDPWR.n335 VDPWR.n212 150
R4756 VDPWR.n311 VDPWR.n218 150
R4757 VDPWR.n294 VDPWR.n222 150
R4758 VDPWR.n385 VDPWR.n187 150
R4759 VDPWR.n200 VDPWR.n199 150
R4760 VDPWR.n355 VDPWR.n209 150
R4761 VDPWR.n344 VDPWR.n342 150
R4762 VDPWR.n325 VDPWR.n320 150
R4763 VDPWR.n304 VDPWR.n220 150
R4764 VDPWR.t93 VDPWR.t97 145.038
R4765 VDPWR.n153 VDPWR.n152 144
R4766 VDPWR.n596 VDPWR.n549 141.712
R4767 VDPWR.n597 VDPWR.n548 141.712
R4768 VDPWR.n598 VDPWR.n547 141.712
R4769 VDPWR.n599 VDPWR.n546 141.712
R4770 VDPWR.n600 VDPWR.n545 141.712
R4771 VDPWR.n601 VDPWR.n544 141.712
R4772 VDPWR.n602 VDPWR.n543 141.712
R4773 VDPWR.n603 VDPWR.n542 141.712
R4774 VDPWR.n316 VDPWR.n310 137.904
R4775 VDPWR.n340 VDPWR.n210 137.904
R4776 VDPWR.n178 VDPWR.t330 126.865
R4777 VDPWR.n262 VDPWR.t230 126.412
R4778 VDPWR.n274 VDPWR.t16 126.412
R4779 VDPWR.n280 VDPWR.t190 126.412
R4780 VDPWR.n293 VDPWR.t109 126.412
R4781 VDPWR.n405 VDPWR.n404 123.987
R4782 VDPWR.n432 VDPWR.n431 123.987
R4783 VDPWR.n434 VDPWR.n433 123.987
R4784 VDPWR.n440 VDPWR.n439 123.987
R4785 VDPWR.t234 VDPWR.n177 123.243
R4786 VDPWR.t271 VDPWR.n559 123.126
R4787 VDPWR.n560 VDPWR.t271 123.126
R4788 VDPWR.n588 VDPWR.t265 123.126
R4789 VDPWR.n584 VDPWR.t265 123.126
R4790 VDPWR.t324 VDPWR.n195 123.126
R4791 VDPWR.n198 VDPWR.t324 123.126
R4792 VDPWR.t152 VDPWR.n192 123.126
R4793 VDPWR.n373 VDPWR.t152 123.126
R4794 VDPWR.n465 VDPWR.n464 120.001
R4795 VDPWR.n464 VDPWR.n408 120.001
R4796 VDPWR.n453 VDPWR.n416 120.001
R4797 VDPWR.n448 VDPWR.n447 120.001
R4798 VDPWR.n287 VDPWR.n226 120.001
R4799 VDPWR.n268 VDPWR.n243 120.001
R4800 VDPWR.n233 VDPWR.n232 120.001
R4801 VDPWR.n278 VDPWR.n239 120.001
R4802 VDPWR.n250 VDPWR.n249 120.001
R4803 VDPWR.n263 VDPWR.n255 120.001
R4804 VDPWR.n261 VDPWR.n257 120.001
R4805 VDPWR.n100 VDPWR.n54 120.001
R4806 VDPWR.n85 VDPWR.n56 120.001
R4807 VDPWR.n75 VDPWR.n67 120.001
R4808 VDPWR.n73 VDPWR.n72 120.001
R4809 VDPWR.t283 VDPWR.n413 119.656
R4810 VDPWR.n436 VDPWR.n435 119.424
R4811 VDPWR.n455 VDPWR.n454 108.779
R4812 VDPWR.t22 VDPWR.n176 107.507
R4813 VDPWR.n364 VDPWR.n350 107.258
R4814 VDPWR.n364 VDPWR.t34 103.427
R4815 VDPWR.n380 VDPWR.t377 103.427
R4816 VDPWR.t151 VDPWR.n380 103.427
R4817 VDPWR.n394 VDPWR.t69 103.427
R4818 VDPWR.n350 VDPWR.t129 95.7666
R4819 VDPWR.t273 VDPWR.t49 94.2753
R4820 VDPWR.t49 VDPWR.t6 94.2753
R4821 VDPWR.t6 VDPWR.t159 94.2753
R4822 VDPWR.t159 VDPWR.t390 94.2753
R4823 VDPWR.t390 VDPWR.t283 94.2753
R4824 VDPWR.t67 VDPWR.t386 94.2753
R4825 VDPWR.t218 VDPWR.t307 94.2753
R4826 VDPWR.n463 VDPWR.t99 94.2753
R4827 VDPWR.t248 VDPWR.t82 94.2753
R4828 VDPWR.t333 VDPWR.t332 94.2753
R4829 VDPWR.n152 VDPWR.n148 92.5005
R4830 VDPWR.n177 VDPWR.n148 92.5005
R4831 VDPWR.n149 VDPWR.n147 92.5005
R4832 VDPWR.n177 VDPWR.n149 92.5005
R4833 VDPWR.t246 VDPWR.t388 91.936
R4834 VDPWR.t24 VDPWR.t115 91.936
R4835 VDPWR.n176 VDPWR.n150 84.8581
R4836 VDPWR.t334 VDPWR.t405 84.2747
R4837 VDPWR.t34 VDPWR.t2 84.2747
R4838 VDPWR.t175 VDPWR.t377 84.2747
R4839 VDPWR.t379 VDPWR.t151 84.2747
R4840 VDPWR.t69 VDPWR.t55 84.2747
R4841 VDPWR.t258 VDPWR.t267 83.3974
R4842 VDPWR.t5 VDPWR.t105 83.3974
R4843 VDPWR.n459 VDPWR.n458 83.2005
R4844 VDPWR.n460 VDPWR.n459 83.2005
R4845 VDPWR.n430 VDPWR.n425 83.2005
R4846 VDPWR.n430 VDPWR.n429 83.2005
R4847 VDPWR.n0 VDPWR.t154 78.8005
R4848 VDPWR.n0 VDPWR.t370 78.8005
R4849 VDPWR.n39 VDPWR.t15 78.8005
R4850 VDPWR.n39 VDPWR.t90 78.8005
R4851 VDPWR.n41 VDPWR.t75 78.8005
R4852 VDPWR.n41 VDPWR.t150 78.8005
R4853 VDPWR.n37 VDPWR.t408 78.8005
R4854 VDPWR.n37 VDPWR.t368 78.8005
R4855 VDPWR.n35 VDPWR.t183 78.8005
R4856 VDPWR.n35 VDPWR.t62 78.8005
R4857 VDPWR.n31 VDPWR.t37 78.8005
R4858 VDPWR.n31 VDPWR.t352 78.8005
R4859 VDPWR.n29 VDPWR.t385 78.8005
R4860 VDPWR.n29 VDPWR.t170 78.8005
R4861 VDPWR.n2 VDPWR.t73 78.8005
R4862 VDPWR.n2 VDPWR.t217 78.8005
R4863 VDPWR.n21 VDPWR.t372 78.8005
R4864 VDPWR.n21 VDPWR.t210 78.8005
R4865 VDPWR.n19 VDPWR.t158 78.8005
R4866 VDPWR.n19 VDPWR.t64 78.8005
R4867 VDPWR.n17 VDPWR.t338 78.8005
R4868 VDPWR.n17 VDPWR.t66 78.8005
R4869 VDPWR.n4 VDPWR.t202 78.8005
R4870 VDPWR.n4 VDPWR.t81 78.8005
R4871 VDPWR.n9 VDPWR.t243 78.8005
R4872 VDPWR.n9 VDPWR.t323 78.8005
R4873 VDPWR.n7 VDPWR.t1 78.8005
R4874 VDPWR.n7 VDPWR.t381 78.8005
R4875 VDPWR.n6 VDPWR.t177 78.8005
R4876 VDPWR.n6 VDPWR.t114 78.8005
R4877 VDPWR.t91 VDPWR.t232 76.1455
R4878 VDPWR.t83 VDPWR.t303 76.1455
R4879 VDPWR.n177 VDPWR.t238 74.46
R4880 VDPWR.n265 VDPWR.n264 72.1074
R4881 VDPWR.n348 VDPWR.n206 71.8576
R4882 VDPWR.n283 VDPWR.n282 71.0449
R4883 VDPWR.n475 VDPWR.n474 69.8479
R4884 VDPWR.n476 VDPWR.n475 69.8479
R4885 VDPWR.n454 VDPWR.n414 69.8479
R4886 VDPWR.n454 VDPWR.n415 69.8479
R4887 VDPWR.n274 VDPWR.n242 69.8479
R4888 VDPWR.n274 VDPWR.n241 69.8479
R4889 VDPWR.n281 VDPWR.n280 69.8479
R4890 VDPWR.n280 VDPWR.n279 69.8479
R4891 VDPWR.n293 VDPWR.n225 69.8479
R4892 VDPWR.n293 VDPWR.n224 69.8479
R4893 VDPWR.n274 VDPWR.n273 69.8479
R4894 VDPWR.n274 VDPWR.n240 69.8479
R4895 VDPWR.n293 VDPWR.n292 69.8479
R4896 VDPWR.n293 VDPWR.n223 69.8479
R4897 VDPWR.n262 VDPWR.n256 69.8479
R4898 VDPWR.n99 VDPWR.n98 69.8479
R4899 VDPWR.n99 VDPWR.n55 69.8479
R4900 VDPWR.n106 VDPWR.n105 69.8479
R4901 VDPWR.n107 VDPWR.n106 69.8479
R4902 VDPWR.n74 VDPWR.n68 69.8479
R4903 VDPWR.t238 VDPWR.t249 69.3248
R4904 VDPWR.t328 VDPWR.t234 69.3248
R4905 VDPWR.t330 VDPWR.t198 69.3248
R4906 VDPWR.t232 VDPWR.t103 68.8936
R4907 VDPWR.n475 VDPWR.t83 68.8936
R4908 VDPWR.n48 VDPWR.n47 68.2005
R4909 VDPWR.n44 VDPWR.n43 68.2005
R4910 VDPWR.n28 VDPWR.n27 68.2005
R4911 VDPWR.n24 VDPWR.n23 68.2005
R4912 VDPWR.n16 VDPWR.n15 68.2005
R4913 VDPWR.n12 VDPWR.n11 68.2005
R4914 VDPWR.n592 VDPWR.n591 65.8183
R4915 VDPWR.n592 VDPWR.n576 65.8183
R4916 VDPWR.n575 VDPWR.n553 65.8183
R4917 VDPWR.n575 VDPWR.n554 65.8183
R4918 VDPWR.n310 VDPWR.n309 65.8183
R4919 VDPWR.n310 VDPWR.n219 65.8183
R4920 VDPWR.n326 VDPWR.n210 65.8183
R4921 VDPWR.n321 VDPWR.n210 65.8183
R4922 VDPWR.n350 VDPWR.n349 65.8183
R4923 VDPWR.n350 VDPWR.n341 65.8183
R4924 VDPWR.n365 VDPWR.n364 65.8183
R4925 VDPWR.n364 VDPWR.n356 65.8183
R4926 VDPWR.n380 VDPWR.n190 65.8183
R4927 VDPWR.n380 VDPWR.n189 65.8183
R4928 VDPWR.n395 VDPWR.n394 65.8183
R4929 VDPWR.n394 VDPWR.n386 65.8183
R4930 VDPWR.n299 VDPWR.n298 65.8183
R4931 VDPWR.n300 VDPWR.n299 65.8183
R4932 VDPWR.n316 VDPWR.n315 65.8183
R4933 VDPWR.n317 VDPWR.n316 65.8183
R4934 VDPWR.n340 VDPWR.n339 65.8183
R4935 VDPWR.n340 VDPWR.n211 65.8183
R4936 VDPWR.n364 VDPWR.n363 65.8183
R4937 VDPWR.n364 VDPWR.n351 65.8183
R4938 VDPWR.n380 VDPWR.n379 65.8183
R4939 VDPWR.n380 VDPWR.n188 65.8183
R4940 VDPWR.n394 VDPWR.n393 65.8183
R4941 VDPWR.n394 VDPWR.n381 65.8183
R4942 VDPWR.t267 VDPWR.t95 61.6417
R4943 VDPWR.t101 VDPWR.t5 61.6417
R4944 VDPWR.n401 VDPWR.t423 58.8005
R4945 VDPWR.n400 VDPWR.t424 58.8005
R4946 VDPWR.n397 VDPWR.n185 58.0576
R4947 VDPWR.n397 VDPWR.n396 58.0576
R4948 VDPWR.n367 VDPWR.n207 58.0576
R4949 VDPWR.n367 VDPWR.n366 58.0576
R4950 VDPWR.n328 VDPWR.n318 58.0576
R4951 VDPWR.n328 VDPWR.n327 58.0576
R4952 VDPWR.n302 VDPWR.n301 58.0576
R4953 VDPWR.n308 VDPWR.n302 58.0576
R4954 VDPWR.n286 VDPWR.n285 57.2449
R4955 VDPWR.n285 VDPWR.n235 57.2449
R4956 VDPWR.n267 VDPWR.n266 57.2449
R4957 VDPWR.n266 VDPWR.n252 57.2449
R4958 VDPWR.n441 VDPWR.n430 56.338
R4959 VDPWR.n334 VDPWR.n333 54.8576
R4960 VDPWR.n371 VDPWR.n194 54.4005
R4961 VDPWR.n205 VDPWR.n194 54.4005
R4962 VDPWR.n371 VDPWR.n370 54.4005
R4963 VDPWR.n370 VDPWR.n205 54.4005
R4964 VDPWR.n585 VDPWR.n576 53.3664
R4965 VDPWR.n591 VDPWR.n578 53.3664
R4966 VDPWR.n576 VDPWR.n552 53.3664
R4967 VDPWR.n556 VDPWR.n553 53.3664
R4968 VDPWR.n568 VDPWR.n554 53.3664
R4969 VDPWR.n569 VDPWR.n553 53.3664
R4970 VDPWR.n561 VDPWR.n554 53.3664
R4971 VDPWR.n386 VDPWR.n385 53.3664
R4972 VDPWR.n200 VDPWR.n189 53.3664
R4973 VDPWR.n356 VDPWR.n355 53.3664
R4974 VDPWR.n309 VDPWR.n220 53.3664
R4975 VDPWR.n304 VDPWR.n219 53.3664
R4976 VDPWR.n326 VDPWR.n325 53.3664
R4977 VDPWR.n321 VDPWR.n320 53.3664
R4978 VDPWR.n349 VDPWR.n342 53.3664
R4979 VDPWR.n344 VDPWR.n341 53.3664
R4980 VDPWR.n365 VDPWR.n209 53.3664
R4981 VDPWR.n199 VDPWR.n190 53.3664
R4982 VDPWR.n395 VDPWR.n187 53.3664
R4983 VDPWR.n298 VDPWR.n294 53.3664
R4984 VDPWR.n300 VDPWR.n222 53.3664
R4985 VDPWR.n315 VDPWR.n311 53.3664
R4986 VDPWR.n317 VDPWR.n218 53.3664
R4987 VDPWR.n339 VDPWR.n212 53.3664
R4988 VDPWR.n335 VDPWR.n211 53.3664
R4989 VDPWR.n363 VDPWR.n357 53.3664
R4990 VDPWR.n359 VDPWR.n351 53.3664
R4991 VDPWR.n379 VDPWR.n191 53.3664
R4992 VDPWR.n374 VDPWR.n188 53.3664
R4993 VDPWR.n393 VDPWR.n387 53.3664
R4994 VDPWR.n389 VDPWR.n381 53.3664
R4995 VDPWR.n459 VDPWR.n410 50.9005
R4996 VDPWR.t97 VDPWR.n463 50.7639
R4997 VDPWR.n411 VDPWR.t387 49.2505
R4998 VDPWR.n411 VDPWR.t233 49.2505
R4999 VDPWR.n409 VDPWR.t219 49.2505
R5000 VDPWR.n409 VDPWR.t308 49.2505
R5001 VDPWR.t268 VDPWR.n412 49.2505
R5002 VDPWR.n412 VDPWR.t68 49.2505
R5003 VDPWR.n421 VDPWR.t7 49.2505
R5004 VDPWR.n421 VDPWR.t160 49.2505
R5005 VDPWR.n426 VDPWR.t391 49.2505
R5006 VDPWR.n426 VDPWR.t284 49.2505
R5007 VDPWR.t274 VDPWR.n422 49.2505
R5008 VDPWR.n422 VDPWR.t50 49.2505
R5009 VDPWR.n400 VDPWR.t425 49.1638
R5010 VDPWR.n402 VDPWR.t429 48.5162
R5011 VDPWR.n476 VDPWR.n408 45.3071
R5012 VDPWR.n474 VDPWR.n465 45.3071
R5013 VDPWR.n416 VDPWR.n414 45.3071
R5014 VDPWR.n447 VDPWR.n415 45.3071
R5015 VDPWR.n448 VDPWR.n414 45.3071
R5016 VDPWR.n232 VDPWR.n224 45.3071
R5017 VDPWR.n249 VDPWR.n241 45.3071
R5018 VDPWR.n250 VDPWR.n242 45.3071
R5019 VDPWR.n281 VDPWR.n239 45.3071
R5020 VDPWR.n279 VDPWR.n278 45.3071
R5021 VDPWR.n233 VDPWR.n225 45.3071
R5022 VDPWR.n273 VDPWR.n243 45.3071
R5023 VDPWR.n268 VDPWR.n240 45.3071
R5024 VDPWR.n292 VDPWR.n226 45.3071
R5025 VDPWR.n287 VDPWR.n223 45.3071
R5026 VDPWR.n256 VDPWR.n255 45.3071
R5027 VDPWR.n257 VDPWR.n256 45.3071
R5028 VDPWR.n98 VDPWR.n56 45.3071
R5029 VDPWR.n85 VDPWR.n55 45.3071
R5030 VDPWR.n105 VDPWR.n100 45.3071
R5031 VDPWR.n107 VDPWR.n54 45.3071
R5032 VDPWR.n68 VDPWR.n67 45.3071
R5033 VDPWR.n72 VDPWR.n68 45.3071
R5034 VDPWR.t82 VDPWR.t93 39.886
R5035 VDPWR.n519 VDPWR.t60 39.4005
R5036 VDPWR.n519 VDPWR.t181 39.4005
R5037 VDPWR.n517 VDPWR.t206 39.4005
R5038 VDPWR.n517 VDPWR.t128 39.4005
R5039 VDPWR.n515 VDPWR.t221 39.4005
R5040 VDPWR.n515 VDPWR.t13 39.4005
R5041 VDPWR.n513 VDPWR.t148 39.4005
R5042 VDPWR.n513 VDPWR.t344 39.4005
R5043 VDPWR.n511 VDPWR.t77 39.4005
R5044 VDPWR.n511 VDPWR.t179 39.4005
R5045 VDPWR.n509 VDPWR.t326 39.4005
R5046 VDPWR.n509 VDPWR.t358 39.4005
R5047 VDPWR.n507 VDPWR.t193 39.4005
R5048 VDPWR.n507 VDPWR.t11 39.4005
R5049 VDPWR.n505 VDPWR.t21 39.4005
R5050 VDPWR.n505 VDPWR.t404 39.4005
R5051 VDPWR.n501 VDPWR.t346 39.4005
R5052 VDPWR.n501 VDPWR.t197 39.4005
R5053 VDPWR.n499 VDPWR.t58 39.4005
R5054 VDPWR.n499 VDPWR.t422 39.4005
R5055 VDPWR.n497 VDPWR.t146 39.4005
R5056 VDPWR.n497 VDPWR.t237 39.4005
R5057 VDPWR.n495 VDPWR.t85 39.4005
R5058 VDPWR.n495 VDPWR.t4 39.4005
R5059 VDPWR.n493 VDPWR.t376 39.4005
R5060 VDPWR.n493 VDPWR.t185 39.4005
R5061 VDPWR.n491 VDPWR.t19 39.4005
R5062 VDPWR.n491 VDPWR.t112 39.4005
R5063 VDPWR.n489 VDPWR.t43 39.4005
R5064 VDPWR.n489 VDPWR.t189 39.4005
R5065 VDPWR.n487 VDPWR.t195 39.4005
R5066 VDPWR.n487 VDPWR.t187 39.4005
R5067 VDPWR.n485 VDPWR.t204 39.4005
R5068 VDPWR.n485 VDPWR.t413 39.4005
R5069 VDPWR.n481 VDPWR.t9 39.4005
R5070 VDPWR.n481 VDPWR.t402 39.4005
R5071 VDPWR.n642 VDPWR.t142 39.4005
R5072 VDPWR.n642 VDPWR.t420 39.4005
R5073 VDPWR.n640 VDPWR.t135 39.4005
R5074 VDPWR.n640 VDPWR.t223 39.4005
R5075 VDPWR.n638 VDPWR.t172 39.4005
R5076 VDPWR.n638 VDPWR.t39 39.4005
R5077 VDPWR.n636 VDPWR.t225 39.4005
R5078 VDPWR.n636 VDPWR.t164 39.4005
R5079 VDPWR.n631 VDPWR.t52 39.4005
R5080 VDPWR.n631 VDPWR.t366 39.4005
R5081 VDPWR.n629 VDPWR.t166 39.4005
R5082 VDPWR.n629 VDPWR.t356 39.4005
R5083 VDPWR.n627 VDPWR.t137 39.4005
R5084 VDPWR.n627 VDPWR.t418 39.4005
R5085 VDPWR.n625 VDPWR.t174 39.4005
R5086 VDPWR.n625 VDPWR.t41 39.4005
R5087 VDPWR.n623 VDPWR.t354 39.4005
R5088 VDPWR.n623 VDPWR.t364 39.4005
R5089 VDPWR.n618 VDPWR.t54 39.4005
R5090 VDPWR.n618 VDPWR.t144 39.4005
R5091 VDPWR.n179 VDPWR.n178 37.0005
R5092 VDPWR.n151 VDPWR.n150 37.0005
R5093 VDPWR.n455 VDPWR.t258 36.26
R5094 VDPWR.t95 VDPWR.t67 32.6341
R5095 VDPWR.t332 VDPWR.t101 32.6341
R5096 VDPWR.n428 VDPWR.n427 30.754
R5097 VDPWR.n424 VDPWR.n423 30.186
R5098 VDPWR.n462 VDPWR.n461 30.18
R5099 VDPWR.n457 VDPWR.n456 29.7151
R5100 VDPWR.t103 VDPWR.t218 25.3822
R5101 VDPWR.t307 VDPWR.t99 25.3822
R5102 VDPWR.n228 VDPWR.t110 24.6255
R5103 VDPWR.n227 VDPWR.t336 24.6255
R5104 VDPWR.n237 VDPWR.t191 24.6255
R5105 VDPWR.n245 VDPWR.t56 24.6255
R5106 VDPWR.n244 VDPWR.t17 24.6255
R5107 VDPWR.n253 VDPWR.t231 24.6255
R5108 VDPWR.n49 VDPWR.t124 24.6255
R5109 VDPWR.n49 VDPWR.t291 24.6255
R5110 VDPWR.n91 VDPWR.t340 24.6255
R5111 VDPWR.n91 VDPWR.t342 24.6255
R5112 VDPWR.t312 VDPWR.n94 24.6255
R5113 VDPWR.n94 VDPWR.t383 24.6255
R5114 VDPWR.n82 VDPWR.t362 24.6255
R5115 VDPWR.n82 VDPWR.t280 24.6255
R5116 VDPWR.n80 VDPWR.t139 24.6255
R5117 VDPWR.n80 VDPWR.t156 24.6255
R5118 VDPWR.n78 VDPWR.t315 24.6255
R5119 VDPWR.n78 VDPWR.t118 24.6255
R5120 VDPWR.t315 VDPWR.n77 24.6255
R5121 VDPWR.n53 VDPWR.t292 24.6255
R5122 VDPWR.n95 VDPWR.t312 24.6255
R5123 VDPWR.n59 VDPWR.t281 24.6255
R5124 VDPWR.n595 VDPWR.n594 22.8576
R5125 VDPWR.n564 VDPWR.n541 22.8576
R5126 VDPWR.n128 VDPWR.n127 21.6365
R5127 VDPWR.n126 VDPWR.n123 21.6365
R5128 VDPWR.n122 VDPWR.n121 21.6365
R5129 VDPWR.n120 VDPWR.n117 21.6365
R5130 VDPWR.n144 VDPWR.n143 21.6365
R5131 VDPWR.n142 VDPWR.n139 21.6365
R5132 VDPWR.n138 VDPWR.n137 21.6365
R5133 VDPWR.n136 VDPWR.n133 21.6365
R5134 VDPWR.n169 VDPWR.n168 21.6365
R5135 VDPWR.n167 VDPWR.n164 21.6365
R5136 VDPWR.n163 VDPWR.n162 21.6365
R5137 VDPWR.n161 VDPWR.n158 21.6365
R5138 VDPWR.n125 VDPWR.n114 21.3338
R5139 VDPWR.n119 VDPWR.n116 21.3338
R5140 VDPWR.n141 VDPWR.n130 21.3338
R5141 VDPWR.n135 VDPWR.n132 21.3338
R5142 VDPWR.n166 VDPWR.n155 21.3338
R5143 VDPWR.n160 VDPWR.n157 21.3338
R5144 VDPWR.n435 VDPWR.t92 19.7005
R5145 VDPWR.n435 VDPWR.t104 19.7005
R5146 VDPWR.n404 VDPWR.t102 19.7005
R5147 VDPWR.n404 VDPWR.t304 19.7005
R5148 VDPWR.n431 VDPWR.t94 19.7005
R5149 VDPWR.n431 VDPWR.t106 19.7005
R5150 VDPWR.n433 VDPWR.t100 19.7005
R5151 VDPWR.n433 VDPWR.t98 19.7005
R5152 VDPWR.n439 VDPWR.t259 19.7005
R5153 VDPWR.n439 VDPWR.t96 19.7005
R5154 VDPWR.t259 VDPWR.n417 19.7005
R5155 VDPWR.n472 VDPWR.t305 19.7005
R5156 VDPWR.n403 VDPWR.t133 18.3076
R5157 VDPWR.t386 VDPWR.t91 18.1303
R5158 VDPWR.t303 VDPWR.t333 18.1303
R5159 VDPWR.n461 VDPWR.n460 16.0005
R5160 VDPWR.n458 VDPWR.n457 16.0005
R5161 VDPWR.n429 VDPWR.n428 16.0005
R5162 VDPWR.n425 VDPWR.n424 16.0005
R5163 VDPWR.n478 VDPWR.n477 15.6449
R5164 VDPWR.n479 VDPWR.n478 14.0505
R5165 VDPWR.n266 VDPWR.n265 13.8005
R5166 VDPWR.n285 VDPWR.n284 13.8005
R5167 VDPWR.n302 VDPWR.n216 13.8005
R5168 VDPWR.n329 VDPWR.n328 13.8005
R5169 VDPWR.n368 VDPWR.n367 13.8005
R5170 VDPWR.n370 VDPWR.n369 13.8005
R5171 VDPWR.n194 VDPWR.n184 13.8005
R5172 VDPWR.n398 VDPWR.n397 13.8005
R5173 VDPWR.n549 VDPWR.t45 13.1338
R5174 VDPWR.n549 VDPWR.t213 13.1338
R5175 VDPWR.n548 VDPWR.t227 13.1338
R5176 VDPWR.n548 VDPWR.t120 13.1338
R5177 VDPWR.n547 VDPWR.t350 13.1338
R5178 VDPWR.n547 VDPWR.t87 13.1338
R5179 VDPWR.n546 VDPWR.t229 13.1338
R5180 VDPWR.n546 VDPWR.t122 13.1338
R5181 VDPWR.n545 VDPWR.t27 13.1338
R5182 VDPWR.n545 VDPWR.t31 13.1338
R5183 VDPWR.n544 VDPWR.t416 13.1338
R5184 VDPWR.n544 VDPWR.t240 13.1338
R5185 VDPWR.n543 VDPWR.t29 13.1338
R5186 VDPWR.n543 VDPWR.t33 13.1338
R5187 VDPWR.n542 VDPWR.t348 13.1338
R5188 VDPWR.n542 VDPWR.t132 13.1338
R5189 VDPWR.n333 VDPWR.n214 12.8005
R5190 VDPWR.n299 VDPWR.t246 11.4924
R5191 VDPWR.n310 VDPWR.t388 11.4924
R5192 VDPWR.n316 VDPWR.t24 11.4924
R5193 VDPWR.t115 VDPWR.n210 11.4924
R5194 VDPWR.t405 VDPWR.n340 11.4924
R5195 VDPWR.n596 VDPWR.n595 11.0575
R5196 VDPWR.t105 VDPWR.t248 10.8784
R5197 VDPWR.n604 VDPWR.n541 10.87
R5198 VDPWR.n123 VDPWR.n122 10.1932
R5199 VDPWR.n139 VDPWR.n138 10.1932
R5200 VDPWR.n164 VDPWR.n163 10.1932
R5201 VDPWR.n152 VDPWR.n146 9.6005
R5202 VDPWR.n527 VDPWR.n503 9.50883
R5203 VDPWR.n537 VDPWR.n483 9.50883
R5204 VDPWR.n573 VDPWR.n572 9.50883
R5205 VDPWR.n565 VDPWR.n564 9.50883
R5206 VDPWR.n590 VDPWR.n579 9.50883
R5207 VDPWR.n594 VDPWR.n551 9.50883
R5208 VDPWR.n614 VDPWR.n606 9.50883
R5209 VDPWR.n477 VDPWR.n406 9.45675
R5210 VDPWR.n469 VDPWR.n406 9.3005
R5211 VDPWR.n470 VDPWR.n468 9.3005
R5212 VDPWR.n446 VDPWR.n419 9.3005
R5213 VDPWR.n450 VDPWR.n449 9.3005
R5214 VDPWR.n444 VDPWR.n443 9.3005
R5215 VDPWR.n527 VDPWR.n526 9.3005
R5216 VDPWR.n537 VDPWR.n536 9.3005
R5217 VDPWR.n583 VDPWR.n551 9.3005
R5218 VDPWR.n586 VDPWR.n582 9.3005
R5219 VDPWR.n587 VDPWR.n581 9.3005
R5220 VDPWR.n580 VDPWR.n579 9.3005
R5221 VDPWR.n565 VDPWR.n562 9.3005
R5222 VDPWR.n567 VDPWR.n566 9.3005
R5223 VDPWR.n570 VDPWR.n558 9.3005
R5224 VDPWR.n572 VDPWR.n571 9.3005
R5225 VDPWR.n614 VDPWR.n613 9.3005
R5226 VDPWR.n333 VDPWR.n332 9.3005
R5227 VDPWR.n215 VDPWR.n214 9.3005
R5228 VDPWR.n119 VDPWR.n118 9.3005
R5229 VDPWR.n116 VDPWR.n115 9.3005
R5230 VDPWR.n125 VDPWR.n124 9.3005
R5231 VDPWR.n114 VDPWR.n113 9.3005
R5232 VDPWR.n135 VDPWR.n134 9.3005
R5233 VDPWR.n132 VDPWR.n131 9.3005
R5234 VDPWR.n141 VDPWR.n140 9.3005
R5235 VDPWR.n130 VDPWR.n129 9.3005
R5236 VDPWR.n160 VDPWR.n159 9.3005
R5237 VDPWR.n157 VDPWR.n156 9.3005
R5238 VDPWR.n166 VDPWR.n165 9.3005
R5239 VDPWR.n155 VDPWR.n154 9.3005
R5240 VDPWR.n170 VDPWR.n153 9.3005
R5241 VDPWR.n146 VDPWR.n145 9.3005
R5242 VDPWR.n181 VDPWR.n180 9.3005
R5243 VDPWR.n173 VDPWR.n172 9.3005
R5244 VDPWR.n52 VDPWR.n51 9.3005
R5245 VDPWR.n109 VDPWR.n108 9.3005
R5246 VDPWR.n71 VDPWR.n70 9.3005
R5247 VDPWR.n69 VDPWR.n64 9.3005
R5248 VDPWR.n587 VDPWR.n580 9.14336
R5249 VDPWR.n587 VDPWR.n586 9.14336
R5250 VDPWR.n586 VDPWR.n583 9.14336
R5251 VDPWR.n571 VDPWR.n570 9.14336
R5252 VDPWR.n570 VDPWR.n567 9.14336
R5253 VDPWR.n567 VDPWR.n562 9.14336
R5254 VDPWR.n336 VDPWR.n213 9.14336
R5255 VDPWR.n390 VDPWR.n388 9.14336
R5256 VDPWR.n384 VDPWR.n383 9.14336
R5257 VDPWR.n360 VDPWR.n358 9.14336
R5258 VDPWR.n354 VDPWR.n353 9.14336
R5259 VDPWR.n345 VDPWR.n343 9.14336
R5260 VDPWR.n313 VDPWR.n312 9.14336
R5261 VDPWR.n324 VDPWR.n323 9.14336
R5262 VDPWR.n296 VDPWR.n295 9.14336
R5263 VDPWR.n305 VDPWR.n303 9.14336
R5264 VDPWR.n127 VDPWR.n114 8.68224
R5265 VDPWR.n126 VDPWR.n125 8.68224
R5266 VDPWR.n121 VDPWR.n116 8.68224
R5267 VDPWR.n120 VDPWR.n119 8.68224
R5268 VDPWR.n143 VDPWR.n130 8.68224
R5269 VDPWR.n142 VDPWR.n141 8.68224
R5270 VDPWR.n137 VDPWR.n132 8.68224
R5271 VDPWR.n136 VDPWR.n135 8.68224
R5272 VDPWR.n168 VDPWR.n155 8.68224
R5273 VDPWR.n167 VDPWR.n166 8.68224
R5274 VDPWR.n162 VDPWR.n157 8.68224
R5275 VDPWR.n161 VDPWR.n160 8.68224
R5276 VDPWR.t129 VDPWR.t334 7.66179
R5277 VDPWR.n454 VDPWR.n413 7.25241
R5278 VDPWR.n470 VDPWR.n469 7.11161
R5279 VDPWR.n449 VDPWR.n446 7.11161
R5280 VDPWR.n291 VDPWR.n290 7.11161
R5281 VDPWR.n288 VDPWR.n286 7.11161
R5282 VDPWR.n235 VDPWR.n234 7.11161
R5283 VDPWR.n231 VDPWR.n230 7.11161
R5284 VDPWR.n282 VDPWR.n238 7.11161
R5285 VDPWR.n277 VDPWR.n275 7.11161
R5286 VDPWR.n272 VDPWR.n271 7.11161
R5287 VDPWR.n269 VDPWR.n267 7.11161
R5288 VDPWR.n252 VDPWR.n251 7.11161
R5289 VDPWR.n248 VDPWR.n247 7.11161
R5290 VDPWR.n264 VDPWR.n254 7.11161
R5291 VDPWR.n260 VDPWR.n259 7.11161
R5292 VDPWR.n108 VDPWR.n52 7.11161
R5293 VDPWR.n71 VDPWR.n64 7.11161
R5294 VDPWR.n375 VDPWR.n193 5.81868
R5295 VDPWR.n201 VDPWR.n196 5.81868
R5296 VDPWR.n172 VDPWR.n171 5.46925
R5297 VDPWR.n663 VDPWR.n662 5.34031
R5298 VDPWR.n590 VDPWR.n589 5.33286
R5299 VDPWR.n594 VDPWR.n550 5.33286
R5300 VDPWR.n573 VDPWR.n557 5.33286
R5301 VDPWR.n564 VDPWR.n563 5.33286
R5302 VDPWR.n337 VDPWR.n334 5.33286
R5303 VDPWR.n391 VDPWR.n185 5.33286
R5304 VDPWR.n396 VDPWR.n186 5.33286
R5305 VDPWR.n361 VDPWR.n207 5.33286
R5306 VDPWR.n366 VDPWR.n208 5.33286
R5307 VDPWR.n348 VDPWR.n347 5.33286
R5308 VDPWR.n318 VDPWR.n217 5.33286
R5309 VDPWR.n327 VDPWR.n319 5.33286
R5310 VDPWR.n301 VDPWR.n221 5.33286
R5311 VDPWR.n308 VDPWR.n307 5.33286
R5312 VDPWR.n79 VDPWR.n62 5.01612
R5313 VDPWR.n644 VDPWR.n643 4.84425
R5314 VDPWR.n666 VDPWR.n48 4.8216
R5315 VDPWR.n90 VDPWR.n89 4.81523
R5316 VDPWR.n442 VDPWR.n441 4.7505
R5317 VDPWR.n646 VDPWR.n645 4.73979
R5318 VDPWR.n650 VDPWR.n633 4.73979
R5319 VDPWR.n656 VDPWR.n655 4.73979
R5320 VDPWR.n660 VDPWR.n620 4.73979
R5321 VDPWR.n664 VDPWR.n398 4.73798
R5322 VDPWR.n111 VDPWR.n110 4.67238
R5323 VDPWR.n182 VDPWR.n181 4.65675
R5324 VDPWR.n145 VDPWR.n112 4.65675
R5325 VDPWR.n171 VDPWR.n170 4.65675
R5326 VDPWR.n645 VDPWR.n634 4.6505
R5327 VDPWR.n650 VDPWR.n649 4.6505
R5328 VDPWR.n655 VDPWR.n621 4.6505
R5329 VDPWR.n660 VDPWR.n659 4.6505
R5330 VDPWR.n635 VDPWR.n634 4.54311
R5331 VDPWR.n646 VDPWR.n635 4.54311
R5332 VDPWR.n622 VDPWR.n621 4.54311
R5333 VDPWR.n656 VDPWR.n622 4.54311
R5334 VDPWR.n437 VDPWR.n436 4.5005
R5335 VDPWR.n438 VDPWR.n410 4.5005
R5336 VDPWR.n662 VDPWR.n661 4.5005
R5337 VDPWR.n654 VDPWR.n653 4.5005
R5338 VDPWR.n652 VDPWR.n651 4.5005
R5339 VDPWR.n332 VDPWR.n331 4.5005
R5340 VDPWR.n330 VDPWR.n215 4.5005
R5341 VDPWR.n526 VDPWR.n525 4.48641
R5342 VDPWR.n525 VDPWR.n503 4.48641
R5343 VDPWR.n536 VDPWR.n535 4.48641
R5344 VDPWR.n535 VDPWR.n483 4.48641
R5345 VDPWR.n613 VDPWR.n612 4.48641
R5346 VDPWR.n612 VDPWR.n606 4.48641
R5347 VDPWR.n649 VDPWR.n648 4.48641
R5348 VDPWR.n648 VDPWR.n633 4.48641
R5349 VDPWR.n659 VDPWR.n658 4.48641
R5350 VDPWR.n658 VDPWR.n620 4.48641
R5351 VDPWR.n480 VDPWR.n479 4.29244
R5352 VDPWR.n664 VDPWR.n663 3.86809
R5353 VDPWR.n183 VDPWR.n182 3.81758
R5354 VDPWR.n665 VDPWR.n183 3.81656
R5355 VDPWR.n589 VDPWR.n580 3.75335
R5356 VDPWR.n583 VDPWR.n550 3.75335
R5357 VDPWR.n571 VDPWR.n557 3.75335
R5358 VDPWR.n563 VDPWR.n562 3.75335
R5359 VDPWR.n338 VDPWR.n213 3.75335
R5360 VDPWR.n337 VDPWR.n336 3.75335
R5361 VDPWR.n392 VDPWR.n388 3.75335
R5362 VDPWR.n391 VDPWR.n390 3.75335
R5363 VDPWR.n383 VDPWR.n186 3.75335
R5364 VDPWR.n384 VDPWR.n382 3.75335
R5365 VDPWR.n362 VDPWR.n358 3.75335
R5366 VDPWR.n361 VDPWR.n360 3.75335
R5367 VDPWR.n353 VDPWR.n208 3.75335
R5368 VDPWR.n354 VDPWR.n352 3.75335
R5369 VDPWR.n347 VDPWR.n343 3.75335
R5370 VDPWR.n346 VDPWR.n345 3.75335
R5371 VDPWR.n314 VDPWR.n313 3.75335
R5372 VDPWR.n312 VDPWR.n217 3.75335
R5373 VDPWR.n324 VDPWR.n319 3.75335
R5374 VDPWR.n323 VDPWR.n322 3.75335
R5375 VDPWR.n297 VDPWR.n296 3.75335
R5376 VDPWR.n295 VDPWR.n221 3.75335
R5377 VDPWR.n307 VDPWR.n303 3.75335
R5378 VDPWR.n306 VDPWR.n305 3.75335
R5379 VDPWR.n468 VDPWR.n466 3.55702
R5380 VDPWR.n451 VDPWR.n450 3.55702
R5381 VDPWR.n103 VDPWR.n51 3.55702
R5382 VDPWR.n70 VDPWR.n65 3.55702
R5383 VDPWR.n471 VDPWR.n467 3.53508
R5384 VDPWR.n469 VDPWR.n407 3.53508
R5385 VDPWR.n471 VDPWR.n470 3.53508
R5386 VDPWR.n477 VDPWR.n407 3.53508
R5387 VDPWR.n420 VDPWR.n418 3.53508
R5388 VDPWR.n446 VDPWR.n445 3.53508
R5389 VDPWR.n449 VDPWR.n420 3.53508
R5390 VDPWR.n445 VDPWR.n444 3.53508
R5391 VDPWR.n290 VDPWR.n289 3.53508
R5392 VDPWR.n289 VDPWR.n288 3.53508
R5393 VDPWR.n234 VDPWR.n229 3.53508
R5394 VDPWR.n231 VDPWR.n229 3.53508
R5395 VDPWR.n276 VDPWR.n238 3.53508
R5396 VDPWR.n277 VDPWR.n276 3.53508
R5397 VDPWR.n271 VDPWR.n270 3.53508
R5398 VDPWR.n270 VDPWR.n269 3.53508
R5399 VDPWR.n251 VDPWR.n246 3.53508
R5400 VDPWR.n248 VDPWR.n246 3.53508
R5401 VDPWR.n258 VDPWR.n254 3.53508
R5402 VDPWR.n259 VDPWR.n258 3.53508
R5403 VDPWR.n102 VDPWR.n101 3.53508
R5404 VDPWR.n101 VDPWR.n52 3.53508
R5405 VDPWR.n66 VDPWR.n63 3.53508
R5406 VDPWR.n71 VDPWR.n63 3.53508
R5407 VDPWR.n609 VDPWR.n608 3.46433
R5408 VDPWR.n522 VDPWR.n521 3.41464
R5409 VDPWR.n532 VDPWR.n531 3.41464
R5410 VDPWR.n378 VDPWR.n377 3.40194
R5411 VDPWR.n376 VDPWR.n372 3.40194
R5412 VDPWR.n204 VDPWR.n203 3.40194
R5413 VDPWR.n202 VDPWR.n197 3.40194
R5414 VDPWR.n97 VDPWR.n58 3.14514
R5415 VDPWR.n523 VDPWR.n522 3.11118
R5416 VDPWR.n533 VDPWR.n532 3.11118
R5417 VDPWR.n87 VDPWR.n86 3.1005
R5418 VDPWR.n60 VDPWR.n58 3.1005
R5419 VDPWR.n89 VDPWR.n88 3.1005
R5420 VDPWR.n522 VDPWR.n504 3.04304
R5421 VDPWR.n532 VDPWR.n484 3.04304
R5422 VDPWR.n610 VDPWR.n609 2.96855
R5423 VDPWR.n609 VDPWR.n607 2.90353
R5424 VDPWR.n473 VDPWR.n466 2.60059
R5425 VDPWR.n452 VDPWR.n451 2.60059
R5426 VDPWR.n104 VDPWR.n103 2.60059
R5427 VDPWR.n76 VDPWR.n65 2.60059
R5428 VDPWR.n467 VDPWR.n466 2.55763
R5429 VDPWR.n451 VDPWR.n418 2.55763
R5430 VDPWR.n103 VDPWR.n102 2.55763
R5431 VDPWR.n66 VDPWR.n65 2.55763
R5432 VDPWR.n377 VDPWR.n193 2.39444
R5433 VDPWR.n376 VDPWR.n375 2.39444
R5434 VDPWR.n203 VDPWR.n196 2.39444
R5435 VDPWR.n202 VDPWR.n201 2.39444
R5436 VDPWR.n372 VDPWR.n371 2.32777
R5437 VDPWR.n205 VDPWR.n204 2.32777
R5438 VDPWR.n96 VDPWR.n60 2.27782
R5439 VDPWR.n84 VDPWR.n60 2.27782
R5440 VDPWR.n88 VDPWR.n61 2.27782
R5441 VDPWR.n86 VDPWR.n84 2.27782
R5442 VDPWR.n97 VDPWR.n96 2.27782
R5443 VDPWR.n86 VDPWR.n61 2.27782
R5444 VDPWR.n183 VDPWR.n111 2.13269
R5445 VDPWR.n608 VDPWR.n605 1.94497
R5446 VDPWR.n616 VDPWR.n615 1.94497
R5447 VDPWR.n521 VDPWR.n520 1.90331
R5448 VDPWR.n403 VDPWR.n402 1.88999
R5449 VDPWR.n529 VDPWR.n528 1.77831
R5450 VDPWR.n531 VDPWR.n530 1.77831
R5451 VDPWR.n539 VDPWR.n538 1.77831
R5452 VDPWR.n617 VDPWR.n616 1.50847
R5453 VDPWR.n540 VDPWR.n539 1.49285
R5454 VDPWR.n369 VDPWR.n368 1.15675
R5455 VDPWR.n398 VDPWR.n184 1.15675
R5456 VDPWR.n43 VDPWR.n42 1.10988
R5457 VDPWR.n40 VDPWR.n1 1.04738
R5458 VDPWR.n30 VDPWR.n28 0.96925
R5459 VDPWR.n11 VDPWR.n10 0.938
R5460 VDPWR.n18 VDPWR.n16 0.938
R5461 VDPWR.n23 VDPWR.n22 0.938
R5462 VDPWR.n653 VDPWR.n652 0.90675
R5463 VDPWR.n42 VDPWR.n40 0.891125
R5464 VDPWR.n171 VDPWR.n112 0.813
R5465 VDPWR.n182 VDPWR.n112 0.813
R5466 VDPWR.n174 VDPWR.n173 0.8005
R5467 VDPWR.n401 VDPWR.n400 0.75233
R5468 VDPWR.n33 VDPWR.n32 0.734875
R5469 VDPWR.n284 VDPWR.n216 0.688
R5470 VDPWR.n81 VDPWR.n79 0.688
R5471 VDPWR.n83 VDPWR.n81 0.688
R5472 VDPWR.n93 VDPWR.n92 0.688
R5473 VDPWR.n92 VDPWR.n50 0.688
R5474 VDPWR.n32 VDPWR.n30 0.688
R5475 VDPWR.n38 VDPWR.n36 0.688
R5476 VDPWR.n43 VDPWR.n38 0.672375
R5477 VDPWR.n48 VDPWR.n1 0.65675
R5478 VDPWR.n402 VDPWR.n401 0.648711
R5479 VDPWR.n437 VDPWR.n434 0.6255
R5480 VDPWR.n434 VDPWR.n432 0.6255
R5481 VDPWR.n432 VDPWR.n405 0.6255
R5482 VDPWR.n284 VDPWR.n283 0.609875
R5483 VDPWR.n10 VDPWR.n5 0.563
R5484 VDPWR.n20 VDPWR.n18 0.563
R5485 VDPWR.n22 VDPWR.n3 0.563
R5486 VDPWR.n11 VDPWR.n8 0.53175
R5487 VDPWR.n16 VDPWR.n5 0.53175
R5488 VDPWR.n23 VDPWR.n20 0.53175
R5489 VDPWR.n28 VDPWR.n3 0.53175
R5490 VDPWR.n329 VDPWR.n216 0.516125
R5491 VDPWR.n440 VDPWR.n438 0.5005
R5492 VDPWR.n90 VDPWR.n83 0.5005
R5493 VDPWR.n93 VDPWR.n90 0.5005
R5494 VDPWR.n368 VDPWR.n206 0.391125
R5495 VDPWR.n36 VDPWR.n34 0.391125
R5496 VDPWR.n662 VDPWR.n619 0.34425
R5497 VDPWR.n624 VDPWR.n619 0.34425
R5498 VDPWR.n626 VDPWR.n624 0.34425
R5499 VDPWR.n628 VDPWR.n626 0.34425
R5500 VDPWR.n630 VDPWR.n628 0.34425
R5501 VDPWR.n653 VDPWR.n630 0.34425
R5502 VDPWR.n652 VDPWR.n632 0.34425
R5503 VDPWR.n637 VDPWR.n632 0.34425
R5504 VDPWR.n639 VDPWR.n637 0.34425
R5505 VDPWR.n641 VDPWR.n639 0.34425
R5506 VDPWR.n643 VDPWR.n641 0.34425
R5507 VDPWR.n111 VDPWR.n50 0.34425
R5508 VDPWR.n34 VDPWR.n33 0.34425
R5509 VDPWR.n530 VDPWR.n529 0.333833
R5510 VDPWR.n605 VDPWR.n604 0.328625
R5511 VDPWR.n283 VDPWR.n236 0.328625
R5512 VDPWR.n330 VDPWR.n329 0.328625
R5513 VDPWR.n441 VDPWR.n440 0.313
R5514 VDPWR.n479 VDPWR.n405 0.313
R5515 VDPWR.n331 VDPWR.n206 0.297375
R5516 VDPWR VDPWR.n666 0.295024
R5517 VDPWR.n617 VDPWR.n540 0.285347
R5518 VDPWR.n265 VDPWR.n236 0.28175
R5519 VDPWR.n528 VDPWR.n527 0.2505
R5520 VDPWR.n538 VDPWR.n537 0.2505
R5521 VDPWR.n369 VDPWR.n184 0.2505
R5522 VDPWR.n181 VDPWR.n128 0.2505
R5523 VDPWR.n145 VDPWR.n144 0.2505
R5524 VDPWR.n170 VDPWR.n169 0.2505
R5525 VDPWR.n615 VDPWR.n614 0.229667
R5526 VDPWR.n616 VDPWR.n605 0.229667
R5527 VDPWR.n572 VDPWR.n558 0.208833
R5528 VDPWR.n566 VDPWR.n558 0.208833
R5529 VDPWR.n566 VDPWR.n565 0.208833
R5530 VDPWR.n581 VDPWR.n579 0.208833
R5531 VDPWR.n582 VDPWR.n581 0.208833
R5532 VDPWR.n582 VDPWR.n551 0.208833
R5533 VDPWR.n122 VDPWR.n115 0.208833
R5534 VDPWR.n118 VDPWR.n115 0.208833
R5535 VDPWR.n118 VDPWR.n117 0.208833
R5536 VDPWR.n128 VDPWR.n113 0.208833
R5537 VDPWR.n124 VDPWR.n113 0.208833
R5538 VDPWR.n124 VDPWR.n123 0.208833
R5539 VDPWR.n138 VDPWR.n131 0.208833
R5540 VDPWR.n134 VDPWR.n131 0.208833
R5541 VDPWR.n134 VDPWR.n133 0.208833
R5542 VDPWR.n144 VDPWR.n129 0.208833
R5543 VDPWR.n140 VDPWR.n129 0.208833
R5544 VDPWR.n140 VDPWR.n139 0.208833
R5545 VDPWR.n163 VDPWR.n156 0.208833
R5546 VDPWR.n159 VDPWR.n156 0.208833
R5547 VDPWR.n159 VDPWR.n158 0.208833
R5548 VDPWR.n169 VDPWR.n154 0.208833
R5549 VDPWR.n165 VDPWR.n154 0.208833
R5550 VDPWR.n165 VDPWR.n164 0.208833
R5551 VDPWR.n480 VDPWR.n403 0.20853
R5552 VDPWR.n443 VDPWR.n442 0.188
R5553 VDPWR.n604 VDPWR.n603 0.188
R5554 VDPWR.n603 VDPWR.n602 0.188
R5555 VDPWR.n602 VDPWR.n601 0.188
R5556 VDPWR.n601 VDPWR.n600 0.188
R5557 VDPWR.n600 VDPWR.n599 0.188
R5558 VDPWR.n599 VDPWR.n598 0.188
R5559 VDPWR.n598 VDPWR.n597 0.188
R5560 VDPWR.n597 VDPWR.n596 0.188
R5561 VDPWR.n110 VDPWR.n109 0.188
R5562 VDPWR.n69 VDPWR.n62 0.188
R5563 VDPWR.n666 VDPWR.n665 0.183005
R5564 VDPWR.n651 VDPWR.n650 0.182048
R5565 VDPWR.n661 VDPWR.n660 0.182048
R5566 VDPWR.n645 VDPWR.n644 0.182048
R5567 VDPWR.n655 VDPWR.n654 0.182048
R5568 VDPWR.n665 VDPWR.n664 0.178305
R5569 VDPWR.t211 VDPWR.t88 0.1603
R5570 VDPWR.t207 VDPWR.t211 0.1603
R5571 VDPWR.t360 VDPWR.t207 0.1603
R5572 VDPWR.t392 VDPWR.t360 0.1603
R5573 VDPWR.t79 VDPWR.t392 0.1603
R5574 VDPWR.t359 VDPWR.t79 0.1603
R5575 VDPWR.t241 VDPWR.t359 0.1603
R5576 VDPWR.t107 VDPWR.t241 0.1603
R5577 VDPWR.t108 VDPWR.t48 0.1603
R5578 VDPWR.t46 VDPWR.t108 0.1603
R5579 VDPWR.t373 VDPWR.t46 0.1603
R5580 VDPWR.t414 VDPWR.t373 0.1603
R5581 VDPWR.t393 VDPWR.t414 0.1603
R5582 VDPWR.t374 VDPWR.t393 0.1603
R5583 VDPWR.t208 VDPWR.t374 0.1603
R5584 VDPWR.t133 VDPWR.t208 0.1603
R5585 VDPWR.t78 VDPWR.n399 0.159278
R5586 VDPWR.n468 VDPWR.n406 0.15675
R5587 VDPWR.n450 VDPWR.n419 0.15675
R5588 VDPWR.n443 VDPWR.n419 0.15675
R5589 VDPWR.n109 VDPWR.n51 0.15675
R5590 VDPWR.n70 VDPWR.n69 0.15675
R5591 VDPWR.t48 VDPWR.t78 0.137822
R5592 VDPWR.n399 VDPWR.t107 0.1368
R5593 VDPWR.n436 VDPWR.n410 0.1255
R5594 VDPWR.n438 VDPWR.n437 0.1255
R5595 VDPWR.n539 VDPWR.n482 0.1255
R5596 VDPWR.n486 VDPWR.n482 0.1255
R5597 VDPWR.n488 VDPWR.n486 0.1255
R5598 VDPWR.n490 VDPWR.n488 0.1255
R5599 VDPWR.n492 VDPWR.n490 0.1255
R5600 VDPWR.n494 VDPWR.n492 0.1255
R5601 VDPWR.n496 VDPWR.n494 0.1255
R5602 VDPWR.n498 VDPWR.n496 0.1255
R5603 VDPWR.n500 VDPWR.n498 0.1255
R5604 VDPWR.n530 VDPWR.n500 0.1255
R5605 VDPWR.n529 VDPWR.n502 0.1255
R5606 VDPWR.n506 VDPWR.n502 0.1255
R5607 VDPWR.n508 VDPWR.n506 0.1255
R5608 VDPWR.n510 VDPWR.n508 0.1255
R5609 VDPWR.n512 VDPWR.n510 0.1255
R5610 VDPWR.n514 VDPWR.n512 0.1255
R5611 VDPWR.n516 VDPWR.n514 0.1255
R5612 VDPWR.n518 VDPWR.n516 0.1255
R5613 VDPWR.n520 VDPWR.n518 0.1255
R5614 VDPWR.n332 VDPWR.n215 0.1255
R5615 VDPWR.n331 VDPWR.n330 0.1255
R5616 VDPWR.n540 VDPWR.n480 0.118442
R5617 VDPWR.n663 VDPWR.n617 0.10278
R5618 VDPWR.n87 VDPWR.n58 0.0451429
R5619 VDPWR.n89 VDPWR.n87 0.0451429
R5620 VDPWR.n399 VDPWR.t47 0.00152174
R5621 a_18930_3150.n5 a_18930_3150.t0 752.333
R5622 a_18930_3150.n4 a_18930_3150.t1 752.333
R5623 a_18930_3150.n0 a_18930_3150.t4 514.134
R5624 a_18930_3150.n3 a_18930_3150.n2 366.856
R5625 a_18930_3150.t2 a_18930_3150.n5 254.333
R5626 a_18930_3150.n3 a_18930_3150.t3 190.123
R5627 a_18930_3150.n4 a_18930_3150.n3 187.201
R5628 a_18930_3150.n2 a_18930_3150.n1 176.733
R5629 a_18930_3150.n1 a_18930_3150.n0 176.733
R5630 a_18930_3150.n0 a_18930_3150.t6 112.468
R5631 a_18930_3150.n1 a_18930_3150.t5 112.468
R5632 a_18930_3150.n2 a_18930_3150.t7 112.468
R5633 a_18930_3150.n5 a_18930_3150.n4 70.4005
R5634 a_19250_3100.n0 a_19250_3100.t1 713.933
R5635 a_19250_3100.t0 a_19250_3100.n0 337
R5636 a_19250_3100.n0 a_19250_3100.t2 314.233
R5637 a_19550_2800.t0 a_19550_2800.t1 96.0005
R5638 a_11200_9430.n1 a_11200_9430.t20 312.798
R5639 a_11200_9430.n8 a_11200_9430.t15 312.781
R5640 a_11200_9430.n14 a_11200_9430.t37 312.5
R5641 a_11200_9430.n8 a_11200_9430.t28 310.401
R5642 a_11200_9430.n9 a_11200_9430.t32 310.401
R5643 a_11200_9430.n10 a_11200_9430.t36 310.401
R5644 a_11200_9430.n11 a_11200_9430.t42 310.401
R5645 a_11200_9430.n12 a_11200_9430.t21 310.401
R5646 a_11200_9430.n13 a_11200_9430.t33 310.401
R5647 a_11200_9430.n5 a_11200_9430.t26 310.401
R5648 a_11200_9430.n4 a_11200_9430.t41 310.401
R5649 a_11200_9430.n3 a_11200_9430.t45 310.401
R5650 a_11200_9430.n2 a_11200_9430.t47 310.401
R5651 a_11200_9430.n1 a_11200_9430.t16 310.401
R5652 a_11200_9430.n16 a_11200_9430.t44 308
R5653 a_11200_9430.n28 a_11200_9430.n26 306.808
R5654 a_11200_9430.n0 a_11200_9430.t46 305.901
R5655 a_11200_9430.n20 a_11200_9430.n19 301.933
R5656 a_11200_9430.n22 a_11200_9430.n21 301.933
R5657 a_11200_9430.n24 a_11200_9430.n23 301.933
R5658 a_11200_9430.n29 a_11200_9430.n25 297.433
R5659 a_11200_9430.n28 a_11200_9430.n27 297.433
R5660 a_11200_9430.t2 a_11200_9430.n50 108.898
R5661 a_11200_9430.n18 a_11200_9430.t10 98.9217
R5662 a_11200_9430.n25 a_11200_9430.t6 39.4005
R5663 a_11200_9430.n25 a_11200_9430.t0 39.4005
R5664 a_11200_9430.n26 a_11200_9430.t11 39.4005
R5665 a_11200_9430.n26 a_11200_9430.t7 39.4005
R5666 a_11200_9430.n27 a_11200_9430.t9 39.4005
R5667 a_11200_9430.n27 a_11200_9430.t12 39.4005
R5668 a_11200_9430.n19 a_11200_9430.t13 39.4005
R5669 a_11200_9430.n19 a_11200_9430.t8 39.4005
R5670 a_11200_9430.n21 a_11200_9430.t4 39.4005
R5671 a_11200_9430.n21 a_11200_9430.t3 39.4005
R5672 a_11200_9430.n23 a_11200_9430.t5 39.4005
R5673 a_11200_9430.n23 a_11200_9430.t1 39.4005
R5674 a_11200_9430.n50 a_11200_9430.n30 13.563
R5675 a_11200_9430.n50 a_11200_9430.n49 12.3446
R5676 a_11200_9430.n20 a_11200_9430.n18 4.90675
R5677 a_11200_9430.n31 a_11200_9430.t17 4.8248
R5678 a_11200_9430.n6 a_11200_9430.n0 4.5005
R5679 a_11200_9430.n17 a_11200_9430.n7 4.5005
R5680 a_11200_9430.n16 a_11200_9430.n15 4.5005
R5681 a_11200_9430.n30 a_11200_9430.n29 4.5005
R5682 a_11200_9430.n39 a_11200_9430.t22 4.5005
R5683 a_11200_9430.n38 a_11200_9430.t49 4.5005
R5684 a_11200_9430.n37 a_11200_9430.t39 4.5005
R5685 a_11200_9430.n36 a_11200_9430.t29 4.5005
R5686 a_11200_9430.n35 a_11200_9430.t34 4.5005
R5687 a_11200_9430.n34 a_11200_9430.t40 4.5005
R5688 a_11200_9430.n33 a_11200_9430.t31 4.5005
R5689 a_11200_9430.n32 a_11200_9430.t35 4.5005
R5690 a_11200_9430.n31 a_11200_9430.t25 4.5005
R5691 a_11200_9430.n40 a_11200_9430.t48 4.5005
R5692 a_11200_9430.n41 a_11200_9430.t38 4.5005
R5693 a_11200_9430.n42 a_11200_9430.t27 4.5005
R5694 a_11200_9430.n43 a_11200_9430.t18 4.5005
R5695 a_11200_9430.n44 a_11200_9430.t23 4.5005
R5696 a_11200_9430.n45 a_11200_9430.t30 4.5005
R5697 a_11200_9430.n46 a_11200_9430.t19 4.5005
R5698 a_11200_9430.n47 a_11200_9430.t24 4.5005
R5699 a_11200_9430.n48 a_11200_9430.t14 4.5005
R5700 a_11200_9430.n49 a_11200_9430.t43 4.5005
R5701 a_11200_9430.n29 a_11200_9430.n28 1.59425
R5702 a_11200_9430.n18 a_11200_9430.n17 1.21925
R5703 a_11200_9430.n30 a_11200_9430.n24 1.1255
R5704 a_11200_9430.n24 a_11200_9430.n22 1.1255
R5705 a_11200_9430.n22 a_11200_9430.n20 1.1255
R5706 a_11200_9430.n39 a_11200_9430.n38 0.3295
R5707 a_11200_9430.n38 a_11200_9430.n37 0.3295
R5708 a_11200_9430.n37 a_11200_9430.n36 0.3295
R5709 a_11200_9430.n36 a_11200_9430.n35 0.3295
R5710 a_11200_9430.n35 a_11200_9430.n34 0.3295
R5711 a_11200_9430.n34 a_11200_9430.n33 0.3295
R5712 a_11200_9430.n33 a_11200_9430.n32 0.3295
R5713 a_11200_9430.n32 a_11200_9430.n31 0.3295
R5714 a_11200_9430.n41 a_11200_9430.n40 0.3295
R5715 a_11200_9430.n42 a_11200_9430.n41 0.3295
R5716 a_11200_9430.n43 a_11200_9430.n42 0.3295
R5717 a_11200_9430.n44 a_11200_9430.n43 0.3295
R5718 a_11200_9430.n45 a_11200_9430.n44 0.3295
R5719 a_11200_9430.n46 a_11200_9430.n45 0.3295
R5720 a_11200_9430.n47 a_11200_9430.n46 0.3295
R5721 a_11200_9430.n48 a_11200_9430.n47 0.3295
R5722 a_11200_9430.n49 a_11200_9430.n48 0.3248
R5723 a_11200_9430.n40 a_11200_9430.n39 0.2825
R5724 a_11200_9430.n2 a_11200_9430.n1 0.28175
R5725 a_11200_9430.n3 a_11200_9430.n2 0.28175
R5726 a_11200_9430.n4 a_11200_9430.n3 0.28175
R5727 a_11200_9430.n5 a_11200_9430.n4 0.28175
R5728 a_11200_9430.n6 a_11200_9430.n5 0.28175
R5729 a_11200_9430.n15 a_11200_9430.n14 0.28175
R5730 a_11200_9430.n14 a_11200_9430.n13 0.28175
R5731 a_11200_9430.n13 a_11200_9430.n12 0.28175
R5732 a_11200_9430.n12 a_11200_9430.n11 0.28175
R5733 a_11200_9430.n11 a_11200_9430.n10 0.28175
R5734 a_11200_9430.n10 a_11200_9430.n9 0.28175
R5735 a_11200_9430.n9 a_11200_9430.n8 0.28175
R5736 a_11200_9430.n7 a_11200_9430.n6 0.141125
R5737 a_11200_9430.n15 a_11200_9430.n7 0.141125
R5738 a_11200_9430.n17 a_11200_9430.n0 0.141125
R5739 a_11200_9430.n17 a_11200_9430.n16 0.141125
R5740 a_11780_7290.n2 a_11780_7290.n0 1319.38
R5741 a_11780_7290.t6 a_11780_7290.t4 1188.93
R5742 a_11780_7290.t4 a_11780_7290.t5 835.467
R5743 a_11780_7290.n0 a_11780_7290.t3 562.333
R5744 a_11780_7290.n2 a_11780_7290.n1 247.917
R5745 a_11780_7290.n0 a_11780_7290.t6 224.934
R5746 a_11780_7290.t1 a_11780_7290.n2 221.411
R5747 a_11780_7290.n1 a_11780_7290.t2 24.0005
R5748 a_11780_7290.n1 a_11780_7290.t0 24.0005
R5749 a_12300_6670.t0 a_12300_6670.t1 39.4005
R5750 a_12070_2860.n4 a_12070_2860.n3 919.244
R5751 a_12070_2860.n9 a_12070_2860.n8 918.702
R5752 a_12070_2860.t10 a_12070_2860.t8 819.4
R5753 a_12070_2860.n10 a_12070_2860.n0 628.734
R5754 a_12070_2860.n3 a_12070_2860.n2 520.361
R5755 a_12070_2860.n8 a_12070_2860.n7 364.178
R5756 a_12070_2860.n1 a_12070_2860.t5 337.401
R5757 a_12070_2860.n9 a_12070_2860.t10 336.25
R5758 a_12070_2860.n1 a_12070_2860.t12 305.267
R5759 a_12070_2860.t0 a_12070_2860.n10 257.534
R5760 a_12070_2860.n5 a_12070_2860.t9 192.8
R5761 a_12070_2860.n2 a_12070_2860.n1 176.733
R5762 a_12070_2860.n7 a_12070_2860.n6 176.733
R5763 a_12070_2860.n5 a_12070_2860.n4 160.667
R5764 a_12070_2860.n4 a_12070_2860.t14 144.601
R5765 a_12070_2860.n3 a_12070_2860.t3 131.976
R5766 a_12070_2860.n1 a_12070_2860.t4 128.534
R5767 a_12070_2860.n2 a_12070_2860.t11 128.534
R5768 a_12070_2860.n6 a_12070_2860.t13 112.468
R5769 a_12070_2860.n7 a_12070_2860.t6 112.468
R5770 a_12070_2860.n8 a_12070_2860.t7 112.468
R5771 a_12070_2860.n6 a_12070_2860.n5 96.4005
R5772 a_12070_2860.n0 a_12070_2860.t1 78.8005
R5773 a_12070_2860.n0 a_12070_2860.t2 78.8005
R5774 a_12070_2860.n10 a_12070_2860.n9 11.2005
R5775 a_12870_2890.t0 a_12870_2890.t1 96.0005
R5776 a_12290_3150.n1 a_12290_3150.t1 685.134
R5777 a_12290_3150.n0 a_12290_3150.t0 685.134
R5778 a_12290_3150.n0 a_12290_3150.t3 534.268
R5779 a_12290_3150.t2 a_12290_3150.n1 340.521
R5780 a_12290_3150.n1 a_12290_3150.n0 105.6
R5781 a_18330_3180.t2 a_18330_3180.t4 1012.2
R5782 a_18330_3180.n0 a_18330_3180.t0 663.801
R5783 a_18330_3180.n2 a_18330_3180.n1 431.401
R5784 a_18330_3180.t3 a_18330_3180.t5 401.668
R5785 a_18330_3180.n0 a_18330_3180.t2 361.692
R5786 a_18330_3180.n1 a_18330_3180.t6 353.467
R5787 a_18330_3180.t1 a_18330_3180.n2 298.921
R5788 a_18330_3180.n1 a_18330_3180.t3 257.067
R5789 a_18330_3180.n2 a_18330_3180.n0 67.2005
R5790 a_9570_16200.n6 a_9570_16200.t9 287.762
R5791 a_9570_16200.n5 a_9570_16200.t7 287.762
R5792 a_9570_16200.n5 a_9570_16200.t10 287.589
R5793 a_9570_16200.n8 a_9570_16200.t11 287.012
R5794 a_9570_16200.n7 a_9570_16200.t8 287.012
R5795 a_9570_16200.t6 a_9570_16200.n9 115.097
R5796 a_9570_16200.n2 a_9570_16200.n0 107.266
R5797 a_9570_16200.n4 a_9570_16200.n3 105.016
R5798 a_9570_16200.n2 a_9570_16200.n1 105.016
R5799 a_9570_16200.n3 a_9570_16200.t3 13.1338
R5800 a_9570_16200.n3 a_9570_16200.t4 13.1338
R5801 a_9570_16200.n1 a_9570_16200.t0 13.1338
R5802 a_9570_16200.n1 a_9570_16200.t1 13.1338
R5803 a_9570_16200.n0 a_9570_16200.t5 13.1338
R5804 a_9570_16200.n0 a_9570_16200.t2 13.1338
R5805 a_9570_16200.n9 a_9570_16200.n4 9.0005
R5806 a_9570_16200.n9 a_9570_16200.n8 6.78086
R5807 a_9570_16200.n4 a_9570_16200.n2 2.2505
R5808 a_9570_16200.n7 a_9570_16200.n6 0.579071
R5809 a_9570_16200.n8 a_9570_16200.n7 0.282643
R5810 a_9570_16200.n6 a_9570_16200.n5 0.2755
R5811 a_9450_16252.n0 a_9450_16252.t11 403.952
R5812 a_9450_16252.n18 a_9450_16252.t27 403.755
R5813 a_9450_16252.n17 a_9450_16252.t16 403.755
R5814 a_9450_16252.n16 a_9450_16252.t24 403.755
R5815 a_9450_16252.n15 a_9450_16252.t14 403.755
R5816 a_9450_16252.n14 a_9450_16252.t22 403.755
R5817 a_9450_16252.n13 a_9450_16252.t12 403.755
R5818 a_9450_16252.n12 a_9450_16252.t18 403.755
R5819 a_9450_16252.n11 a_9450_16252.t25 403.755
R5820 a_9450_16252.n10 a_9450_16252.t21 403.755
R5821 a_9450_16252.n9 a_9450_16252.t10 403.755
R5822 a_9450_16252.n8 a_9450_16252.t29 403.755
R5823 a_9450_16252.n7 a_9450_16252.t19 403.755
R5824 a_9450_16252.n6 a_9450_16252.t26 403.755
R5825 a_9450_16252.n5 a_9450_16252.t15 403.755
R5826 a_9450_16252.n4 a_9450_16252.t23 403.755
R5827 a_9450_16252.n3 a_9450_16252.t13 403.755
R5828 a_9450_16252.n2 a_9450_16252.t20 403.755
R5829 a_9450_16252.n1 a_9450_16252.t28 403.755
R5830 a_9450_16252.n0 a_9450_16252.t17 403.755
R5831 a_9450_16252.n26 a_9450_16252.n25 301.933
R5832 a_9450_16252.n24 a_9450_16252.n23 301.933
R5833 a_9450_16252.n22 a_9450_16252.n21 301.933
R5834 a_9450_16252.n20 a_9450_16252.n19 301.933
R5835 a_9450_16252.t2 a_9450_16252.n27 117.008
R5836 a_9450_16252.n20 a_9450_16252.t6 103.828
R5837 a_9450_16252.n25 a_9450_16252.t1 39.4005
R5838 a_9450_16252.n25 a_9450_16252.t4 39.4005
R5839 a_9450_16252.n23 a_9450_16252.t8 39.4005
R5840 a_9450_16252.n23 a_9450_16252.t3 39.4005
R5841 a_9450_16252.n21 a_9450_16252.t0 39.4005
R5842 a_9450_16252.n21 a_9450_16252.t7 39.4005
R5843 a_9450_16252.n19 a_9450_16252.t5 39.4005
R5844 a_9450_16252.n19 a_9450_16252.t9 39.4005
R5845 a_9450_16252.n27 a_9450_16252.n18 10.3335
R5846 a_9450_16252.n27 a_9450_16252.n26 5.313
R5847 a_9450_16252.n9 a_9450_16252.n8 1.6255
R5848 a_9450_16252.n22 a_9450_16252.n20 1.1255
R5849 a_9450_16252.n24 a_9450_16252.n22 1.1255
R5850 a_9450_16252.n26 a_9450_16252.n24 1.1255
R5851 a_9450_16252.n1 a_9450_16252.n0 0.196929
R5852 a_9450_16252.n2 a_9450_16252.n1 0.196929
R5853 a_9450_16252.n3 a_9450_16252.n2 0.196929
R5854 a_9450_16252.n4 a_9450_16252.n3 0.196929
R5855 a_9450_16252.n5 a_9450_16252.n4 0.196929
R5856 a_9450_16252.n6 a_9450_16252.n5 0.196929
R5857 a_9450_16252.n7 a_9450_16252.n6 0.196929
R5858 a_9450_16252.n8 a_9450_16252.n7 0.196929
R5859 a_9450_16252.n10 a_9450_16252.n9 0.196929
R5860 a_9450_16252.n11 a_9450_16252.n10 0.196929
R5861 a_9450_16252.n12 a_9450_16252.n11 0.196929
R5862 a_9450_16252.n13 a_9450_16252.n12 0.196929
R5863 a_9450_16252.n14 a_9450_16252.n13 0.196929
R5864 a_9450_16252.n15 a_9450_16252.n14 0.196929
R5865 a_9450_16252.n16 a_9450_16252.n15 0.196929
R5866 a_9450_16252.n17 a_9450_16252.n16 0.196929
R5867 a_9450_16252.n18 a_9450_16252.n17 0.196929
R5868 a_10480_13480.n0 a_10480_13480.t6 238.322
R5869 a_10480_13480.n0 a_10480_13480.t7 238.322
R5870 a_10480_13480.n4 a_10480_13480.n0 168.8
R5871 a_10480_13480.n1 a_10480_13480.t1 130.001
R5872 a_10480_13480.n3 a_10480_13480.n2 105.171
R5873 a_10480_13480.n5 a_10480_13480.n4 105.171
R5874 a_10480_13480.n1 a_10480_13480.t0 81.7085
R5875 a_10480_13480.n3 a_10480_13480.n1 46.5739
R5876 a_10480_13480.n2 a_10480_13480.t3 13.1338
R5877 a_10480_13480.n2 a_10480_13480.t4 13.1338
R5878 a_10480_13480.t5 a_10480_13480.n5 13.1338
R5879 a_10480_13480.n5 a_10480_13480.t2 13.1338
R5880 a_10480_13480.n4 a_10480_13480.n3 3.3755
R5881 a_9450_17070.t6 a_9450_17070.t13 138.543
R5882 a_9450_17070.t20 a_9450_17070.t8 0.1603
R5883 a_9450_17070.t4 a_9450_17070.t20 0.1603
R5884 a_9450_17070.t18 a_9450_17070.t4 0.1603
R5885 a_9450_17070.t7 a_9450_17070.t18 0.1603
R5886 a_9450_17070.t5 a_9450_17070.t7 0.1603
R5887 a_9450_17070.t16 a_9450_17070.t5 0.1603
R5888 a_9450_17070.t15 a_9450_17070.t16 0.1603
R5889 a_9450_17070.t12 a_9450_17070.t15 0.1603
R5890 a_9450_17070.t9 a_9450_17070.t14 0.1603
R5891 a_9450_17070.t17 a_9450_17070.t9 0.1603
R5892 a_9450_17070.t2 a_9450_17070.t17 0.1603
R5893 a_9450_17070.t10 a_9450_17070.t2 0.1603
R5894 a_9450_17070.t19 a_9450_17070.t10 0.1603
R5895 a_9450_17070.t3 a_9450_17070.t19 0.1603
R5896 a_9450_17070.t11 a_9450_17070.t3 0.1603
R5897 a_9450_17070.t13 a_9450_17070.t11 0.1603
R5898 a_9450_17070.t0 a_9450_17070.n0 0.159278
R5899 a_9450_17070.t14 a_9450_17070.t0 0.137822
R5900 a_9450_17070.n0 a_9450_17070.t12 0.1368
R5901 a_9450_17070.n0 a_9450_17070.t1 0.00152174
R5902 a_13200_10990.n15 a_13200_10990.t21 310.488
R5903 a_13200_10990.n9 a_13200_10990.t22 310.488
R5904 a_13200_10990.n4 a_13200_10990.t20 310.488
R5905 a_13200_10990.n13 a_13200_10990.n12 297.433
R5906 a_13200_10990.n8 a_13200_10990.n7 297.433
R5907 a_13200_10990.n19 a_13200_10990.n18 297.433
R5908 a_13200_10990.n2 a_13200_10990.t16 248.133
R5909 a_13200_10990.n2 a_13200_10990.n1 199.383
R5910 a_13200_10990.n3 a_13200_10990.n0 194.883
R5911 a_13200_10990.n17 a_13200_10990.t10 184.097
R5912 a_13200_10990.n11 a_13200_10990.t6 184.097
R5913 a_13200_10990.n6 a_13200_10990.t8 184.097
R5914 a_13200_10990.n16 a_13200_10990.n15 167.094
R5915 a_13200_10990.n10 a_13200_10990.n9 167.094
R5916 a_13200_10990.n5 a_13200_10990.n4 167.094
R5917 a_13200_10990.n18 a_13200_10990.n17 161.3
R5918 a_13200_10990.n13 a_13200_10990.n11 161.3
R5919 a_13200_10990.n8 a_13200_10990.n6 161.3
R5920 a_13200_10990.n15 a_13200_10990.t18 120.501
R5921 a_13200_10990.n16 a_13200_10990.t2 120.501
R5922 a_13200_10990.n9 a_13200_10990.t19 120.501
R5923 a_13200_10990.n10 a_13200_10990.t0 120.501
R5924 a_13200_10990.n4 a_13200_10990.t17 120.501
R5925 a_13200_10990.n5 a_13200_10990.t4 120.501
R5926 a_13200_10990.n1 a_13200_10990.t13 48.0005
R5927 a_13200_10990.n1 a_13200_10990.t12 48.0005
R5928 a_13200_10990.n0 a_13200_10990.t15 48.0005
R5929 a_13200_10990.n0 a_13200_10990.t14 48.0005
R5930 a_13200_10990.n17 a_13200_10990.n16 40.7027
R5931 a_13200_10990.n11 a_13200_10990.n10 40.7027
R5932 a_13200_10990.n6 a_13200_10990.n5 40.7027
R5933 a_13200_10990.n12 a_13200_10990.t7 39.4005
R5934 a_13200_10990.n12 a_13200_10990.t1 39.4005
R5935 a_13200_10990.n7 a_13200_10990.t9 39.4005
R5936 a_13200_10990.n7 a_13200_10990.t5 39.4005
R5937 a_13200_10990.t11 a_13200_10990.n19 39.4005
R5938 a_13200_10990.n19 a_13200_10990.t3 39.4005
R5939 a_13200_10990.n14 a_13200_10990.n13 6.6255
R5940 a_13200_10990.n14 a_13200_10990.n8 6.6255
R5941 a_13200_10990.n3 a_13200_10990.n2 5.2505
R5942 a_13200_10990.n18 a_13200_10990.n14 4.5005
R5943 a_13200_10990.n18 a_13200_10990.n3 0.78175
R5944 a_10000_15820.n3 a_10000_15820.t6 291.502
R5945 a_10000_15820.n3 a_10000_15820.t9 291.288
R5946 a_10000_15820.n4 a_10000_15820.t7 291.288
R5947 a_10000_15820.n5 a_10000_15820.t8 291.288
R5948 a_10000_15820.n6 a_10000_15820.t10 291.288
R5949 a_10000_15820.n8 a_10000_15820.t5 148.653
R5950 a_10000_15820.t0 a_10000_15820.n8 125.371
R5951 a_10000_15820.n2 a_10000_15820.n0 105.609
R5952 a_10000_15820.n2 a_10000_15820.n1 104.484
R5953 a_10000_15820.n8 a_10000_15820.n7 21.4246
R5954 a_10000_15820.n7 a_10000_15820.n2 14.2349
R5955 a_10000_15820.n0 a_10000_15820.t2 13.1338
R5956 a_10000_15820.n0 a_10000_15820.t4 13.1338
R5957 a_10000_15820.n1 a_10000_15820.t3 13.1338
R5958 a_10000_15820.n1 a_10000_15820.t1 13.1338
R5959 a_10000_15820.n7 a_10000_15820.n6 6.43621
R5960 a_10000_15820.n6 a_10000_15820.n5 0.643357
R5961 a_10000_15820.n4 a_10000_15820.n3 0.643357
R5962 a_10000_15820.n5 a_10000_15820.n4 0.214786
R5963 a_13360_11960.n0 a_13360_11960.n4 199.935
R5964 a_13360_11960.n0 a_13360_11960.n3 199.53
R5965 a_13360_11960.n0 a_13360_11960.n2 199.53
R5966 a_13360_11960.n0 a_13360_11960.n1 199.53
R5967 a_13360_11960.n5 a_13360_11960.n0 199.53
R5968 a_13360_11960.n0 a_13360_11960.t7 56.2681
R5969 a_13360_11960.n4 a_13360_11960.t4 48.0005
R5970 a_13360_11960.n4 a_13360_11960.t10 48.0005
R5971 a_13360_11960.n3 a_13360_11960.t2 48.0005
R5972 a_13360_11960.n3 a_13360_11960.t1 48.0005
R5973 a_13360_11960.n2 a_13360_11960.t8 48.0005
R5974 a_13360_11960.n2 a_13360_11960.t5 48.0005
R5975 a_13360_11960.n1 a_13360_11960.t3 48.0005
R5976 a_13360_11960.n1 a_13360_11960.t9 48.0005
R5977 a_13360_11960.t0 a_13360_11960.n5 48.0005
R5978 a_13360_11960.n5 a_13360_11960.t6 48.0005
R5979 a_13070_11250.n12 a_13070_11250.t26 363.909
R5980 a_13070_11250.n11 a_13070_11250.t16 351.974
R5981 a_13070_11250.n21 a_13070_11250.n13 299.252
R5982 a_13070_11250.n11 a_13070_11250.n14 299.25
R5983 a_13070_11250.n11 a_13070_11250.n16 299.25
R5984 a_13070_11250.n9 a_13070_11250.t6 242.968
R5985 a_13070_11250.n19 a_13070_11250.n17 200.477
R5986 a_13070_11250.n19 a_13070_11250.n18 199.727
R5987 a_13070_11250.n20 a_13070_11250.t32 194.809
R5988 a_13070_11250.n20 a_13070_11250.t14 194.809
R5989 a_13070_11250.n15 a_13070_11250.t30 194.809
R5990 a_13070_11250.n15 a_13070_11250.t23 194.809
R5991 a_13070_11250.n11 a_13070_11250.n15 163.097
R5992 a_13070_11250.n9 a_13070_11250.n20 161.653
R5993 a_13070_11250.n17 a_13070_11250.t7 48.0005
R5994 a_13070_11250.n17 a_13070_11250.t10 48.0005
R5995 a_13070_11250.n18 a_13070_11250.t8 48.0005
R5996 a_13070_11250.n18 a_13070_11250.t9 48.0005
R5997 a_13070_11250.n14 a_13070_11250.t3 39.4005
R5998 a_13070_11250.n14 a_13070_11250.t0 39.4005
R5999 a_13070_11250.n16 a_13070_11250.t4 39.4005
R6000 a_13070_11250.n16 a_13070_11250.t1 39.4005
R6001 a_13070_11250.t5 a_13070_11250.n21 39.4005
R6002 a_13070_11250.n21 a_13070_11250.t2 39.4005
R6003 a_13070_11250.n12 a_13070_11250.n8 11.6665
R6004 a_13070_11250.n9 a_13070_11250.n19 5.2505
R6005 a_13070_11250.n3 a_13070_11250.t36 4.8248
R6006 a_13070_11250.n10 a_13070_11250.t13 4.5005
R6007 a_13070_11250.n1 a_13070_11250.t34 4.5005
R6008 a_13070_11250.n1 a_13070_11250.t28 4.5005
R6009 a_13070_11250.n0 a_13070_11250.t20 4.5005
R6010 a_13070_11250.n0 a_13070_11250.t24 4.5005
R6011 a_13070_11250.n2 a_13070_11250.t29 4.5005
R6012 a_13070_11250.n2 a_13070_11250.t22 4.5005
R6013 a_13070_11250.n3 a_13070_11250.t25 4.5005
R6014 a_13070_11250.n3 a_13070_11250.t18 4.5005
R6015 a_13070_11250.n10 a_13070_11250.t33 4.5005
R6016 a_13070_11250.n4 a_13070_11250.t27 4.5005
R6017 a_13070_11250.n5 a_13070_11250.t19 4.5005
R6018 a_13070_11250.n5 a_13070_11250.t11 4.5005
R6019 a_13070_11250.n6 a_13070_11250.t15 4.5005
R6020 a_13070_11250.n6 a_13070_11250.t21 4.5005
R6021 a_13070_11250.n7 a_13070_11250.t12 4.5005
R6022 a_13070_11250.n7 a_13070_11250.t17 4.5005
R6023 a_13070_11250.n8 a_13070_11250.t35 4.5005
R6024 a_13070_11250.n8 a_13070_11250.t31 4.5005
R6025 a_13070_11250.n13 a_13070_11250.n9 1.74185
R6026 a_13070_11250.n7 a_13070_11250.n6 0.6585
R6027 a_13070_11250.n6 a_13070_11250.n5 0.6585
R6028 a_13070_11250.n5 a_13070_11250.n4 0.6585
R6029 a_13070_11250.n2 a_13070_11250.n3 0.6585
R6030 a_13070_11250.n0 a_13070_11250.n2 0.6585
R6031 a_13070_11250.n1 a_13070_11250.n0 0.6585
R6032 a_13070_11250.n10 a_13070_11250.n1 0.6585
R6033 a_13070_11250.n8 a_13070_11250.n7 0.6538
R6034 a_13070_11250.n13 a_13070_11250.n11 0.6255
R6035 a_13070_11250.n4 a_13070_11250.n10 0.6115
R6036 a_13070_11250.n13 a_13070_11250.n12 0.34425
R6037 a_20230_3150.n5 a_20230_3150.t2 752.333
R6038 a_20230_3150.n4 a_20230_3150.t1 752.333
R6039 a_20230_3150.n0 a_20230_3150.t6 514.134
R6040 a_20230_3150.n3 a_20230_3150.n2 366.856
R6041 a_20230_3150.t0 a_20230_3150.n5 254.333
R6042 a_20230_3150.n3 a_20230_3150.t4 190.123
R6043 a_20230_3150.n4 a_20230_3150.n3 187.201
R6044 a_20230_3150.n2 a_20230_3150.n1 176.733
R6045 a_20230_3150.n1 a_20230_3150.n0 176.733
R6046 a_20230_3150.n0 a_20230_3150.t3 112.468
R6047 a_20230_3150.n1 a_20230_3150.t5 112.468
R6048 a_20230_3150.n2 a_20230_3150.t7 112.468
R6049 a_20230_3150.n5 a_20230_3150.n4 70.4005
R6050 a_20140_2930.n0 a_20140_2930.t3 750.201
R6051 a_20140_2930.n1 a_20140_2930.t4 349.433
R6052 a_20140_2930.n0 a_20140_2930.t0 276.733
R6053 a_20140_2930.n2 a_20140_2930.n1 206.333
R6054 a_20140_2930.n1 a_20140_2930.n0 48.0005
R6055 a_20140_2930.n2 a_20140_2930.t1 48.0005
R6056 a_20140_2930.t2 a_20140_2930.n2 48.0005
R6057 a_17950_3100.n0 a_17950_3100.t0 713.933
R6058 a_17950_3100.t1 a_17950_3100.n0 337
R6059 a_17950_3100.n0 a_17950_3100.t2 314.233
R6060 a_17540_2930.n2 a_17540_2930.t0 750.201
R6061 a_17540_2930.n1 a_17540_2930.t4 349.433
R6062 a_17540_2930.t1 a_17540_2930.n2 276.733
R6063 a_17540_2930.n1 a_17540_2930.n0 206.333
R6064 a_17540_2930.n0 a_17540_2930.t3 48.0005
R6065 a_17540_2930.n0 a_17540_2930.t2 48.0005
R6066 a_17540_2930.n2 a_17540_2930.n1 48.0005
R6067 a_15320_6670.n0 a_15320_6670.t5 1028.27
R6068 a_15320_6670.n2 a_15320_6670.n1 569.734
R6069 a_15320_6670.n1 a_15320_6670.n0 465.933
R6070 a_15320_6670.n1 a_15320_6670.t3 401.668
R6071 a_15320_6670.n1 a_15320_6670.t4 385.601
R6072 a_15320_6670.n0 a_15320_6670.t2 385.601
R6073 a_15320_6670.t1 a_15320_6670.n2 211.847
R6074 a_15320_6670.n2 a_15320_6670.t0 173.055
R6075 a_12960_8860.n5 a_12960_8860.n4 1269.42
R6076 a_12960_8860.n0 a_12960_8860.n9 299.368
R6077 a_12960_8860.n0 a_12960_8860.n10 299.252
R6078 a_12960_8860.n0 a_12960_8860.n11 299.252
R6079 a_12960_8860.n1 a_12960_8860.n12 299.252
R6080 a_12960_8860.n1 a_12960_8860.n13 299.252
R6081 a_12960_8860.n15 a_12960_8860.n14 299.252
R6082 a_12960_8860.t11 a_12960_8860.n5 275.325
R6083 a_12960_8860.n2 a_12960_8860.t0 238.891
R6084 a_12960_8860.n6 a_12960_8860.t11 178.34
R6085 a_12960_8860.n6 a_12960_8860.t13 178.34
R6086 a_12960_8860.n2 a_12960_8860.t17 161.371
R6087 a_12960_8860.n7 a_12960_8860.n6 152
R6088 a_12960_8860.n4 a_12960_8860.t18 151.792
R6089 a_12960_8860.n5 a_12960_8860.t13 80.3338
R6090 a_12960_8860.n8 a_12960_8860.n2 73.5729
R6091 a_12960_8860.n7 a_12960_8860.n3 68.0438
R6092 a_12960_8860.n4 a_12960_8860.t19 44.2902
R6093 a_12960_8860.n9 a_12960_8860.t1 39.4005
R6094 a_12960_8860.n9 a_12960_8860.t16 39.4005
R6095 a_12960_8860.n10 a_12960_8860.t3 39.4005
R6096 a_12960_8860.n10 a_12960_8860.t6 39.4005
R6097 a_12960_8860.n11 a_12960_8860.t4 39.4005
R6098 a_12960_8860.n11 a_12960_8860.t8 39.4005
R6099 a_12960_8860.n12 a_12960_8860.t5 39.4005
R6100 a_12960_8860.n12 a_12960_8860.t9 39.4005
R6101 a_12960_8860.n13 a_12960_8860.t7 39.4005
R6102 a_12960_8860.n13 a_12960_8860.t2 39.4005
R6103 a_12960_8860.n15 a_12960_8860.t15 39.4005
R6104 a_12960_8860.t10 a_12960_8860.n15 39.4005
R6105 a_12960_8860.n8 a_12960_8860.n7 15.7979
R6106 a_12960_8860.n3 a_12960_8860.t14 15.0005
R6107 a_12960_8860.n3 a_12960_8860.t12 15.0005
R6108 a_12960_8860.n14 a_12960_8860.n8 4.48377
R6109 a_12960_8860.n1 a_12960_8860.n0 0.229667
R6110 a_12960_8860.n14 a_12960_8860.n1 0.229667
R6111 a_16000_6670.t5 a_16000_6670.t3 377.567
R6112 a_16000_6670.n2 a_16000_6670.n1 237.353
R6113 a_16000_6670.t1 a_16000_6670.n3 229.127
R6114 a_16000_6670.n0 a_16000_6670.t4 220.505
R6115 a_16000_6670.n1 a_16000_6670.n0 196.817
R6116 a_16000_6670.n3 a_16000_6670.t0 158.335
R6117 a_16000_6670.n2 a_16000_6670.t2 151.935
R6118 a_16000_6670.n3 a_16000_6670.n2 121.6
R6119 a_16000_6670.t3 a_16000_6670.n0 92.3838
R6120 a_16000_6670.n1 a_16000_6670.t5 92.3838
R6121 pll_bgr_magic_3_0.VV1 pll_bgr_magic_3_0.VV1.n6 1052.95
R6122 pll_bgr_magic_3_0.VV1.n2 pll_bgr_magic_3_0.VV1.n0 297.988
R6123 pll_bgr_magic_3_0.VV1.n3 pll_bgr_magic_3_0.VV1.n2 264.61
R6124 pll_bgr_magic_3_0.VV1.n3 pll_bgr_magic_3_0.VV1.t6 208.868
R6125 pll_bgr_magic_3_0.VV1.n4 pll_bgr_magic_3_0.VV1.t7 208.868
R6126 pll_bgr_magic_3_0.VV1.n5 pll_bgr_magic_3_0.VV1.t8 208.868
R6127 pll_bgr_magic_3_0.VV1.n6 pll_bgr_magic_3_0.VV1.t5 208.868
R6128 pll_bgr_magic_3_0.VV1.n6 pll_bgr_magic_3_0.VV1.n5 208.868
R6129 pll_bgr_magic_3_0.VV1.n5 pll_bgr_magic_3_0.VV1.n4 208.868
R6130 pll_bgr_magic_3_0.VV1.n4 pll_bgr_magic_3_0.VV1.n3 208.868
R6131 pll_bgr_magic_3_0.VV1.n2 pll_bgr_magic_3_0.VV1.n1 195.035
R6132 pll_bgr_magic_3_0.VV1.n1 pll_bgr_magic_3_0.VV1.t1 60.0005
R6133 pll_bgr_magic_3_0.VV1.n1 pll_bgr_magic_3_0.VV1.t2 60.0005
R6134 pll_bgr_magic_3_0.VV1 pll_bgr_magic_3_0.VV1.t3 59.81
R6135 pll_bgr_magic_3_0.VV1.n0 pll_bgr_magic_3_0.VV1.t4 49.2505
R6136 pll_bgr_magic_3_0.VV1.n0 pll_bgr_magic_3_0.VV1.t0 49.2505
R6137 a_15870_5490.n2 a_15870_5490.n1 424.447
R6138 a_15870_5490.n2 a_15870_5490.n0 354.046
R6139 a_15870_5490.n14 a_15870_5490.n13 313
R6140 a_15870_5490.n6 a_15870_5490.t13 297.233
R6141 a_15870_5490.n7 a_15870_5490.t13 297.233
R6142 a_15870_5490.t15 a_15870_5490.n4 297.233
R6143 a_15870_5490.n5 a_15870_5490.t15 297.233
R6144 a_15870_5490.n9 a_15870_5490.t4 281.596
R6145 a_15870_5490.n15 a_15870_5490.n14 242.601
R6146 a_15870_5490.n3 a_15870_5490.n2 220.8
R6147 a_15870_5490.n14 a_15870_5490.n12 220.8
R6148 a_15870_5490.n6 a_15870_5490.n5 216.9
R6149 a_15870_5490.n10 a_15870_5490.n8 167.644
R6150 a_15870_5490.n9 a_15870_5490.t1 118.666
R6151 a_15870_5490.n8 a_15870_5490.n7 81.6727
R6152 a_15870_5490.n8 a_15870_5490.n4 81.6727
R6153 a_15870_5490.n7 a_15870_5490.t11 80.3338
R6154 a_15870_5490.t11 a_15870_5490.n6 80.3338
R6155 a_15870_5490.t10 a_15870_5490.n4 80.3338
R6156 a_15870_5490.n5 a_15870_5490.t10 80.3338
R6157 a_15870_5490.n12 a_15870_5490.t12 70.0829
R6158 a_15870_5490.n11 a_15870_5490.n3 64.0005
R6159 a_15870_5490.n12 a_15870_5490.n11 64.0005
R6160 a_15870_5490.n3 a_15870_5490.t14 63.6829
R6161 a_15870_5490.n10 a_15870_5490.n9 60.4288
R6162 a_15870_5490.n13 a_15870_5490.t6 60.0005
R6163 a_15870_5490.n13 a_15870_5490.t7 60.0005
R6164 a_15870_5490.t8 a_15870_5490.n15 60.0005
R6165 a_15870_5490.n15 a_15870_5490.t5 60.0005
R6166 a_15870_5490.n11 a_15870_5490.n10 52.113
R6167 a_15870_5490.n0 a_15870_5490.t2 49.2505
R6168 a_15870_5490.n0 a_15870_5490.t0 49.2505
R6169 a_15870_5490.n1 a_15870_5490.t3 49.2505
R6170 a_15870_5490.n1 a_15870_5490.t9 49.2505
R6171 a_12760_5460.n0 a_12760_5460.t3 517.347
R6172 a_12760_5460.n2 a_12760_5460.n0 417.574
R6173 a_12760_5460.n2 a_12760_5460.n1 244.716
R6174 a_12760_5460.n0 a_12760_5460.t4 228.148
R6175 a_12760_5460.t0 a_12760_5460.n2 221.411
R6176 a_12760_5460.n1 a_12760_5460.t2 24.0005
R6177 a_12760_5460.n1 a_12760_5460.t1 24.0005
R6178 a_12680_5910.t0 a_12680_5910.t1 39.4005
R6179 a_12380_5460.n4 a_12380_5460.n0 1319.38
R6180 a_12380_5460.n0 a_12380_5460.t3 562.333
R6181 a_12380_5460.n2 a_12380_5460.t5 388.813
R6182 a_12380_5460.n2 a_12380_5460.t6 356.68
R6183 a_12380_5460.n3 a_12380_5460.n2 232
R6184 a_12380_5460.n0 a_12380_5460.t4 224.934
R6185 a_12380_5460.t0 a_12380_5460.n4 221.411
R6186 a_12380_5460.n3 a_12380_5460.n1 157.278
R6187 a_12380_5460.n4 a_12380_5460.n3 90.64
R6188 a_12380_5460.n1 a_12380_5460.t1 24.0005
R6189 a_12380_5460.n1 a_12380_5460.t2 24.0005
R6190 a_11040_2860.n4 a_11040_2860.t0 777.4
R6191 a_11040_2860.t8 a_11040_2860.t10 514.134
R6192 a_11040_2860.n3 a_11040_2860.n2 364.178
R6193 a_11040_2860.n0 a_11040_2860.t3 353.467
R6194 a_11040_2860.t5 a_11040_2860.n5 353.467
R6195 a_11040_2860.n6 a_11040_2860.t5 318.702
R6196 a_11040_2860.n6 a_11040_2860.t8 307.909
R6197 a_11040_2860.n5 a_11040_2860.t11 289.2
R6198 a_11040_2860.n4 a_11040_2860.n3 257.079
R6199 a_11040_2860.t1 a_11040_2860.n7 233
R6200 a_11040_2860.n0 a_11040_2860.t9 192.8
R6201 a_11040_2860.n2 a_11040_2860.n1 176.733
R6202 a_11040_2860.n1 a_11040_2860.t2 112.468
R6203 a_11040_2860.n2 a_11040_2860.t7 112.468
R6204 a_11040_2860.n3 a_11040_2860.t4 112.468
R6205 a_11040_2860.n5 a_11040_2860.t6 112.468
R6206 a_11040_2860.n1 a_11040_2860.n0 96.4005
R6207 a_11040_2860.n7 a_11040_2860.n6 38.2642
R6208 a_11040_2860.n7 a_11040_2860.n4 21.3338
R6209 a_10910_3020.n0 a_10910_3020.t3 761.4
R6210 a_10910_3020.n1 a_10910_3020.t4 349.433
R6211 a_10910_3020.n0 a_10910_3020.t1 254.333
R6212 a_10910_3020.n2 a_10910_3020.n1 206.333
R6213 a_10910_3020.n1 a_10910_3020.n0 70.4005
R6214 a_10910_3020.t2 a_10910_3020.n2 48.0005
R6215 a_10910_3020.n2 a_10910_3020.t0 48.0005
R6216 a_16240_3020.n0 a_16240_3020.t1 721.4
R6217 a_16240_3020.n1 a_16240_3020.t4 350.349
R6218 a_16240_3020.n0 a_16240_3020.t2 276.733
R6219 a_16240_3020.n2 a_16240_3020.n1 206.333
R6220 a_16240_3020.n1 a_16240_3020.n0 48.0005
R6221 a_16240_3020.t0 a_16240_3020.n2 48.0005
R6222 a_16240_3020.n2 a_16240_3020.t3 48.0005
R6223 a_15820_2860.n1 a_15820_2860.n0 701.467
R6224 a_15820_2860.n1 a_15820_2860.t1 694.201
R6225 a_15820_2860.n0 a_15820_2860.t2 321.334
R6226 a_15820_2860.t0 a_15820_2860.n1 314.921
R6227 a_15820_2860.n0 a_15820_2860.t3 144.601
R6228 a_17630_3150.n4 a_17630_3150.t0 752.333
R6229 a_17630_3150.t1 a_17630_3150.n5 752.333
R6230 a_17630_3150.n0 a_17630_3150.t7 514.134
R6231 a_17630_3150.n3 a_17630_3150.n2 366.856
R6232 a_17630_3150.n5 a_17630_3150.t2 254.333
R6233 a_17630_3150.n3 a_17630_3150.t5 190.123
R6234 a_17630_3150.n4 a_17630_3150.n3 187.201
R6235 a_17630_3150.n2 a_17630_3150.n1 176.733
R6236 a_17630_3150.n1 a_17630_3150.n0 176.733
R6237 a_17630_3150.n0 a_17630_3150.t4 112.468
R6238 a_17630_3150.n1 a_17630_3150.t6 112.468
R6239 a_17630_3150.n2 a_17630_3150.t3 112.468
R6240 a_17630_3150.n5 a_17630_3150.n4 70.4005
R6241 a_11960_2860.n0 a_11960_2860.t3 723.534
R6242 a_11960_2860.n1 a_11960_2860.t4 553.534
R6243 a_11960_2860.n0 a_11960_2860.t1 254.333
R6244 a_11960_2860.n2 a_11960_2860.n1 206.333
R6245 a_11960_2860.n1 a_11960_2860.n0 70.4005
R6246 a_11960_2860.t2 a_11960_2860.n2 48.0005
R6247 a_11960_2860.n2 a_11960_2860.t0 48.0005
R6248 a_18390_5940.n3 a_18390_5940.t9 377.567
R6249 a_18390_5940.n2 a_18390_5940.t7 297.233
R6250 a_18390_5940.n4 a_18390_5940.n2 231.575
R6251 a_18390_5940.n4 a_18390_5940.n3 228.778
R6252 a_18390_5940.n3 a_18390_5940.t6 216.9
R6253 a_18390_5940.n0 a_18390_5940.n5 153.401
R6254 a_18390_5940.n6 a_18390_5940.n0 153.4
R6255 a_18390_5940.n2 a_18390_5940.t8 136.567
R6256 a_18390_5940.n0 a_18390_5940.n1 54.9641
R6257 a_18390_5940.n5 a_18390_5940.t2 24.6255
R6258 a_18390_5940.n5 a_18390_5940.t1 24.6255
R6259 a_18390_5940.n6 a_18390_5940.t0 24.6255
R6260 a_18390_5940.t3 a_18390_5940.n6 24.6255
R6261 a_18390_5940.n0 a_18390_5940.n4 22.2974
R6262 a_18390_5940.n1 a_18390_5940.t5 15.0005
R6263 a_18390_5940.n1 a_18390_5940.t4 15.0005
R6264 a_15790_17280.t20 a_15790_17280.t0 130.1
R6265 a_15790_17280.t1 a_15790_17280.t4 0.1603
R6266 a_15790_17280.t15 a_15790_17280.t1 0.1603
R6267 a_15790_17280.t18 a_15790_17280.t15 0.1603
R6268 a_15790_17280.t11 a_15790_17280.t18 0.1603
R6269 a_15790_17280.t16 a_15790_17280.t11 0.1603
R6270 a_15790_17280.t19 a_15790_17280.t16 0.1603
R6271 a_15790_17280.t13 a_15790_17280.t19 0.1603
R6272 a_15790_17280.t7 a_15790_17280.t13 0.1603
R6273 a_15790_17280.t6 a_15790_17280.t2 0.1603
R6274 a_15790_17280.t12 a_15790_17280.t6 0.1603
R6275 a_15790_17280.t9 a_15790_17280.t12 0.1603
R6276 a_15790_17280.t5 a_15790_17280.t9 0.1603
R6277 a_15790_17280.t10 a_15790_17280.t5 0.1603
R6278 a_15790_17280.t8 a_15790_17280.t10 0.1603
R6279 a_15790_17280.t14 a_15790_17280.t8 0.1603
R6280 a_15790_17280.t0 a_15790_17280.t14 0.1603
R6281 a_15790_17280.t17 a_15790_17280.n0 0.159278
R6282 a_15790_17280.t2 a_15790_17280.t17 0.137822
R6283 a_15790_17280.n0 a_15790_17280.t7 0.1368
R6284 a_15790_17280.n0 a_15790_17280.t3 0.00152174
R6285 a_10160_10990.n15 a_10160_10990.t22 310.488
R6286 a_10160_10990.n9 a_10160_10990.t17 310.488
R6287 a_10160_10990.n0 a_10160_10990.t18 310.488
R6288 a_10160_10990.n13 a_10160_10990.n12 297.433
R6289 a_10160_10990.n4 a_10160_10990.n3 297.433
R6290 a_10160_10990.n19 a_10160_10990.n18 297.433
R6291 a_10160_10990.n7 a_10160_10990.t3 248.133
R6292 a_10160_10990.n7 a_10160_10990.n6 199.383
R6293 a_10160_10990.n8 a_10160_10990.n5 194.883
R6294 a_10160_10990.n17 a_10160_10990.t7 184.097
R6295 a_10160_10990.n11 a_10160_10990.t9 184.097
R6296 a_10160_10990.n2 a_10160_10990.t5 184.097
R6297 a_10160_10990.n16 a_10160_10990.n15 167.094
R6298 a_10160_10990.n10 a_10160_10990.n9 167.094
R6299 a_10160_10990.n1 a_10160_10990.n0 167.094
R6300 a_10160_10990.n18 a_10160_10990.n17 161.3
R6301 a_10160_10990.n13 a_10160_10990.n11 161.3
R6302 a_10160_10990.n4 a_10160_10990.n2 161.3
R6303 a_10160_10990.n15 a_10160_10990.t19 120.501
R6304 a_10160_10990.n16 a_10160_10990.t15 120.501
R6305 a_10160_10990.n9 a_10160_10990.t20 120.501
R6306 a_10160_10990.n10 a_10160_10990.t11 120.501
R6307 a_10160_10990.n0 a_10160_10990.t21 120.501
R6308 a_10160_10990.n1 a_10160_10990.t13 120.501
R6309 a_10160_10990.n6 a_10160_10990.t4 48.0005
R6310 a_10160_10990.n6 a_10160_10990.t1 48.0005
R6311 a_10160_10990.n5 a_10160_10990.t0 48.0005
R6312 a_10160_10990.n5 a_10160_10990.t2 48.0005
R6313 a_10160_10990.n17 a_10160_10990.n16 40.7027
R6314 a_10160_10990.n11 a_10160_10990.n10 40.7027
R6315 a_10160_10990.n2 a_10160_10990.n1 40.7027
R6316 a_10160_10990.n12 a_10160_10990.t12 39.4005
R6317 a_10160_10990.n12 a_10160_10990.t10 39.4005
R6318 a_10160_10990.n3 a_10160_10990.t14 39.4005
R6319 a_10160_10990.n3 a_10160_10990.t6 39.4005
R6320 a_10160_10990.t16 a_10160_10990.n19 39.4005
R6321 a_10160_10990.n19 a_10160_10990.t8 39.4005
R6322 a_10160_10990.n14 a_10160_10990.n4 6.6255
R6323 a_10160_10990.n18 a_10160_10990.n14 6.6255
R6324 a_10160_10990.n8 a_10160_10990.n7 5.2505
R6325 a_10160_10990.n14 a_10160_10990.n13 4.5005
R6326 a_10160_10990.n13 a_10160_10990.n8 0.78175
R6327 a_10030_11260.n14 a_10030_11260.t18 362.341
R6328 a_10030_11260.n11 a_10030_11260.t17 355.094
R6329 a_10030_11260.n16 a_10030_11260.n15 302.183
R6330 a_10030_11260.n11 a_10030_11260.n10 302.183
R6331 a_10030_11260.n25 a_10030_11260.n24 302.183
R6332 a_10030_11260.n20 a_10030_11260.t9 242.968
R6333 a_10030_11260.n19 a_10030_11260.n17 200.477
R6334 a_10030_11260.n19 a_10030_11260.n18 199.727
R6335 a_10030_11260.n21 a_10030_11260.t27 194.809
R6336 a_10030_11260.n21 a_10030_11260.t13 194.809
R6337 a_10030_11260.n12 a_10030_11260.t21 194.809
R6338 a_10030_11260.n12 a_10030_11260.t32 194.809
R6339 a_10030_11260.n13 a_10030_11260.n12 166.03
R6340 a_10030_11260.n22 a_10030_11260.n21 161.53
R6341 a_10030_11260.n18 a_10030_11260.t2 48.0005
R6342 a_10030_11260.n18 a_10030_11260.t1 48.0005
R6343 a_10030_11260.n17 a_10030_11260.t0 48.0005
R6344 a_10030_11260.n17 a_10030_11260.t10 48.0005
R6345 a_10030_11260.n14 a_10030_11260.n8 40.0796
R6346 a_10030_11260.n15 a_10030_11260.t7 39.4005
R6347 a_10030_11260.n15 a_10030_11260.t4 39.4005
R6348 a_10030_11260.n10 a_10030_11260.t3 39.4005
R6349 a_10030_11260.n10 a_10030_11260.t6 39.4005
R6350 a_10030_11260.t8 a_10030_11260.n25 39.4005
R6351 a_10030_11260.n25 a_10030_11260.t5 39.4005
R6352 a_10030_11260.n20 a_10030_11260.n19 5.2505
R6353 a_10030_11260.n3 a_10030_11260.t24 4.8248
R6354 a_10030_11260.n9 a_10030_11260.t28 4.5005
R6355 a_10030_11260.n1 a_10030_11260.t22 4.5005
R6356 a_10030_11260.n1 a_10030_11260.t15 4.5005
R6357 a_10030_11260.n0 a_10030_11260.t34 4.5005
R6358 a_10030_11260.n0 a_10030_11260.t11 4.5005
R6359 a_10030_11260.n2 a_10030_11260.t16 4.5005
R6360 a_10030_11260.n2 a_10030_11260.t36 4.5005
R6361 a_10030_11260.n3 a_10030_11260.t12 4.5005
R6362 a_10030_11260.n3 a_10030_11260.t31 4.5005
R6363 a_10030_11260.n9 a_10030_11260.t20 4.5005
R6364 a_10030_11260.n4 a_10030_11260.t14 4.5005
R6365 a_10030_11260.n5 a_10030_11260.t33 4.5005
R6366 a_10030_11260.n5 a_10030_11260.t25 4.5005
R6367 a_10030_11260.n6 a_10030_11260.t29 4.5005
R6368 a_10030_11260.n6 a_10030_11260.t35 4.5005
R6369 a_10030_11260.n7 a_10030_11260.t26 4.5005
R6370 a_10030_11260.n7 a_10030_11260.t30 4.5005
R6371 a_10030_11260.n8 a_10030_11260.t23 4.5005
R6372 a_10030_11260.n8 a_10030_11260.t19 4.5005
R6373 a_10030_11260.n23 a_10030_11260.n22 4.5005
R6374 a_10030_11260.n16 a_10030_11260.n14 2.90725
R6375 a_10030_11260.n13 a_10030_11260.n11 0.7505
R6376 a_10030_11260.n24 a_10030_11260.n23 0.7505
R6377 a_10030_11260.n7 a_10030_11260.n6 0.6585
R6378 a_10030_11260.n6 a_10030_11260.n5 0.6585
R6379 a_10030_11260.n5 a_10030_11260.n4 0.6585
R6380 a_10030_11260.n2 a_10030_11260.n3 0.6585
R6381 a_10030_11260.n0 a_10030_11260.n2 0.6585
R6382 a_10030_11260.n1 a_10030_11260.n0 0.6585
R6383 a_10030_11260.n9 a_10030_11260.n1 0.6585
R6384 a_10030_11260.n8 a_10030_11260.n7 0.6538
R6385 a_10030_11260.n4 a_10030_11260.n9 0.6115
R6386 a_10030_11260.n22 a_10030_11260.n20 0.422375
R6387 a_10030_11260.n24 a_10030_11260.n13 0.3755
R6388 a_10030_11260.n23 a_10030_11260.n16 0.3755
R6389 a_10751_12090.n2 a_10751_12090.n0 302.507
R6390 a_10751_12090.n10 a_10751_12090.n9 302.163
R6391 a_10751_12090.n8 a_10751_12090.n7 302.163
R6392 a_10751_12090.n6 a_10751_12090.n5 302.163
R6393 a_10751_12090.n4 a_10751_12090.n3 302.163
R6394 a_10751_12090.n2 a_10751_12090.n1 302.163
R6395 a_10751_12090.n11 a_10751_12090.t14 291.502
R6396 a_10751_12090.n14 a_10751_12090.t15 291.288
R6397 a_10751_12090.n13 a_10751_12090.t16 291.288
R6398 a_10751_12090.n12 a_10751_12090.t13 291.288
R6399 a_10751_12090.n11 a_10751_12090.t17 291.288
R6400 a_10751_12090.t0 a_10751_12090.n15 133.005
R6401 a_10751_12090.n9 a_10751_12090.t1 39.4005
R6402 a_10751_12090.n9 a_10751_12090.t12 39.4005
R6403 a_10751_12090.n7 a_10751_12090.t3 39.4005
R6404 a_10751_12090.n7 a_10751_12090.t7 39.4005
R6405 a_10751_12090.n5 a_10751_12090.t4 39.4005
R6406 a_10751_12090.n5 a_10751_12090.t8 39.4005
R6407 a_10751_12090.n3 a_10751_12090.t6 39.4005
R6408 a_10751_12090.n3 a_10751_12090.t9 39.4005
R6409 a_10751_12090.n1 a_10751_12090.t5 39.4005
R6410 a_10751_12090.n1 a_10751_12090.t2 39.4005
R6411 a_10751_12090.n0 a_10751_12090.t11 39.4005
R6412 a_10751_12090.n0 a_10751_12090.t10 39.4005
R6413 a_10751_12090.n15 a_10751_12090.n10 12.0474
R6414 a_10751_12090.n15 a_10751_12090.n14 6.4005
R6415 a_10751_12090.n12 a_10751_12090.n11 0.643357
R6416 a_10751_12090.n14 a_10751_12090.n13 0.643357
R6417 a_10751_12090.n4 a_10751_12090.n2 0.34425
R6418 a_10751_12090.n6 a_10751_12090.n4 0.34425
R6419 a_10751_12090.n8 a_10751_12090.n6 0.34425
R6420 a_10751_12090.n10 a_10751_12090.n8 0.34425
R6421 a_10751_12090.n13 a_10751_12090.n12 0.214786
R6422 a_20550_3100.n0 a_20550_3100.t0 713.933
R6423 a_20550_3100.t1 a_20550_3100.n0 337
R6424 a_20550_3100.n0 a_20550_3100.t2 314.233
R6425 a_20850_2800.t0 a_20850_2800.t1 96.0005
R6426 a_19630_3180.t2 a_19630_3180.t4 1012.2
R6427 a_19630_3180.n0 a_19630_3180.t0 663.801
R6428 a_19630_3180.n2 a_19630_3180.n1 431.401
R6429 a_19630_3180.t3 a_19630_3180.t5 401.668
R6430 a_19630_3180.n0 a_19630_3180.t2 361.692
R6431 a_19630_3180.n1 a_19630_3180.t6 353.467
R6432 a_19630_3180.t1 a_19630_3180.n2 298.921
R6433 a_19630_3180.n1 a_19630_3180.t3 257.067
R6434 a_19630_3180.n2 a_19630_3180.n0 67.2005
R6435 a_14930_5490.n0 a_14930_5490.t2 441.834
R6436 a_14930_5490.n0 a_14930_5490.t3 313.3
R6437 a_14930_5490.n1 a_14930_5490.n0 235.201
R6438 a_14930_5490.t0 a_14930_5490.n1 219.528
R6439 a_14930_5490.n1 a_14930_5490.t1 167.935
R6440 a_15320_5490.n0 a_15320_5490.t4 1205
R6441 a_15320_5490.n2 a_15320_5490.t3 522.168
R6442 a_15320_5490.n1 a_15320_5490.n0 441.834
R6443 a_15320_5490.n3 a_15320_5490.n2 235.201
R6444 a_15320_5490.t0 a_15320_5490.n3 229.127
R6445 a_15320_5490.n1 a_15320_5490.t5 217.905
R6446 a_15320_5490.n0 a_15320_5490.t2 208.868
R6447 a_15320_5490.n3 a_15320_5490.t1 158.335
R6448 a_15320_5490.n2 a_15320_5490.n1 15.063
R6449 a_12760_6640.n0 a_12760_6640.t3 517.347
R6450 a_12760_6640.n2 a_12760_6640.n0 417.574
R6451 a_12760_6640.n2 a_12760_6640.n1 244.716
R6452 a_12760_6640.n0 a_12760_6640.t4 228.148
R6453 a_12760_6640.t1 a_12760_6640.n2 221.411
R6454 a_12760_6640.n1 a_12760_6640.t0 24.0005
R6455 a_12760_6640.n1 a_12760_6640.t2 24.0005
R6456 a_12680_6670.t0 a_12680_6670.t1 39.4005
R6457 a_12380_6640.n4 a_12380_6640.n0 1319.38
R6458 a_12380_6640.n0 a_12380_6640.t3 562.333
R6459 a_12380_6640.n2 a_12380_6640.t5 388.813
R6460 a_12380_6640.n2 a_12380_6640.t4 356.68
R6461 a_12380_6640.n3 a_12380_6640.n2 232
R6462 a_12380_6640.n0 a_12380_6640.t6 224.934
R6463 a_12380_6640.t0 a_12380_6640.n4 221.411
R6464 a_12380_6640.n3 a_12380_6640.n1 157.278
R6465 a_12380_6640.n4 a_12380_6640.n3 90.64
R6466 a_12380_6640.n1 a_12380_6640.t1 24.0005
R6467 a_12380_6640.n1 a_12380_6640.t2 24.0005
R6468 a_12700_3340.n0 a_12700_3340.t1 723
R6469 a_12700_3340.t3 a_12700_3340.t2 514.134
R6470 a_12700_3340.n0 a_12700_3340.t3 335.983
R6471 a_12700_3340.t0 a_12700_3340.n0 314.921
R6472 a_12540_2890.n0 a_12540_2890.t1 531.067
R6473 a_12540_2890.t0 a_12540_2890.n0 48.0005
R6474 a_12540_2890.n0 a_12540_2890.t2 48.0005
R6475 a_10060_12570.n1 a_10060_12570.n2 199.935
R6476 a_10060_12570.n0 a_10060_12570.n4 199.53
R6477 a_10060_12570.n0 a_10060_12570.n5 199.53
R6478 a_10060_12570.n1 a_10060_12570.n3 199.53
R6479 a_10060_12570.n6 a_10060_12570.n1 199.53
R6480 a_10060_12570.n0 a_10060_12570.t10 97.8998
R6481 a_10060_12570.n4 a_10060_12570.t5 48.0005
R6482 a_10060_12570.n4 a_10060_12570.t2 48.0005
R6483 a_10060_12570.n5 a_10060_12570.t1 48.0005
R6484 a_10060_12570.n5 a_10060_12570.t8 48.0005
R6485 a_10060_12570.n3 a_10060_12570.t0 48.0005
R6486 a_10060_12570.n3 a_10060_12570.t9 48.0005
R6487 a_10060_12570.n2 a_10060_12570.t6 48.0005
R6488 a_10060_12570.n2 a_10060_12570.t3 48.0005
R6489 a_10060_12570.n6 a_10060_12570.t7 48.0005
R6490 a_10060_12570.t4 a_10060_12570.n6 48.0005
R6491 a_10060_12570.n1 a_10060_12570.n0 1.09425
R6492 a_14010_6640.t1 a_14010_6640.n2 500.086
R6493 a_14010_6640.n1 a_14010_6640.n0 473.334
R6494 a_14010_6640.n0 a_14010_6640.t2 465.933
R6495 a_14010_6640.t1 a_14010_6640.n2 461.389
R6496 a_14010_6640.n0 a_14010_6640.t3 321.334
R6497 a_14010_6640.n1 a_14010_6640.t0 177.577
R6498 a_14010_6640.n2 a_14010_6640.n1 48.3899
R6499 a_13680_6640.t0 a_13680_6640.n2 500.086
R6500 a_13680_6640.n1 a_13680_6640.n0 473.334
R6501 a_13680_6640.n0 a_13680_6640.t3 465.933
R6502 a_13680_6640.t0 a_13680_6640.n2 461.389
R6503 a_13680_6640.n0 a_13680_6640.t2 321.334
R6504 a_13680_6640.n1 a_13680_6640.t1 177.577
R6505 a_13680_6640.n2 a_13680_6640.n1 48.3899
R6506 a_13200_5910.t0 a_13200_5910.t1 39.4005
R6507 a_19530_10890.n1 a_19530_10890.t6 401.668
R6508 a_19530_10890.n5 a_19530_10890.n4 297.394
R6509 a_19530_10890.n3 a_19530_10890.t2 252.248
R6510 a_19530_10890.n2 a_19530_10890.n1 208.868
R6511 a_19530_10890.n4 a_19530_10890.n0 195.582
R6512 a_19530_10890.n1 a_19530_10890.t7 192.8
R6513 a_19530_10890.n2 a_19530_10890.t0 192.8
R6514 a_19530_10890.n4 a_19530_10890.n3 161.3
R6515 a_19530_10890.n0 a_19530_10890.t5 60.0005
R6516 a_19530_10890.n0 a_19530_10890.t4 60.0005
R6517 a_19530_10890.n3 a_19530_10890.n2 59.4472
R6518 a_19530_10890.n5 a_19530_10890.t1 49.2505
R6519 a_19530_10890.t3 a_19530_10890.n5 49.2505
R6520 a_18510_9670.n7 a_18510_9670.n5 482.582
R6521 a_18510_9670.n3 a_18510_9670.t8 304.634
R6522 a_18510_9670.n0 a_18510_9670.t11 304.634
R6523 a_18510_9670.n3 a_18510_9670.t10 279.134
R6524 a_18510_9670.t12 a_18510_9670.n0 277
R6525 a_18510_9670.n8 a_18510_9670.n1 204.201
R6526 a_18510_9670.n4 a_18510_9670.n2 204.201
R6527 a_18510_9670.n10 a_18510_9670.n9 204.201
R6528 a_18510_9670.n7 a_18510_9670.n6 120.981
R6529 a_18510_9670.n8 a_18510_9670.n4 74.6672
R6530 a_18510_9670.n9 a_18510_9670.n8 74.6672
R6531 a_18510_9670.n1 a_18510_9670.t3 60.0005
R6532 a_18510_9670.n1 a_18510_9670.t7 60.0005
R6533 a_18510_9670.n2 a_18510_9670.t6 60.0005
R6534 a_18510_9670.n2 a_18510_9670.t9 60.0005
R6535 a_18510_9670.t12 a_18510_9670.n10 60.0005
R6536 a_18510_9670.n10 a_18510_9670.t2 60.0005
R6537 a_18510_9670.n8 a_18510_9670.n7 28.5443
R6538 a_18510_9670.n5 a_18510_9670.t5 24.0005
R6539 a_18510_9670.n5 a_18510_9670.t4 24.0005
R6540 a_18510_9670.n6 a_18510_9670.t0 24.0005
R6541 a_18510_9670.n6 a_18510_9670.t1 24.0005
R6542 a_18510_9670.n4 a_18510_9670.n3 16.0005
R6543 a_18510_9670.n9 a_18510_9670.n0 16.0005
R6544 a_10900_14480.t0 a_10900_14480.n129 172.969
R6545 a_10900_14480.n119 a_10900_14480.n118 83.5719
R6546 a_10900_14480.n121 a_10900_14480.n120 83.5719
R6547 a_10900_14480.n123 a_10900_14480.n122 83.5719
R6548 a_10900_14480.n109 a_10900_14480.n108 83.5719
R6549 a_10900_14480.n101 a_10900_14480.n11 83.5719
R6550 a_10900_14480.n94 a_10900_14480.n12 83.5719
R6551 a_10900_14480.n96 a_10900_14480.n95 83.5719
R6552 a_10900_14480.n88 a_10900_14480.n16 83.5719
R6553 a_10900_14480.n83 a_10900_14480.n17 83.5719
R6554 a_10900_14480.n75 a_10900_14480.n74 83.5719
R6555 a_10900_14480.n73 a_10900_14480.n72 83.5719
R6556 a_10900_14480.n71 a_10900_14480.n70 83.5719
R6557 a_10900_14480.n41 a_10900_14480.n40 83.5719
R6558 a_10900_14480.n48 a_10900_14480.n47 83.5719
R6559 a_10900_14480.n34 a_10900_14480.n31 83.5719
R6560 a_10900_14480.n53 a_10900_14480.n30 83.5719
R6561 a_10900_14480.n60 a_10900_14480.n59 83.5719
R6562 a_10900_14480.n28 a_10900_14480.n26 83.5719
R6563 a_10900_14480.n119 a_10900_14480.n117 73.3165
R6564 a_10900_14480.n103 a_10900_14480.n11 73.3165
R6565 a_10900_14480.n90 a_10900_14480.n16 73.3165
R6566 a_10900_14480.n76 a_10900_14480.n75 73.3165
R6567 a_10900_14480.n47 a_10900_14480.n46 73.3165
R6568 a_10900_14480.n59 a_10900_14480.n58 73.3165
R6569 a_10900_14480.n122 a_10900_14480.n6 73.19
R6570 a_10900_14480.n108 a_10900_14480.n107 73.19
R6571 a_10900_14480.n95 a_10900_14480.n93 73.19
R6572 a_10900_14480.n71 a_10900_14480.n23 73.19
R6573 a_10900_14480.n40 a_10900_14480.n35 73.19
R6574 a_10900_14480.n55 a_10900_14480.n30 73.19
R6575 a_10900_14480.n84 a_10900_14480.t4 65.0299
R6576 a_10900_14480.t2 a_10900_14480.n24 65.0299
R6577 a_10900_14480.n111 a_10900_14480.t1 36.6639
R6578 a_10900_14480.t6 a_10900_14480.n39 36.6639
R6579 a_10900_14480.n121 a_10900_14480.n119 26.074
R6580 a_10900_14480.n94 a_10900_14480.n11 26.074
R6581 a_10900_14480.n83 a_10900_14480.n16 26.074
R6582 a_10900_14480.n75 a_10900_14480.n73 26.074
R6583 a_10900_14480.n47 a_10900_14480.n34 26.074
R6584 a_10900_14480.n59 a_10900_14480.n28 26.074
R6585 a_10900_14480.n122 a_10900_14480.t7 25.7843
R6586 a_10900_14480.n108 a_10900_14480.t1 25.7843
R6587 a_10900_14480.n95 a_10900_14480.t8 25.7843
R6588 a_10900_14480.t3 a_10900_14480.n71 25.7843
R6589 a_10900_14480.n40 a_10900_14480.t6 25.7843
R6590 a_10900_14480.t5 a_10900_14480.n30 25.7843
R6591 a_10900_14480.n77 a_10900_14480.n65 9.3005
R6592 a_10900_14480.n65 a_10900_14480.n21 9.3005
R6593 a_10900_14480.n65 a_10900_14480.n22 9.3005
R6594 a_10900_14480.n81 a_10900_14480.n65 9.3005
R6595 a_10900_14480.n67 a_10900_14480.n21 9.3005
R6596 a_10900_14480.n67 a_10900_14480.n22 9.3005
R6597 a_10900_14480.n67 a_10900_14480.n19 9.3005
R6598 a_10900_14480.n81 a_10900_14480.n67 9.3005
R6599 a_10900_14480.n82 a_10900_14480.n21 9.3005
R6600 a_10900_14480.n82 a_10900_14480.n20 9.3005
R6601 a_10900_14480.n82 a_10900_14480.n22 9.3005
R6602 a_10900_14480.n82 a_10900_14480.n19 9.3005
R6603 a_10900_14480.n82 a_10900_14480.n81 9.3005
R6604 a_10900_14480.n81 a_10900_14480.n69 9.3005
R6605 a_10900_14480.n69 a_10900_14480.n19 9.3005
R6606 a_10900_14480.n69 a_10900_14480.n22 9.3005
R6607 a_10900_14480.n69 a_10900_14480.n20 9.3005
R6608 a_10900_14480.n81 a_10900_14480.n64 9.3005
R6609 a_10900_14480.n64 a_10900_14480.n19 9.3005
R6610 a_10900_14480.n64 a_10900_14480.n22 9.3005
R6611 a_10900_14480.n64 a_10900_14480.n20 9.3005
R6612 a_10900_14480.n77 a_10900_14480.n64 9.3005
R6613 a_10900_14480.n80 a_10900_14480.n21 9.3005
R6614 a_10900_14480.n80 a_10900_14480.n20 9.3005
R6615 a_10900_14480.n80 a_10900_14480.n22 9.3005
R6616 a_10900_14480.n81 a_10900_14480.n80 9.3005
R6617 a_10900_14480.n128 a_10900_14480.n3 9.3005
R6618 a_10900_14480.n128 a_10900_14480.n4 9.3005
R6619 a_10900_14480.n128 a_10900_14480.n2 9.3005
R6620 a_10900_14480.n128 a_10900_14480.n5 9.3005
R6621 a_10900_14480.n128 a_10900_14480.n127 9.3005
R6622 a_10900_14480.n115 a_10900_14480.n4 9.3005
R6623 a_10900_14480.n115 a_10900_14480.n2 9.3005
R6624 a_10900_14480.n115 a_10900_14480.n5 9.3005
R6625 a_10900_14480.n127 a_10900_14480.n115 9.3005
R6626 a_10900_14480.n113 a_10900_14480.n4 9.3005
R6627 a_10900_14480.n113 a_10900_14480.n2 9.3005
R6628 a_10900_14480.n113 a_10900_14480.n5 9.3005
R6629 a_10900_14480.n124 a_10900_14480.n113 9.3005
R6630 a_10900_14480.n127 a_10900_14480.n113 9.3005
R6631 a_10900_14480.n127 a_10900_14480.n126 9.3005
R6632 a_10900_14480.n126 a_10900_14480.n124 9.3005
R6633 a_10900_14480.n126 a_10900_14480.n5 9.3005
R6634 a_10900_14480.n126 a_10900_14480.n2 9.3005
R6635 a_10900_14480.n127 a_10900_14480.n7 9.3005
R6636 a_10900_14480.n124 a_10900_14480.n7 9.3005
R6637 a_10900_14480.n7 a_10900_14480.n5 9.3005
R6638 a_10900_14480.n7 a_10900_14480.n2 9.3005
R6639 a_10900_14480.n7 a_10900_14480.n3 9.3005
R6640 a_10900_14480.n4 a_10900_14480.n0 9.3005
R6641 a_10900_14480.n2 a_10900_14480.n0 9.3005
R6642 a_10900_14480.n5 a_10900_14480.n0 9.3005
R6643 a_10900_14480.n124 a_10900_14480.n0 9.3005
R6644 a_10900_14480.n127 a_10900_14480.n0 9.3005
R6645 a_10900_14480.n79 a_10900_14480.n19 4.64654
R6646 a_10900_14480.n66 a_10900_14480.n20 4.64654
R6647 a_10900_14480.n77 a_10900_14480.n18 4.64654
R6648 a_10900_14480.n68 a_10900_14480.n21 4.64654
R6649 a_10900_14480.n78 a_10900_14480.n77 4.64654
R6650 a_10900_14480.n124 a_10900_14480.n1 4.64654
R6651 a_10900_14480.n114 a_10900_14480.n3 4.64654
R6652 a_10900_14480.n116 a_10900_14480.n4 4.64654
R6653 a_10900_14480.n125 a_10900_14480.n3 4.64654
R6654 a_10900_14480.n107 a_10900_14480.n106 2.36206
R6655 a_10900_14480.n93 a_10900_14480.n92 2.36206
R6656 a_10900_14480.n44 a_10900_14480.n35 2.36206
R6657 a_10900_14480.n56 a_10900_14480.n55 2.36206
R6658 a_10900_14480.n104 a_10900_14480.n103 2.19742
R6659 a_10900_14480.n91 a_10900_14480.n90 2.19742
R6660 a_10900_14480.n46 a_10900_14480.n45 2.19742
R6661 a_10900_14480.n58 a_10900_14480.n57 2.19742
R6662 a_10900_14480.n111 a_10900_14480.n110 1.80838
R6663 a_10900_14480.n39 a_10900_14480.n37 1.80838
R6664 a_10900_14480.n84 a_10900_14480.n17 1.56363
R6665 a_10900_14480.n26 a_10900_14480.n24 1.56363
R6666 a_10900_14480.n27 a_10900_14480.n25 1.5505
R6667 a_10900_14480.n62 a_10900_14480.n61 1.5505
R6668 a_10900_14480.n33 a_10900_14480.n32 1.5505
R6669 a_10900_14480.n50 a_10900_14480.n49 1.5505
R6670 a_10900_14480.n52 a_10900_14480.n51 1.5505
R6671 a_10900_14480.n54 a_10900_14480.n29 1.5505
R6672 a_10900_14480.n43 a_10900_14480.n42 1.5505
R6673 a_10900_14480.n37 a_10900_14480.n36 1.5505
R6674 a_10900_14480.n89 a_10900_14480.n15 1.5505
R6675 a_10900_14480.n87 a_10900_14480.n86 1.5505
R6676 a_10900_14480.n102 a_10900_14480.n10 1.5505
R6677 a_10900_14480.n100 a_10900_14480.n99 1.5505
R6678 a_10900_14480.n98 a_10900_14480.n97 1.5505
R6679 a_10900_14480.n14 a_10900_14480.n13 1.5505
R6680 a_10900_14480.n110 a_10900_14480.n8 1.5505
R6681 a_10900_14480.n105 a_10900_14480.n9 1.5505
R6682 a_10900_14480.n124 a_10900_14480.n123 1.25468
R6683 a_10900_14480.n109 a_10900_14480.n9 1.25468
R6684 a_10900_14480.n96 a_10900_14480.n14 1.25468
R6685 a_10900_14480.n70 a_10900_14480.n19 1.25468
R6686 a_10900_14480.n42 a_10900_14480.n41 1.25468
R6687 a_10900_14480.n54 a_10900_14480.n53 1.25468
R6688 a_10900_14480.n117 a_10900_14480.n4 1.19225
R6689 a_10900_14480.n103 a_10900_14480.n102 1.19225
R6690 a_10900_14480.n90 a_10900_14480.n89 1.19225
R6691 a_10900_14480.n76 a_10900_14480.n21 1.19225
R6692 a_10900_14480.n46 a_10900_14480.n33 1.19225
R6693 a_10900_14480.n58 a_10900_14480.n27 1.19225
R6694 a_10900_14480.n120 a_10900_14480.n5 1.07024
R6695 a_10900_14480.n97 a_10900_14480.n12 1.07024
R6696 a_10900_14480.n72 a_10900_14480.n22 1.07024
R6697 a_10900_14480.n52 a_10900_14480.n31 1.07024
R6698 a_10900_14480.n39 a_10900_14480.n38 1.04968
R6699 a_10900_14480.n112 a_10900_14480.n111 1.04968
R6700 a_10900_14480.n124 a_10900_14480.n6 1.0237
R6701 a_10900_14480.n107 a_10900_14480.n9 1.0237
R6702 a_10900_14480.n93 a_10900_14480.n14 1.0237
R6703 a_10900_14480.n23 a_10900_14480.n19 1.0237
R6704 a_10900_14480.n42 a_10900_14480.n35 1.0237
R6705 a_10900_14480.n55 a_10900_14480.n54 1.0237
R6706 a_10900_14480.n118 a_10900_14480.n4 0.959578
R6707 a_10900_14480.n102 a_10900_14480.n101 0.959578
R6708 a_10900_14480.n89 a_10900_14480.n88 0.959578
R6709 a_10900_14480.n74 a_10900_14480.n21 0.959578
R6710 a_10900_14480.n48 a_10900_14480.n33 0.959578
R6711 a_10900_14480.n60 a_10900_14480.n27 0.959578
R6712 a_10900_14480.n118 a_10900_14480.n2 0.885803
R6713 a_10900_14480.n101 a_10900_14480.n100 0.885803
R6714 a_10900_14480.n88 a_10900_14480.n87 0.885803
R6715 a_10900_14480.n74 a_10900_14480.n20 0.885803
R6716 a_10900_14480.n49 a_10900_14480.n48 0.885803
R6717 a_10900_14480.n61 a_10900_14480.n60 0.885803
R6718 a_10900_14480.n127 a_10900_14480.n6 0.812055
R6719 a_10900_14480.n81 a_10900_14480.n23 0.812055
R6720 a_10900_14480.n120 a_10900_14480.n2 0.77514
R6721 a_10900_14480.n100 a_10900_14480.n12 0.77514
R6722 a_10900_14480.n87 a_10900_14480.n17 0.77514
R6723 a_10900_14480.n72 a_10900_14480.n20 0.77514
R6724 a_10900_14480.n49 a_10900_14480.n31 0.77514
R6725 a_10900_14480.n61 a_10900_14480.n26 0.77514
R6726 a_10900_14480.n117 a_10900_14480.n3 0.647417
R6727 a_10900_14480.n77 a_10900_14480.n76 0.647417
R6728 a_10900_14480.n123 a_10900_14480.n5 0.590702
R6729 a_10900_14480.n110 a_10900_14480.n109 0.590702
R6730 a_10900_14480.n97 a_10900_14480.n96 0.590702
R6731 a_10900_14480.n70 a_10900_14480.n22 0.590702
R6732 a_10900_14480.n41 a_10900_14480.n37 0.590702
R6733 a_10900_14480.n53 a_10900_14480.n52 0.590702
R6734 a_10900_14480.n63 a_10900_14480.n24 0.530034
R6735 a_10900_14480.n85 a_10900_14480.n84 0.530034
R6736 a_10900_14480.t7 a_10900_14480.n121 0.290206
R6737 a_10900_14480.t8 a_10900_14480.n94 0.290206
R6738 a_10900_14480.t4 a_10900_14480.n83 0.290206
R6739 a_10900_14480.n73 a_10900_14480.t3 0.290206
R6740 a_10900_14480.n34 a_10900_14480.t5 0.290206
R6741 a_10900_14480.n28 a_10900_14480.t2 0.290206
R6742 a_10900_14480.n57 a_10900_14480.n56 0.154071
R6743 a_10900_14480.n45 a_10900_14480.n44 0.154071
R6744 a_10900_14480.n92 a_10900_14480.n91 0.154071
R6745 a_10900_14480.n106 a_10900_14480.n104 0.154071
R6746 a_10900_14480.n85 a_10900_14480.n82 0.137464
R6747 a_10900_14480.n113 a_10900_14480.n112 0.137464
R6748 a_10900_14480.n64 a_10900_14480.n63 0.134964
R6749 a_10900_14480.n38 a_10900_14480.n7 0.134964
R6750 a_10900_14480.n62 a_10900_14480.n25 0.0183571
R6751 a_10900_14480.n57 a_10900_14480.n25 0.0183571
R6752 a_10900_14480.n56 a_10900_14480.n29 0.0183571
R6753 a_10900_14480.n51 a_10900_14480.n29 0.0183571
R6754 a_10900_14480.n51 a_10900_14480.n50 0.0183571
R6755 a_10900_14480.n50 a_10900_14480.n32 0.0183571
R6756 a_10900_14480.n45 a_10900_14480.n32 0.0183571
R6757 a_10900_14480.n44 a_10900_14480.n43 0.0183571
R6758 a_10900_14480.n43 a_10900_14480.n36 0.0183571
R6759 a_10900_14480.n86 a_10900_14480.n15 0.0183571
R6760 a_10900_14480.n91 a_10900_14480.n15 0.0183571
R6761 a_10900_14480.n92 a_10900_14480.n13 0.0183571
R6762 a_10900_14480.n98 a_10900_14480.n13 0.0183571
R6763 a_10900_14480.n99 a_10900_14480.n98 0.0183571
R6764 a_10900_14480.n99 a_10900_14480.n10 0.0183571
R6765 a_10900_14480.n104 a_10900_14480.n10 0.0183571
R6766 a_10900_14480.n106 a_10900_14480.n105 0.0183571
R6767 a_10900_14480.n105 a_10900_14480.n8 0.0183571
R6768 a_10900_14480.n38 a_10900_14480.n36 0.0106786
R6769 a_10900_14480.n112 a_10900_14480.n8 0.0106786
R6770 a_10900_14480.n129 a_10900_14480.n0 0.0106786
R6771 a_10900_14480.n69 a_10900_14480.n68 0.00992001
R6772 a_10900_14480.n80 a_10900_14480.n78 0.00992001
R6773 a_10900_14480.n79 a_10900_14480.n65 0.00992001
R6774 a_10900_14480.n67 a_10900_14480.n66 0.00992001
R6775 a_10900_14480.n82 a_10900_14480.n18 0.00992001
R6776 a_10900_14480.n66 a_10900_14480.n65 0.00992001
R6777 a_10900_14480.n67 a_10900_14480.n18 0.00992001
R6778 a_10900_14480.n78 a_10900_14480.n69 0.00992001
R6779 a_10900_14480.n68 a_10900_14480.n64 0.00992001
R6780 a_10900_14480.n80 a_10900_14480.n79 0.00992001
R6781 a_10900_14480.n126 a_10900_14480.n116 0.00992001
R6782 a_10900_14480.n125 a_10900_14480.n0 0.00992001
R6783 a_10900_14480.n115 a_10900_14480.n1 0.00992001
R6784 a_10900_14480.n114 a_10900_14480.n113 0.00992001
R6785 a_10900_14480.n128 a_10900_14480.n1 0.00992001
R6786 a_10900_14480.n115 a_10900_14480.n114 0.00992001
R6787 a_10900_14480.n126 a_10900_14480.n125 0.00992001
R6788 a_10900_14480.n116 a_10900_14480.n7 0.00992001
R6789 a_10900_14480.n63 a_10900_14480.n62 0.00817857
R6790 a_10900_14480.n86 a_10900_14480.n85 0.00817857
R6791 a_10900_14480.n129 a_10900_14480.n128 0.00817857
R6792 a_10120_15820.t0 a_10120_15820.t1 178.133
R6793 a_21720_2700.n0 a_21720_2700.t2 399.724
R6794 a_21720_2700.t1 a_21720_2700.n1 359.615
R6795 a_21720_2700.n0 a_21720_2700.t3 319.39
R6796 a_21720_2700.n1 a_21720_2700.t0 243.16
R6797 a_21720_2700.n1 a_21720_2700.n0 3.08327
R6798 a_22130_3360.n0 a_22130_3360.t1 236.913
R6799 a_22130_3360.n0 a_22130_3360.t0 359.865
R6800 a_22130_3360.t2 a_22130_3360.n0 235.453
R6801 a_22240_2700.n0 a_22240_2700.t3 399.724
R6802 a_22240_2700.t1 a_22240_2700.n1 359.615
R6803 a_22240_2700.n0 a_22240_2700.t2 319.39
R6804 a_22240_2700.n1 a_22240_2700.t0 243.16
R6805 a_22240_2700.n1 a_22240_2700.n0 3.08327
R6806 a_22650_1940.t1 a_22650_1940.n0 134.684
R6807 a_22650_1940.n0 a_22650_1940.t0 243.054
R6808 a_22650_1940.n0 a_22650_1940.t2 135.409
R6809 ua1.t3 ua1.t6 401.668
R6810 ua1.n1 ua1.t5 399.724
R6811 ua1.n0 ua1.n2 366.81
R6812 ua1.t1 ua1.n3 359.615
R6813 ua1.n2 ua1.t2 353.467
R6814 ua1.n1 ua1.t4 319.39
R6815 ua1.n2 ua1.t3 257.067
R6816 ua1.n3 ua1.t0 243.16
R6817 ua1.n0 ua1.n1 2.03856
R6818 ua1.n3 ua1.n0 5.94143
R6819 a_22130_1940.t1 a_22130_1940.n0 134.684
R6820 a_22130_1940.n0 a_22130_1940.t0 243.054
R6821 a_22130_1940.n0 a_22130_1940.t2 135.409
R6822 a_13200_6670.t0 a_13200_6670.t1 39.4005
R6823 a_10780_3220.n3 a_10780_3220.t5 772.196
R6824 a_10780_3220.n1 a_10780_3220.t0 756.067
R6825 a_10780_3220.n4 a_10780_3220.n3 607.465
R6826 a_10780_3220.n0 a_10780_3220.t3 514.134
R6827 a_10780_3220.t5 a_10780_3220.t4 514.134
R6828 a_10780_3220.n1 a_10780_3220.n0 437.913
R6829 a_10780_3220.n2 a_10780_3220.t6 289.2
R6830 a_10780_3220.n0 a_10780_3220.t2 273.134
R6831 a_10780_3220.t1 a_10780_3220.n4 233
R6832 a_10780_3220.n3 a_10780_3220.n2 208.868
R6833 a_10780_3220.n2 a_10780_3220.t7 176.733
R6834 a_10780_3220.n4 a_10780_3220.n1 31.7872
R6835 a_18840_2930.n0 a_18840_2930.t3 750.201
R6836 a_18840_2930.n1 a_18840_2930.t4 349.433
R6837 a_18840_2930.n0 a_18840_2930.t0 276.733
R6838 a_18840_2930.n2 a_18840_2930.n1 206.333
R6839 a_18840_2930.n1 a_18840_2930.n0 48.0005
R6840 a_18840_2930.t2 a_18840_2930.n2 48.0005
R6841 a_18840_2930.n2 a_18840_2930.t1 48.0005
R6842 a_11860_5460.t7 a_11860_5460.t6 835.467
R6843 a_11860_5460.n2 a_11860_5460.t8 517.347
R6844 a_11860_5460.n0 a_11860_5460.t3 465.933
R6845 a_11860_5460.n1 a_11860_5460.n0 458.469
R6846 a_11860_5460.n1 a_11860_5460.t7 398.767
R6847 a_11860_5460.n0 a_11860_5460.t5 321.334
R6848 a_11860_5460.n5 a_11860_5460.n4 244.716
R6849 a_11860_5460.n2 a_11860_5460.t4 228.148
R6850 a_11860_5460.t2 a_11860_5460.n5 221.411
R6851 a_11860_5460.n3 a_11860_5460.n2 216
R6852 a_11860_5460.n5 a_11860_5460.n3 201.573
R6853 a_11860_5460.n3 a_11860_5460.n1 121.451
R6854 a_11860_5460.n4 a_11860_5460.t0 24.0005
R6855 a_11860_5460.n4 a_11860_5460.t1 24.0005
R6856 a_12650_3210.t0 a_12650_3210.t1 157.601
R6857 a_11780_5490.n2 a_11780_5490.n0 1319.38
R6858 a_11780_5490.t3 a_11780_5490.t5 1188.93
R6859 a_11780_5490.t5 a_11780_5490.t4 835.467
R6860 a_11780_5490.n0 a_11780_5490.t6 562.333
R6861 a_11780_5490.n2 a_11780_5490.n1 247.917
R6862 a_11780_5490.n0 a_11780_5490.t3 224.934
R6863 a_11780_5490.t1 a_11780_5490.n2 221.411
R6864 a_11780_5490.n1 a_11780_5490.t2 24.0005
R6865 a_11780_5490.n1 a_11780_5490.t0 24.0005
R6866 a_18390_10330.n1 a_18390_10330.t7 321.334
R6867 a_18390_10330.n5 a_18390_10330.n4 298.503
R6868 a_18390_10330.n2 a_18390_10330.n1 208.868
R6869 a_18390_10330.n4 a_18390_10330.n0 194.488
R6870 a_18390_10330.n3 a_18390_10330.t0 174.056
R6871 a_18390_10330.n4 a_18390_10330.n3 161.3
R6872 a_18390_10330.n2 a_18390_10330.t2 112.468
R6873 a_18390_10330.n1 a_18390_10330.t6 112.468
R6874 a_18390_10330.n3 a_18390_10330.n2 61.5894
R6875 a_18390_10330.n0 a_18390_10330.t3 60.0005
R6876 a_18390_10330.n0 a_18390_10330.t1 60.0005
R6877 a_18390_10330.n5 a_18390_10330.t4 49.2505
R6878 a_18390_10330.t5 a_18390_10330.n5 49.2505
R6879 a_11840_9460.n4 a_11840_9460.n3 314.526
R6880 a_11840_9460.n5 a_11840_9460.t12 287.762
R6881 a_11840_9460.n6 a_11840_9460.t10 287.762
R6882 a_11840_9460.n5 a_11840_9460.t9 287.589
R6883 a_11840_9460.n7 a_11840_9460.t11 287.012
R6884 a_11840_9460.n8 a_11840_9460.t8 287.012
R6885 a_11840_9460.t0 a_11840_9460.n10 117.817
R6886 a_11840_9460.n2 a_11840_9460.n0 107.079
R6887 a_11840_9460.n2 a_11840_9460.n1 104.829
R6888 a_11840_9460.n10 a_11840_9460.t7 47.7922
R6889 a_11840_9460.n3 a_11840_9460.t1 39.4005
R6890 a_11840_9460.n3 a_11840_9460.t2 39.4005
R6891 a_11840_9460.n0 a_11840_9460.t4 13.1338
R6892 a_11840_9460.n0 a_11840_9460.t6 13.1338
R6893 a_11840_9460.n1 a_11840_9460.t3 13.1338
R6894 a_11840_9460.n1 a_11840_9460.t5 13.1338
R6895 a_11840_9460.n10 a_11840_9460.n9 13.0943
R6896 a_11840_9460.n9 a_11840_9460.n4 10.7505
R6897 a_11840_9460.n9 a_11840_9460.n8 6.78086
R6898 a_11840_9460.n4 a_11840_9460.n2 2.0005
R6899 a_11840_9460.n7 a_11840_9460.n6 0.579071
R6900 a_11840_9460.n8 a_11840_9460.n7 0.282643
R6901 a_11840_9460.n6 a_11840_9460.n5 0.2755
R6902 a_21690_4400.n1 a_21690_4400.t1 247.257
R6903 a_21690_4400.n0 a_21690_4400.t2 240.543
R6904 a_21690_4400.n0 a_21690_4400.t3 198.746
R6905 a_21690_4400.n0 a_21690_4400.t5 197.934
R6906 a_21690_4400.n0 a_21690_4400.t4 197.934
R6907 a_21690_4400.t0 a_21690_4400.n1 139.434
R6908 a_21690_4400.n1 a_21690_4400.n0 6.1255
R6909 a_13720_5910.n1 a_13720_5910.n0 481.334
R6910 a_13720_5910.n0 a_13720_5910.t3 465.933
R6911 a_13720_5910.n0 a_13720_5910.t4 321.334
R6912 a_13720_5910.n2 a_13720_5910.n1 226.888
R6913 a_13720_5910.n1 a_13720_5910.t1 172.458
R6914 a_13720_5910.n2 a_13720_5910.t2 19.7005
R6915 a_13720_5910.t0 a_13720_5910.n2 19.7005
R6916 a_14160_5490.t0 a_14160_5490.n2 500.086
R6917 a_14160_5490.n1 a_14160_5490.n0 473.334
R6918 a_14160_5490.n0 a_14160_5490.t2 465.933
R6919 a_14160_5490.t0 a_14160_5490.n2 461.389
R6920 a_14160_5490.n0 a_14160_5490.t3 321.334
R6921 a_14160_5490.n1 a_14160_5490.t1 177.577
R6922 a_14160_5490.n2 a_14160_5490.n1 48.3898
R6923 a_21610_3360.n0 a_21610_3360.t1 236.913
R6924 a_21610_3360.n0 a_21610_3360.t2 359.865
R6925 a_21610_3360.t0 a_21610_3360.n0 235.453
R6926 a_15710_6670.n0 a_15710_6670.t3 605.311
R6927 a_15710_6670.t3 a_15710_6670.t0 420.202
R6928 a_15710_6670.t1 a_15710_6670.n0 240.327
R6929 a_15710_6670.n0 a_15710_6670.t2 148.734
R6930 a_13280_3020.n2 a_13280_3020.t3 761.4
R6931 a_13280_3020.n1 a_13280_3020.t4 350.349
R6932 a_13280_3020.t2 a_13280_3020.n2 254.333
R6933 a_13280_3020.n1 a_13280_3020.n0 206.333
R6934 a_13280_3020.n2 a_13280_3020.n1 70.4005
R6935 a_13280_3020.n0 a_13280_3020.t0 48.0005
R6936 a_13280_3020.n0 a_13280_3020.t1 48.0005
R6937 a_18410_9620.n10 a_18410_9620.t8 486.038
R6938 a_18410_9620.n6 a_18410_9620.t12 317.317
R6939 a_18410_9620.n0 a_18410_9620.t11 317.317
R6940 a_18410_9620.n7 a_18410_9620.n6 257.067
R6941 a_18410_9620.n1 a_18410_9620.n0 257.067
R6942 a_18410_9620.n5 a_18410_9620.n4 257.067
R6943 a_18410_9620.n9 a_18410_9620.n8 152
R6944 a_18410_9620.n11 a_18410_9620.n2 152
R6945 a_18410_9620.n9 a_18410_9620.n3 117.781
R6946 a_18410_9620.n12 a_18410_9620.n11 117.781
R6947 a_18410_9620.n8 a_18410_9620.n7 85.6894
R6948 a_18410_9620.n2 a_18410_9620.n1 85.6894
R6949 a_18410_9620.n4 a_18410_9620.n2 85.6894
R6950 a_18410_9620.n8 a_18410_9620.n5 85.6894
R6951 a_18410_9620.n6 a_18410_9620.t10 60.2505
R6952 a_18410_9620.n7 a_18410_9620.t0 60.2505
R6953 a_18410_9620.n0 a_18410_9620.t9 60.2505
R6954 a_18410_9620.n1 a_18410_9620.t2 60.2505
R6955 a_18410_9620.n4 a_18410_9620.t6 60.2505
R6956 a_18410_9620.n5 a_18410_9620.t4 60.2505
R6957 a_18410_9620.n11 a_18410_9620.n10 25.6005
R6958 a_18410_9620.n3 a_18410_9620.t5 24.0005
R6959 a_18410_9620.n3 a_18410_9620.t1 24.0005
R6960 a_18410_9620.n10 a_18410_9620.n9 24.0005
R6961 a_18410_9620.n12 a_18410_9620.t3 24.0005
R6962 a_18410_9620.t7 a_18410_9620.n12 24.0005
R6963 a_14340_6640.n0 a_14340_6640.t3 465.933
R6964 a_14340_6640.n1 a_14340_6640.n0 431.824
R6965 a_14340_6640.n0 a_14340_6640.t2 321.334
R6966 a_14340_6640.t0 a_14340_6640.n1 288.37
R6967 a_14340_6640.n1 a_14340_6640.t1 177.577
R6968 a_13800_2890.n0 a_13800_2890.t1 663.801
R6969 a_13800_2890.t0 a_13800_2890.n0 397.053
R6970 a_13800_2890.n0 a_13800_2890.t2 348.851
R6971 a_13910_2890.t0 a_13910_2890.t1 96.0005
R6972 a_16000_5490.n4 a_16000_5490.t3 297.233
R6973 a_16000_5490.t6 a_16000_5490.n5 297.233
R6974 a_16000_5490.n3 a_16000_5490.n1 257.067
R6975 a_16000_5490.n0 a_16000_5490.t2 241.928
R6976 a_16000_5490.n7 a_16000_5490.n6 237.728
R6977 a_16000_5490.t1 a_16000_5490.n7 235.528
R6978 a_16000_5490.n6 a_16000_5490.n1 226.942
R6979 a_16000_5490.n3 a_16000_5490.n2 226.942
R6980 a_16000_5490.n2 a_16000_5490.t7 220.505
R6981 a_16000_5490.n5 a_16000_5490.n4 216.9
R6982 a_16000_5490.n0 a_16000_5490.t0 145.536
R6983 a_16000_5490.n7 a_16000_5490.n0 121.6
R6984 a_16000_5490.n2 a_16000_5490.t3 92.3838
R6985 a_16000_5490.n6 a_16000_5490.t6 92.3838
R6986 a_16000_5490.t4 a_16000_5490.n3 80.3338
R6987 a_16000_5490.n4 a_16000_5490.t4 80.3338
R6988 a_16000_5490.t5 a_16000_5490.n1 80.3338
R6989 a_16000_5490.n5 a_16000_5490.t5 80.3338
R6990 a_14890_17428.t0 a_14890_17428.t1 178.133
R6991 a_14770_15820.t0 a_14770_15820.t1 178.133
R6992 a_11430_2890.n0 a_11430_2890.t1 663.801
R6993 a_11430_2890.t0 a_11430_2890.n0 397.053
R6994 a_11430_2890.n0 a_11430_2890.t2 355.378
R6995 a_11540_2890.t0 a_11540_2890.t1 96.0005
R6996 a_10000_17428.t0 a_10000_17428.t1 178.133
R6997 a_17030_3180.t5 a_17030_3180.t2 1012.2
R6998 a_17030_3180.n0 a_17030_3180.t0 663.801
R6999 a_17030_3180.n2 a_17030_3180.n1 431.401
R7000 a_17030_3180.t6 a_17030_3180.t3 401.668
R7001 a_17030_3180.n0 a_17030_3180.t5 361.692
R7002 a_17030_3180.t1 a_17030_3180.n2 298.921
R7003 a_17030_3180.n1 a_17030_3180.t6 257.067
R7004 a_17030_3180.n1 a_17030_3180.t4 208.868
R7005 a_17030_3180.n2 a_17030_3180.n0 67.2005
R7006 a_18250_2800.t0 a_18250_2800.t1 96.0005
R7007 pll_bgr_magic_3_0.VV3.n7 pll_bgr_magic_3_0.VV3.n6 959.696
R7008 pll_bgr_magic_3_0.VV3.n2 pll_bgr_magic_3_0.VV3.n0 297.503
R7009 pll_bgr_magic_3_0.VV3.n6 pll_bgr_magic_3_0.VV3.t7 289.2
R7010 pll_bgr_magic_3_0.VV3.n5 pll_bgr_magic_3_0.VV3.t6 289.2
R7011 pll_bgr_magic_3_0.VV3.n4 pll_bgr_magic_3_0.VV3.t5 289.2
R7012 pll_bgr_magic_3_0.VV3.n3 pll_bgr_magic_3_0.VV3.t8 232.968
R7013 pll_bgr_magic_3_0.VV3.n6 pll_bgr_magic_3_0.VV3.n5 208.868
R7014 pll_bgr_magic_3_0.VV3.n5 pll_bgr_magic_3_0.VV3.n4 208.868
R7015 pll_bgr_magic_3_0.VV3.n4 pll_bgr_magic_3_0.VV3.n3 199.829
R7016 pll_bgr_magic_3_0.VV3.n2 pll_bgr_magic_3_0.VV3.n1 195.55
R7017 pll_bgr_magic_3_0.VV3.n3 pll_bgr_magic_3_0.VV3.n2 172.582
R7018 pll_bgr_magic_3_0.VV3.n1 pll_bgr_magic_3_0.VV3.t0 60.0005
R7019 pll_bgr_magic_3_0.VV3.n1 pll_bgr_magic_3_0.VV3.t1 60.0005
R7020 pll_bgr_magic_3_0.VV3.n7 pll_bgr_magic_3_0.VV3.t2 50.6672
R7021 pll_bgr_magic_3_0.VV3.n0 pll_bgr_magic_3_0.VV3.t4 49.2505
R7022 pll_bgr_magic_3_0.VV3.n0 pll_bgr_magic_3_0.VV3.t3 49.2505
R7023 pll_bgr_magic_3_0.VV3 pll_bgr_magic_3_0.VV3.n7 1.82907
R7024 a_15160_2860.n4 a_15160_2860.n3 742.51
R7025 a_15160_2860.n0 a_15160_2860.t0 723.534
R7026 a_15160_2860.t1 a_15160_2860.n9 723.534
R7027 a_15160_2860.n3 a_15160_2860.n2 684.806
R7028 a_15160_2860.n8 a_15160_2860.n7 366.856
R7029 a_15160_2860.n1 a_15160_2860.t11 337.401
R7030 a_15160_2860.n1 a_15160_2860.t5 305.267
R7031 a_15160_2860.n0 a_15160_2860.t2 254.333
R7032 a_15160_2860.n5 a_15160_2860.n4 224.934
R7033 a_15160_2860.n8 a_15160_2860.t8 190.123
R7034 a_15160_2860.n9 a_15160_2860.n8 187.201
R7035 a_15160_2860.n2 a_15160_2860.n1 176.733
R7036 a_15160_2860.n7 a_15160_2860.n6 176.733
R7037 a_15160_2860.n6 a_15160_2860.n5 176.733
R7038 a_15160_2860.n4 a_15160_2860.t9 144.601
R7039 a_15160_2860.n3 a_15160_2860.t4 131.976
R7040 a_15160_2860.n1 a_15160_2860.t10 128.534
R7041 a_15160_2860.n2 a_15160_2860.t3 128.534
R7042 a_15160_2860.n5 a_15160_2860.t7 112.468
R7043 a_15160_2860.n6 a_15160_2860.t12 112.468
R7044 a_15160_2860.n7 a_15160_2860.t6 112.468
R7045 a_15160_2860.n9 a_15160_2860.n0 70.4005
R7046 a_15050_2860.n2 a_15050_2860.t0 723.534
R7047 a_15050_2860.n1 a_15050_2860.t4 553.534
R7048 a_15050_2860.t3 a_15050_2860.n2 254.333
R7049 a_15050_2860.n1 a_15050_2860.n0 206.333
R7050 a_15050_2860.n2 a_15050_2860.n1 70.4005
R7051 a_15050_2860.n0 a_15050_2860.t1 48.0005
R7052 a_15050_2860.n0 a_15050_2860.t2 48.0005
R7053 a_21610_1940.t0 a_21610_1940.n0 134.684
R7054 a_21610_1940.n0 a_21610_1940.t2 243.054
R7055 a_21610_1940.n0 a_21610_1940.t1 135.409
R7056 a_22650_3360.n0 a_22650_3360.t2 236.913
R7057 a_22650_3360.n0 a_22650_3360.t0 359.865
R7058 a_22650_3360.t1 a_22650_3360.n0 235.453
R7059 a_16650_3100.n0 a_16650_3100.t1 713.933
R7060 a_16650_3100.n0 a_16650_3100.t2 314.233
R7061 a_16650_3100.t0 a_16650_3100.n0 308.2
R7062 a_9570_17278.t0 a_9570_17278.t1 178.133
R7063 a_15288_18640.t0 a_15288_18640.t1 165.826
R7064 a_15850_2890.t0 a_15850_2890.t1 96.0005
R7065 a_15380_3150.n0 a_15380_3150.t2 685.134
R7066 a_15380_3150.n1 a_15380_3150.t0 663.801
R7067 a_15380_3150.n0 a_15380_3150.t3 534.268
R7068 a_15380_3150.t1 a_15380_3150.n1 362.921
R7069 a_15380_3150.n1 a_15380_3150.n0 91.7338
R7070 a_16950_2890.t0 a_16950_2890.t1 96.0005
R7071 a_13990_2860.t1 a_13990_2860.n2 755.534
R7072 a_13990_2860.n2 a_13990_2860.t0 685.134
R7073 a_13990_2860.n1 a_13990_2860.n0 389.733
R7074 a_13990_2860.n1 a_13990_2860.t2 340.2
R7075 a_13990_2860.n0 a_13990_2860.t3 321.334
R7076 a_13990_2860.n0 a_13990_2860.t4 144.601
R7077 a_13990_2860.n2 a_13990_2860.n1 19.2005
R7078 pll_bgr_magic_3_0.VV2.n0 pll_bgr_magic_3_0.VV2.t0 133.959
R7079 pll_bgr_magic_3_0.VV2.n0 pll_bgr_magic_3_0.VV2.t1 50.6672
R7080 pll_bgr_magic_3_0.VV2 pll_bgr_magic_3_0.VV2.n0 7.31479
R7081 a_12560_13480.t0 a_12560_13480.t1 178.194
R7082 a_13280_5460.n1 a_13280_5460.t3 562.333
R7083 a_13280_5460.t0 a_13280_5460.n4 500.086
R7084 a_13280_5460.t0 a_13280_5460.n4 461.389
R7085 a_13280_5460.n2 a_13280_5460.n1 453.315
R7086 a_13280_5460.n0 a_13280_5460.t4 417.733
R7087 a_13280_5460.n2 a_13280_5460.n0 388.639
R7088 a_13280_5460.n0 a_13280_5460.t2 369.534
R7089 a_13280_5460.n1 a_13280_5460.t5 224.934
R7090 a_13280_5460.n3 a_13280_5460.t1 172.458
R7091 a_13280_5460.n4 a_13280_5460.n3 43.2699
R7092 a_13280_5460.n3 a_13280_5460.n2 13.4217
R7093 a_15710_5490.n1 a_15710_5490.n0 409.067
R7094 a_15710_5490.n0 a_15710_5490.t2 403.38
R7095 a_15710_5490.n0 a_15710_5490.t3 369.534
R7096 a_15710_5490.t0 a_15710_5490.n1 209.928
R7097 a_15710_5490.n1 a_15710_5490.t1 177.536
R7098 a_12300_5910.t0 a_12300_5910.t1 39.4005
R7099 a_14690_3160.n0 a_14690_3160.t0 663.801
R7100 a_14690_3160.t4 a_14690_3160.t2 514.134
R7101 a_14690_3160.n0 a_14690_3160.t4 479.284
R7102 a_14690_3160.n3 a_14690_3160.n2 344.8
R7103 a_14690_3160.n1 a_14690_3160.t3 289.2
R7104 a_14690_3160.t1 a_14690_3160.n3 275.454
R7105 a_14690_3160.n2 a_14690_3160.t5 241
R7106 a_14690_3160.n1 a_14690_3160.t6 112.468
R7107 a_14690_3160.n3 a_14690_3160.n0 97.9205
R7108 a_14690_3160.n2 a_14690_3160.n1 64.2672
R7109 a_15740_2890.t0 a_15740_2890.t1 96.0005
R7110 ua[0].n0 ua[0].t0 514.134
R7111 ua[0] ua[0].n0 462.964
R7112 ua[0].n0 ua[0].t1 273.134
R7113 a_11780_5910.t0 a_11780_5910.t1 39.4005
R7114 a_11780_6670.t0 a_11780_6670.t1 39.4005
R7115 a_9690_16200.t0 a_9690_16200.t1 178.133
R7116 a_13720_5490.t0 a_13720_5490.t1 48.0005
R7117 pll_bgr_magic_3_0.VV4.n0 pll_bgr_magic_3_0.VV4.t0 178.577
R7118 pll_bgr_magic_3_0.VV4.n0 pll_bgr_magic_3_0.VV4.t1 50.6672
R7119 pll_bgr_magic_3_0.VV4 pll_bgr_magic_3_0.VV4.n0 2.92621
C0 pll_bgr_magic_3_0.VV2 V_CONT 0.455425f
C1 pll_bgr_magic_3_0.VV1 VDPWR 0.063069f
C2 pll_bgr_magic_3_0.VV4 VDPWR 0.08361f
C3 pll_bgr_magic_3_0.VV1 V_CONT 0.496053f
C4 pll_bgr_magic_3_0.VV3 VDPWR 1.07562f
C5 pll_bgr_magic_3_0.VV4 V_CONT 0.397769f
C6 pll_bgr_magic_3_0.VV1 pll_bgr_magic_3_0.VV2 0.034878f
C7 pll_bgr_magic_3_0.VV2 pll_bgr_magic_3_0.VV4 0.362952f
C8 VDPWR ua[0] 0.352654f
C9 V_CONT VDPWR 1.43423f
C10 pll_bgr_magic_3_0.VV1 pll_bgr_magic_3_0.VV3 0.389599f
C11 pll_bgr_magic_3_0.VV4 pll_bgr_magic_3_0.VV3 0.023643f
C12 V_CONT ua[0] 0.050598f
C13 ua[0] VGND 14.351799f
C14 VDPWR VGND 0.174356p
C15 pll_bgr_magic_3_0.VV2 VGND 3.31398f
C16 pll_bgr_magic_3_0.VV1 VGND 2.26609f
C17 pll_bgr_magic_3_0.VV3 VGND 1.23229f
C18 pll_bgr_magic_3_0.VV4 VGND 3.44556f
C19 V_CONT VGND 38.102207f
C20 a_15710_5490.t1 VGND 0.023659f
C21 a_15710_5490.t2 VGND 2.0362f
C22 a_15710_5490.n0 VGND 0.026464f
C23 a_15710_5490.n1 VGND 0.060553f
C24 a_15710_5490.t0 VGND 0.044187f
C25 a_15288_18640.t1 VGND 5.9975f
C26 a_15710_6670.t2 VGND 0.034319f
C27 a_15710_6670.t0 VGND 1.73994f
C28 a_15710_6670.t3 VGND 0.042516f
C29 a_15710_6670.n0 VGND 0.102101f
C30 a_15710_6670.t1 VGND 0.08112f
C31 a_21690_4400.n0 VGND 1.04311f
C32 a_21690_4400.t3 VGND 0.499058f
C33 a_21690_4400.t4 VGND 0.498316f
C34 a_21690_4400.t5 VGND 0.498316f
C35 a_21690_4400.t2 VGND 0.094724f
C36 a_21690_4400.t1 VGND 0.492622f
C37 a_21690_4400.n1 VGND 0.706776f
C38 a_21690_4400.t0 VGND 0.067077f
C39 a_11840_9460.t4 VGND 0.044358f
C40 a_11840_9460.t6 VGND 0.044358f
C41 a_11840_9460.n0 VGND 0.11867f
C42 a_11840_9460.t3 VGND 0.044358f
C43 a_11840_9460.t5 VGND 0.044358f
C44 a_11840_9460.n1 VGND 0.107634f
C45 a_11840_9460.n2 VGND 1.21683f
C46 a_11840_9460.t1 VGND 0.014786f
C47 a_11840_9460.t2 VGND 0.014786f
C48 a_11840_9460.n3 VGND 0.041682f
C49 a_11840_9460.n4 VGND 0.860437f
C50 a_11840_9460.t9 VGND 0.024477f
C51 a_11840_9460.t12 VGND 0.023979f
C52 a_11840_9460.n5 VGND 0.186829f
C53 a_11840_9460.t10 VGND 0.023979f
C54 a_11840_9460.n6 VGND 0.099745f
C55 a_11840_9460.t11 VGND 0.024302f
C56 a_11840_9460.n7 VGND 0.100457f
C57 a_11840_9460.t8 VGND 0.024302f
C58 a_11840_9460.n8 VGND 0.34311f
C59 a_11840_9460.n9 VGND 0.545948f
C60 a_11840_9460.t7 VGND 3.3892f
C61 a_11840_9460.n10 VGND 3.47416f
C62 a_11840_9460.t0 VGND 0.187264f
C63 a_10751_12090.t11 VGND 0.022048f
C64 a_10751_12090.t10 VGND 0.022048f
C65 a_10751_12090.n0 VGND 0.048589f
C66 a_10751_12090.t5 VGND 0.022048f
C67 a_10751_12090.t2 VGND 0.022048f
C68 a_10751_12090.n1 VGND 0.048287f
C69 a_10751_12090.n2 VGND 0.562362f
C70 a_10751_12090.t6 VGND 0.022048f
C71 a_10751_12090.t9 VGND 0.022048f
C72 a_10751_12090.n3 VGND 0.048287f
C73 a_10751_12090.n4 VGND 0.296766f
C74 a_10751_12090.t4 VGND 0.022048f
C75 a_10751_12090.t8 VGND 0.022048f
C76 a_10751_12090.n5 VGND 0.048287f
C77 a_10751_12090.n6 VGND 0.296766f
C78 a_10751_12090.t3 VGND 0.022048f
C79 a_10751_12090.t7 VGND 0.022048f
C80 a_10751_12090.n7 VGND 0.048287f
C81 a_10751_12090.n8 VGND 0.296766f
C82 a_10751_12090.t1 VGND 0.022048f
C83 a_10751_12090.t12 VGND 0.022048f
C84 a_10751_12090.n9 VGND 0.048287f
C85 a_10751_12090.n10 VGND 1.16667f
C86 a_10751_12090.t14 VGND 0.033898f
C87 a_10751_12090.t17 VGND 0.033832f
C88 a_10751_12090.n11 VGND 0.237966f
C89 a_10751_12090.t13 VGND 0.033832f
C90 a_10751_12090.n12 VGND 0.147954f
C91 a_10751_12090.t16 VGND 0.033832f
C92 a_10751_12090.n13 VGND 0.147954f
C93 a_10751_12090.t15 VGND 0.033832f
C94 a_10751_12090.n14 VGND 0.489729f
C95 a_10751_12090.n15 VGND 5.43823f
C96 a_10751_12090.t0 VGND 0.695008f
C97 a_10030_11260.n0 VGND 0.360667f
C98 a_10030_11260.n1 VGND 0.360667f
C99 a_10030_11260.n2 VGND 0.360667f
C100 a_10030_11260.n3 VGND 0.454298f
C101 a_10030_11260.n4 VGND 0.180333f
C102 a_10030_11260.n5 VGND 0.360667f
C103 a_10030_11260.n6 VGND 0.360667f
C104 a_10030_11260.n7 VGND 0.360667f
C105 a_10030_11260.n8 VGND 1.23779f
C106 a_10030_11260.n9 VGND 0.360667f
C107 a_10030_11260.t17 VGND 0.024727f
C108 a_10030_11260.t3 VGND 0.010305f
C109 a_10030_11260.t6 VGND 0.010305f
C110 a_10030_11260.n10 VGND 0.022597f
C111 a_10030_11260.n11 VGND 0.245331f
C112 a_10030_11260.t32 VGND 0.015954f
C113 a_10030_11260.t21 VGND 0.015954f
C114 a_10030_11260.n12 VGND 0.030906f
C115 a_10030_11260.n13 VGND 0.119581f
C116 a_10030_11260.t18 VGND 0.024402f
C117 a_10030_11260.t28 VGND 0.41219f
C118 a_10030_11260.t24 VGND 0.419031f
C119 a_10030_11260.t31 VGND 0.41219f
C120 a_10030_11260.t12 VGND 0.41219f
C121 a_10030_11260.t36 VGND 0.41219f
C122 a_10030_11260.t16 VGND 0.41219f
C123 a_10030_11260.t11 VGND 0.41219f
C124 a_10030_11260.t34 VGND 0.41219f
C125 a_10030_11260.t15 VGND 0.41219f
C126 a_10030_11260.t22 VGND 0.41219f
C127 a_10030_11260.t20 VGND 0.41219f
C128 a_10030_11260.t14 VGND 0.41219f
C129 a_10030_11260.t33 VGND 0.41219f
C130 a_10030_11260.t25 VGND 0.41219f
C131 a_10030_11260.t29 VGND 0.41219f
C132 a_10030_11260.t35 VGND 0.41219f
C133 a_10030_11260.t26 VGND 0.41219f
C134 a_10030_11260.t30 VGND 0.41219f
C135 a_10030_11260.t23 VGND 0.41219f
C136 a_10030_11260.t19 VGND 0.41219f
C137 a_10030_11260.n14 VGND 0.949966f
C138 a_10030_11260.t7 VGND 0.010305f
C139 a_10030_11260.t4 VGND 0.010305f
C140 a_10030_11260.n15 VGND 0.022597f
C141 a_10030_11260.n16 VGND 0.215201f
C142 a_10030_11260.t9 VGND 0.018148f
C143 a_10030_11260.n17 VGND 0.013021f
C144 a_10030_11260.n18 VGND 0.012563f
C145 a_10030_11260.n19 VGND 0.335083f
C146 a_10030_11260.n20 VGND 0.110146f
C147 a_10030_11260.t13 VGND 0.015954f
C148 a_10030_11260.t27 VGND 0.015954f
C149 a_10030_11260.n21 VGND 0.029642f
C150 a_10030_11260.n22 VGND 0.06623f
C151 a_10030_11260.n23 VGND 0.074194f
C152 a_10030_11260.n24 VGND 0.169072f
C153 a_10030_11260.t5 VGND 0.010305f
C154 a_10030_11260.n25 VGND 0.022597f
C155 a_10030_11260.t8 VGND 0.010305f
C156 a_10160_10990.t13 VGND 0.02f
C157 a_10160_10990.t21 VGND 0.02f
C158 a_10160_10990.t18 VGND 0.032283f
C159 a_10160_10990.n0 VGND 0.036051f
C160 a_10160_10990.n1 VGND 0.024627f
C161 a_10160_10990.t5 VGND 0.025389f
C162 a_10160_10990.n2 VGND 0.039854f
C163 a_10160_10990.t14 VGND 0.016667f
C164 a_10160_10990.t6 VGND 0.016667f
C165 a_10160_10990.n3 VGND 0.034125f
C166 a_10160_10990.n4 VGND 0.176664f
C167 a_10160_10990.n5 VGND 0.017774f
C168 a_10160_10990.t3 VGND 0.031554f
C169 a_10160_10990.n6 VGND 0.019781f
C170 a_10160_10990.n7 VGND 0.511999f
C171 a_10160_10990.n8 VGND 0.172226f
C172 a_10160_10990.t11 VGND 0.02f
C173 a_10160_10990.t20 VGND 0.02f
C174 a_10160_10990.t17 VGND 0.032283f
C175 a_10160_10990.n9 VGND 0.036051f
C176 a_10160_10990.n10 VGND 0.024627f
C177 a_10160_10990.t9 VGND 0.025389f
C178 a_10160_10990.n11 VGND 0.039854f
C179 a_10160_10990.t12 VGND 0.016667f
C180 a_10160_10990.t10 VGND 0.016667f
C181 a_10160_10990.n12 VGND 0.034125f
C182 a_10160_10990.n13 VGND 0.221004f
C183 a_10160_10990.n14 VGND 0.242013f
C184 a_10160_10990.t15 VGND 0.02f
C185 a_10160_10990.t19 VGND 0.02f
C186 a_10160_10990.t22 VGND 0.032283f
C187 a_10160_10990.n15 VGND 0.036051f
C188 a_10160_10990.n16 VGND 0.024627f
C189 a_10160_10990.t7 VGND 0.025389f
C190 a_10160_10990.n17 VGND 0.039854f
C191 a_10160_10990.n18 VGND 0.176664f
C192 a_10160_10990.t8 VGND 0.016667f
C193 a_10160_10990.n19 VGND 0.034125f
C194 a_10160_10990.t16 VGND 0.016667f
C195 a_15790_17280.t4 VGND 0.31433f
C196 a_15790_17280.t1 VGND 0.331199f
C197 a_15790_17280.t15 VGND 0.331199f
C198 a_15790_17280.t18 VGND 0.331199f
C199 a_15790_17280.t11 VGND 0.331199f
C200 a_15790_17280.t16 VGND 0.331199f
C201 a_15790_17280.t19 VGND 0.331199f
C202 a_15790_17280.t13 VGND 0.331199f
C203 a_15790_17280.t7 VGND 0.315469f
C204 a_15790_17280.t3 VGND 0.151964f
C205 a_15790_17280.n0 VGND 0.19601f
C206 a_15790_17280.t17 VGND 0.344559f
C207 a_15790_17280.t2 VGND 0.316794f
C208 a_15790_17280.t6 VGND 0.331199f
C209 a_15790_17280.t12 VGND 0.331199f
C210 a_15790_17280.t9 VGND 0.331199f
C211 a_15790_17280.t5 VGND 0.331199f
C212 a_15790_17280.t10 VGND 0.331199f
C213 a_15790_17280.t8 VGND 0.331199f
C214 a_15790_17280.t14 VGND 0.331199f
C215 a_15790_17280.t0 VGND 0.722653f
C216 a_15790_17280.t20 VGND 0.101437f
C217 a_18390_5940.n0 VGND 1.21839f
C218 a_18390_5940.t0 VGND 0.020492f
C219 a_18390_5940.t5 VGND 0.020492f
C220 a_18390_5940.t4 VGND 0.020492f
C221 a_18390_5940.n1 VGND 0.070101f
C222 a_18390_5940.n2 VGND 0.020862f
C223 a_18390_5940.t9 VGND 0.011978f
C224 a_18390_5940.n3 VGND 0.022994f
C225 a_18390_5940.n4 VGND 0.620084f
C226 a_18390_5940.t2 VGND 0.020492f
C227 a_18390_5940.t1 VGND 0.020492f
C228 a_18390_5940.n5 VGND 0.046427f
C229 a_18390_5940.n6 VGND 0.046427f
C230 a_18390_5940.t3 VGND 0.020492f
C231 a_15870_5490.t12 VGND 3.02742f
C232 a_15870_5490.t14 VGND 3.02613f
C233 a_15870_5490.n1 VGND 0.012413f
C234 a_15870_5490.n2 VGND 0.040951f
C235 a_15870_5490.n3 VGND 0.027173f
C236 a_15870_5490.n4 VGND 0.019604f
C237 a_15870_5490.t13 VGND 0.040684f
C238 a_15870_5490.t15 VGND 0.040684f
C239 a_15870_5490.t10 VGND 0.017772f
C240 a_15870_5490.n5 VGND 0.021423f
C241 a_15870_5490.n6 VGND 0.021423f
C242 a_15870_5490.t11 VGND 0.017772f
C243 a_15870_5490.n7 VGND 0.019604f
C244 a_15870_5490.t4 VGND 0.038007f
C245 a_15870_5490.t1 VGND 0.012002f
C246 a_15870_5490.n9 VGND 0.059042f
C247 a_15870_5490.n10 VGND 0.712029f
C248 a_15870_5490.n11 VGND 0.336097f
C249 a_15870_5490.n12 VGND 0.026477f
C250 a_15870_5490.n14 VGND 0.030457f
C251 a_12960_8860.n0 VGND 0.733925f
C252 a_12960_8860.n1 VGND 0.517552f
C253 a_12960_8860.t15 VGND 0.010076f
C254 a_12960_8860.t0 VGND 0.073183f
C255 a_12960_8860.t17 VGND 0.089231f
C256 a_12960_8860.n2 VGND 0.154524f
C257 a_12960_8860.t14 VGND 0.025191f
C258 a_12960_8860.t12 VGND 0.025191f
C259 a_12960_8860.n3 VGND 0.100278f
C260 a_12960_8860.t13 VGND 0.084832f
C261 a_12960_8860.t19 VGND 0.10958f
C262 a_12960_8860.t18 VGND 0.147001f
C263 a_12960_8860.n4 VGND 0.109992f
C264 a_12960_8860.n5 VGND 0.114936f
C265 a_12960_8860.t11 VGND 0.122253f
C266 a_12960_8860.n6 VGND 0.059573f
C267 a_12960_8860.n7 VGND 0.162248f
C268 a_12960_8860.n8 VGND 1.6251f
C269 a_12960_8860.t1 VGND 0.010076f
C270 a_12960_8860.t16 VGND 0.010076f
C271 a_12960_8860.n9 VGND 0.021428f
C272 a_12960_8860.t3 VGND 0.010076f
C273 a_12960_8860.t6 VGND 0.010076f
C274 a_12960_8860.n10 VGND 0.021345f
C275 a_12960_8860.t4 VGND 0.010076f
C276 a_12960_8860.t8 VGND 0.010076f
C277 a_12960_8860.n11 VGND 0.021345f
C278 a_12960_8860.t5 VGND 0.010076f
C279 a_12960_8860.t9 VGND 0.010076f
C280 a_12960_8860.n12 VGND 0.021345f
C281 a_12960_8860.t7 VGND 0.010076f
C282 a_12960_8860.t2 VGND 0.010076f
C283 a_12960_8860.n13 VGND 0.021345f
C284 a_12960_8860.n14 VGND 2.29634f
C285 a_12960_8860.n15 VGND 0.021345f
C286 a_12960_8860.t10 VGND 0.010076f
C287 a_13070_11250.n0 VGND 0.314325f
C288 a_13070_11250.n1 VGND 0.314325f
C289 a_13070_11250.n2 VGND 0.314325f
C290 a_13070_11250.n3 VGND 0.395925f
C291 a_13070_11250.n4 VGND 0.157163f
C292 a_13070_11250.n5 VGND 0.314325f
C293 a_13070_11250.n6 VGND 0.314325f
C294 a_13070_11250.n7 VGND 0.314325f
C295 a_13070_11250.n8 VGND 0.704522f
C296 a_13070_11250.n9 VGND 0.153679f
C297 a_13070_11250.n10 VGND 0.314325f
C298 a_13070_11250.n11 VGND 1.04942f
C299 a_13070_11250.n12 VGND 2.35472f
C300 a_13070_11250.n13 VGND 0.483896f
C301 a_13070_11250.t13 VGND 0.359229f
C302 a_13070_11250.t36 VGND 0.36519f
C303 a_13070_11250.t18 VGND 0.359229f
C304 a_13070_11250.t25 VGND 0.359229f
C305 a_13070_11250.t22 VGND 0.359229f
C306 a_13070_11250.t29 VGND 0.359229f
C307 a_13070_11250.t24 VGND 0.359229f
C308 a_13070_11250.t20 VGND 0.359229f
C309 a_13070_11250.t28 VGND 0.359229f
C310 a_13070_11250.t34 VGND 0.359229f
C311 a_13070_11250.t33 VGND 0.359229f
C312 a_13070_11250.t27 VGND 0.359229f
C313 a_13070_11250.t19 VGND 0.359229f
C314 a_13070_11250.t11 VGND 0.359229f
C315 a_13070_11250.t15 VGND 0.359229f
C316 a_13070_11250.t21 VGND 0.359229f
C317 a_13070_11250.t12 VGND 0.359229f
C318 a_13070_11250.t17 VGND 0.359229f
C319 a_13070_11250.t35 VGND 0.359229f
C320 a_13070_11250.t31 VGND 0.359229f
C321 a_13070_11250.t26 VGND 0.021589f
C322 a_13070_11250.t16 VGND 0.021247f
C323 a_13070_11250.n14 VGND 0.019024f
C324 a_13070_11250.t23 VGND 0.013904f
C325 a_13070_11250.t30 VGND 0.013904f
C326 a_13070_11250.n15 VGND 0.026482f
C327 a_13070_11250.n16 VGND 0.019024f
C328 a_13070_11250.t6 VGND 0.015816f
C329 a_13070_11250.n17 VGND 0.011348f
C330 a_13070_11250.n18 VGND 0.010949f
C331 a_13070_11250.n19 VGND 0.292028f
C332 a_13070_11250.t14 VGND 0.013904f
C333 a_13070_11250.t32 VGND 0.013904f
C334 a_13070_11250.n20 VGND 0.025867f
C335 a_13070_11250.n21 VGND 0.019024f
C336 a_10000_15820.t2 VGND 0.051177f
C337 a_10000_15820.t4 VGND 0.051177f
C338 a_10000_15820.n0 VGND 0.127304f
C339 a_10000_15820.t3 VGND 0.051177f
C340 a_10000_15820.t1 VGND 0.051177f
C341 a_10000_15820.n1 VGND 0.122338f
C342 a_10000_15820.n2 VGND 1.74488f
C343 a_10000_15820.t6 VGND 0.026228f
C344 a_10000_15820.t9 VGND 0.026176f
C345 a_10000_15820.n3 VGND 0.184117f
C346 a_10000_15820.t7 VGND 0.026176f
C347 a_10000_15820.n4 VGND 0.114474f
C348 a_10000_15820.t8 VGND 0.026176f
C349 a_10000_15820.n5 VGND 0.114474f
C350 a_10000_15820.t10 VGND 0.026176f
C351 a_10000_15820.n6 VGND 0.383297f
C352 a_10000_15820.n7 VGND 0.903315f
C353 a_10000_15820.t5 VGND 0.148895f
C354 a_10000_15820.n8 VGND 2.17873f
C355 a_10000_15820.t0 VGND 0.342532f
C356 a_13200_10990.n0 VGND 0.019256f
C357 a_13200_10990.t16 VGND 0.034183f
C358 a_13200_10990.n1 VGND 0.021429f
C359 a_13200_10990.n2 VGND 0.554666f
C360 a_13200_10990.n3 VGND 0.186578f
C361 a_13200_10990.t8 VGND 0.027505f
C362 a_13200_10990.t4 VGND 0.021667f
C363 a_13200_10990.t17 VGND 0.021667f
C364 a_13200_10990.t20 VGND 0.034973f
C365 a_13200_10990.n4 VGND 0.039055f
C366 a_13200_10990.n5 VGND 0.02668f
C367 a_13200_10990.n6 VGND 0.043175f
C368 a_13200_10990.t9 VGND 0.018056f
C369 a_13200_10990.t5 VGND 0.018056f
C370 a_13200_10990.n7 VGND 0.036969f
C371 a_13200_10990.n8 VGND 0.191386f
C372 a_13200_10990.t6 VGND 0.027505f
C373 a_13200_10990.t0 VGND 0.021667f
C374 a_13200_10990.t19 VGND 0.021667f
C375 a_13200_10990.t22 VGND 0.034973f
C376 a_13200_10990.n9 VGND 0.039055f
C377 a_13200_10990.n10 VGND 0.02668f
C378 a_13200_10990.n11 VGND 0.043175f
C379 a_13200_10990.t7 VGND 0.018056f
C380 a_13200_10990.t1 VGND 0.018056f
C381 a_13200_10990.n12 VGND 0.036969f
C382 a_13200_10990.n13 VGND 0.191386f
C383 a_13200_10990.n14 VGND 0.26218f
C384 a_13200_10990.t10 VGND 0.027505f
C385 a_13200_10990.t2 VGND 0.021667f
C386 a_13200_10990.t18 VGND 0.021667f
C387 a_13200_10990.t21 VGND 0.034973f
C388 a_13200_10990.n15 VGND 0.039055f
C389 a_13200_10990.n16 VGND 0.02668f
C390 a_13200_10990.n17 VGND 0.043175f
C391 a_13200_10990.n18 VGND 0.239421f
C392 a_13200_10990.t3 VGND 0.018056f
C393 a_13200_10990.n19 VGND 0.036969f
C394 a_13200_10990.t11 VGND 0.018056f
C395 a_9450_17070.t8 VGND 0.44893f
C396 a_9450_17070.t20 VGND 0.473023f
C397 a_9450_17070.t4 VGND 0.473023f
C398 a_9450_17070.t18 VGND 0.473023f
C399 a_9450_17070.t7 VGND 0.473023f
C400 a_9450_17070.t5 VGND 0.473023f
C401 a_9450_17070.t16 VGND 0.473023f
C402 a_9450_17070.t15 VGND 0.473023f
C403 a_9450_17070.t12 VGND 0.450557f
C404 a_9450_17070.t1 VGND 0.217037f
C405 a_9450_17070.n0 VGND 0.279945f
C406 a_9450_17070.t0 VGND 0.492104f
C407 a_9450_17070.t14 VGND 0.45245f
C408 a_9450_17070.t9 VGND 0.473023f
C409 a_9450_17070.t17 VGND 0.473023f
C410 a_9450_17070.t2 VGND 0.473023f
C411 a_9450_17070.t10 VGND 0.473023f
C412 a_9450_17070.t19 VGND 0.473023f
C413 a_9450_17070.t3 VGND 0.473023f
C414 a_9450_17070.t11 VGND 0.473023f
C415 a_9450_17070.t13 VGND 1.73608f
C416 a_9450_17070.t6 VGND 0.300567f
C417 a_10480_13480.t7 VGND 0.016248f
C418 a_10480_13480.t6 VGND 0.016248f
C419 a_10480_13480.n0 VGND 0.053414f
C420 a_10480_13480.t0 VGND 1.72364f
C421 a_10480_13480.t1 VGND 0.04531f
C422 a_10480_13480.n1 VGND 1.47476f
C423 a_10480_13480.t3 VGND 0.04324f
C424 a_10480_13480.t4 VGND 0.04324f
C425 a_10480_13480.n2 VGND 0.106515f
C426 a_10480_13480.n3 VGND 2.1672f
C427 a_10480_13480.n4 VGND 1.2172f
C428 a_10480_13480.t2 VGND 0.04324f
C429 a_10480_13480.n5 VGND 0.106515f
C430 a_10480_13480.t5 VGND 0.04324f
C431 a_9450_16252.t11 VGND 0.049701f
C432 a_9450_16252.t17 VGND 0.049641f
C433 a_9450_16252.n0 VGND 0.259634f
C434 a_9450_16252.t28 VGND 0.049641f
C435 a_9450_16252.n1 VGND 0.136128f
C436 a_9450_16252.t20 VGND 0.049641f
C437 a_9450_16252.n2 VGND 0.136128f
C438 a_9450_16252.t13 VGND 0.049641f
C439 a_9450_16252.n3 VGND 0.136128f
C440 a_9450_16252.t23 VGND 0.049641f
C441 a_9450_16252.n4 VGND 0.136128f
C442 a_9450_16252.t15 VGND 0.049641f
C443 a_9450_16252.n5 VGND 0.136128f
C444 a_9450_16252.t26 VGND 0.049641f
C445 a_9450_16252.n6 VGND 0.136128f
C446 a_9450_16252.t19 VGND 0.049641f
C447 a_9450_16252.n7 VGND 0.136128f
C448 a_9450_16252.t29 VGND 0.049641f
C449 a_9450_16252.n8 VGND 0.337114f
C450 a_9450_16252.t10 VGND 0.049641f
C451 a_9450_16252.n9 VGND 0.337114f
C452 a_9450_16252.t21 VGND 0.049641f
C453 a_9450_16252.n10 VGND 0.136128f
C454 a_9450_16252.t25 VGND 0.049641f
C455 a_9450_16252.n11 VGND 0.136128f
C456 a_9450_16252.t18 VGND 0.049641f
C457 a_9450_16252.n12 VGND 0.136128f
C458 a_9450_16252.t12 VGND 0.049641f
C459 a_9450_16252.n13 VGND 0.136128f
C460 a_9450_16252.t22 VGND 0.049641f
C461 a_9450_16252.n14 VGND 0.136128f
C462 a_9450_16252.t14 VGND 0.049641f
C463 a_9450_16252.n15 VGND 0.136128f
C464 a_9450_16252.t24 VGND 0.049641f
C465 a_9450_16252.n16 VGND 0.136128f
C466 a_9450_16252.t16 VGND 0.049641f
C467 a_9450_16252.n17 VGND 0.136128f
C468 a_9450_16252.t27 VGND 0.049641f
C469 a_9450_16252.n18 VGND 0.992373f
C470 a_9450_16252.t6 VGND 0.43431f
C471 a_9450_16252.t5 VGND 0.028712f
C472 a_9450_16252.t9 VGND 0.028712f
C473 a_9450_16252.n19 VGND 0.062021f
C474 a_9450_16252.n20 VGND 1.41734f
C475 a_9450_16252.t0 VGND 0.028712f
C476 a_9450_16252.t7 VGND 0.028712f
C477 a_9450_16252.n21 VGND 0.062021f
C478 a_9450_16252.n22 VGND 0.627074f
C479 a_9450_16252.t8 VGND 0.028712f
C480 a_9450_16252.t3 VGND 0.028712f
C481 a_9450_16252.n23 VGND 0.062021f
C482 a_9450_16252.n24 VGND 0.614154f
C483 a_9450_16252.t1 VGND 0.028712f
C484 a_9450_16252.t4 VGND 0.028712f
C485 a_9450_16252.n25 VGND 0.062021f
C486 a_9450_16252.n26 VGND 0.715576f
C487 a_9450_16252.n27 VGND 4.11339f
C488 a_9450_16252.t2 VGND 0.439339f
C489 a_9570_16200.t5 VGND 0.10095f
C490 a_9570_16200.t2 VGND 0.10095f
C491 a_9570_16200.n0 VGND 0.281599f
C492 a_9570_16200.t0 VGND 0.10095f
C493 a_9570_16200.t1 VGND 0.10095f
C494 a_9570_16200.n1 VGND 0.253459f
C495 a_9570_16200.n2 VGND 3.1126f
C496 a_9570_16200.t3 VGND 0.10095f
C497 a_9570_16200.t4 VGND 0.10095f
C498 a_9570_16200.n3 VGND 0.253459f
C499 a_9570_16200.n4 VGND 2.34993f
C500 a_9570_16200.t10 VGND 0.055705f
C501 a_9570_16200.t7 VGND 0.05457f
C502 a_9570_16200.n5 VGND 0.425181f
C503 a_9570_16200.t9 VGND 0.05457f
C504 a_9570_16200.n6 VGND 0.226997f
C505 a_9570_16200.t8 VGND 0.055305f
C506 a_9570_16200.n7 VGND 0.228617f
C507 a_9570_16200.t11 VGND 0.055305f
C508 a_9570_16200.n8 VGND 0.780841f
C509 a_9570_16200.n9 VGND 4.03498f
C510 a_9570_16200.t6 VGND 0.471183f
C511 a_11200_9430.t10 VGND 0.175143f
C512 a_11200_9430.t46 VGND 0.176134f
C513 a_11200_9430.n0 VGND 0.078499f
C514 a_11200_9430.t20 VGND 0.176493f
C515 a_11200_9430.t16 VGND 0.177254f
C516 a_11200_9430.n1 VGND 0.223018f
C517 a_11200_9430.t47 VGND 0.177254f
C518 a_11200_9430.n2 VGND 0.122165f
C519 a_11200_9430.t45 VGND 0.177254f
C520 a_11200_9430.n3 VGND 0.122165f
C521 a_11200_9430.t41 VGND 0.177254f
C522 a_11200_9430.n4 VGND 0.122165f
C523 a_11200_9430.t26 VGND 0.177254f
C524 a_11200_9430.n5 VGND 0.122165f
C525 a_11200_9430.n6 VGND 0.034548f
C526 a_11200_9430.n7 VGND 0.023032f
C527 a_11200_9430.t15 VGND 0.175981f
C528 a_11200_9430.t28 VGND 0.177254f
C529 a_11200_9430.n8 VGND 0.22257f
C530 a_11200_9430.t32 VGND 0.177254f
C531 a_11200_9430.n9 VGND 0.122165f
C532 a_11200_9430.t36 VGND 0.177254f
C533 a_11200_9430.n10 VGND 0.122165f
C534 a_11200_9430.t42 VGND 0.177254f
C535 a_11200_9430.n11 VGND 0.122165f
C536 a_11200_9430.t21 VGND 0.177254f
C537 a_11200_9430.n12 VGND 0.122165f
C538 a_11200_9430.t33 VGND 0.177254f
C539 a_11200_9430.n13 VGND 0.122165f
C540 a_11200_9430.t37 VGND 0.175891f
C541 a_11200_9430.n14 VGND 0.115851f
C542 a_11200_9430.n15 VGND 0.034548f
C543 a_11200_9430.t44 VGND 0.174871f
C544 a_11200_9430.n16 VGND 0.072085f
C545 a_11200_9430.n17 VGND 0.122838f
C546 a_11200_9430.n18 VGND 0.479119f
C547 a_11200_9430.t13 VGND 0.012796f
C548 a_11200_9430.t8 VGND 0.012796f
C549 a_11200_9430.n19 VGND 0.02764f
C550 a_11200_9430.n20 VGND 0.260499f
C551 a_11200_9430.t4 VGND 0.012796f
C552 a_11200_9430.t3 VGND 0.012796f
C553 a_11200_9430.n21 VGND 0.02764f
C554 a_11200_9430.n22 VGND 0.279456f
C555 a_11200_9430.t5 VGND 0.012796f
C556 a_11200_9430.t1 VGND 0.012796f
C557 a_11200_9430.n23 VGND 0.02764f
C558 a_11200_9430.n24 VGND 0.271779f
C559 a_11200_9430.t6 VGND 0.012796f
C560 a_11200_9430.t0 VGND 0.012796f
C561 a_11200_9430.n25 VGND 0.026199f
C562 a_11200_9430.t11 VGND 0.012796f
C563 a_11200_9430.t7 VGND 0.012796f
C564 a_11200_9430.n26 VGND 0.029778f
C565 a_11200_9430.t9 VGND 0.012796f
C566 a_11200_9430.t12 VGND 0.012796f
C567 a_11200_9430.n27 VGND 0.026199f
C568 a_11200_9430.n28 VGND 0.350925f
C569 a_11200_9430.n29 VGND 0.216918f
C570 a_11200_9430.n30 VGND 0.657119f
C571 a_11200_9430.t22 VGND 0.511827f
C572 a_11200_9430.t17 VGND 0.520321f
C573 a_11200_9430.t25 VGND 0.511827f
C574 a_11200_9430.n31 VGND 0.340188f
C575 a_11200_9430.t35 VGND 0.511827f
C576 a_11200_9430.n32 VGND 0.223924f
C577 a_11200_9430.t31 VGND 0.511827f
C578 a_11200_9430.n33 VGND 0.223924f
C579 a_11200_9430.t40 VGND 0.511827f
C580 a_11200_9430.n34 VGND 0.223924f
C581 a_11200_9430.t34 VGND 0.511827f
C582 a_11200_9430.n35 VGND 0.223924f
C583 a_11200_9430.t29 VGND 0.511827f
C584 a_11200_9430.n36 VGND 0.223924f
C585 a_11200_9430.t39 VGND 0.511827f
C586 a_11200_9430.n37 VGND 0.223924f
C587 a_11200_9430.t49 VGND 0.511827f
C588 a_11200_9430.n38 VGND 0.223924f
C589 a_11200_9430.n39 VGND 0.223924f
C590 a_11200_9430.t48 VGND 0.511827f
C591 a_11200_9430.n40 VGND 0.223924f
C592 a_11200_9430.t38 VGND 0.511827f
C593 a_11200_9430.n41 VGND 0.223924f
C594 a_11200_9430.t27 VGND 0.511827f
C595 a_11200_9430.n42 VGND 0.223924f
C596 a_11200_9430.t18 VGND 0.511827f
C597 a_11200_9430.n43 VGND 0.223924f
C598 a_11200_9430.t23 VGND 0.511827f
C599 a_11200_9430.n44 VGND 0.223924f
C600 a_11200_9430.t30 VGND 0.511827f
C601 a_11200_9430.n45 VGND 0.223924f
C602 a_11200_9430.t19 VGND 0.511827f
C603 a_11200_9430.n46 VGND 0.223924f
C604 a_11200_9430.t24 VGND 0.511827f
C605 a_11200_9430.n47 VGND 0.223924f
C606 a_11200_9430.t14 VGND 0.511827f
C607 a_11200_9430.n48 VGND 0.222325f
C608 a_11200_9430.t43 VGND 0.511827f
C609 a_11200_9430.n49 VGND 0.39273f
C610 a_11200_9430.n50 VGND 1.20725f
C611 a_11200_9430.t2 VGND 0.144453f
C612 VDPWR.n1 VGND 0.047692f
C613 VDPWR.t367 VGND 0.02994f
C614 VDPWR.n3 VGND 0.03643f
C615 VDPWR.t63 VGND 0.023876f
C616 VDPWR.n5 VGND 0.03643f
C617 VDPWR.t176 VGND 0.028803f
C618 VDPWR.t113 VGND 0.027287f
C619 VDPWR.t0 VGND 0.027287f
C620 VDPWR.t380 VGND 0.023876f
C621 VDPWR.n8 VGND 0.065328f
C622 VDPWR.n10 VGND 0.043938f
C623 VDPWR.n11 VGND 0.036559f
C624 VDPWR.n13 VGND 0.022922f
C625 VDPWR.t399 VGND 0.047373f
C626 VDPWR.t242 VGND 0.045479f
C627 VDPWR.t322 VGND 0.027287f
C628 VDPWR.t201 VGND 0.027287f
C629 VDPWR.t80 VGND 0.023876f
C630 VDPWR.t157 VGND 0.027287f
C631 VDPWR.t65 VGND 0.027287f
C632 VDPWR.t337 VGND 0.045479f
C633 VDPWR.t214 VGND 0.047373f
C634 VDPWR.n14 VGND 0.022922f
C635 VDPWR.n16 VGND 0.036559f
C636 VDPWR.n18 VGND 0.043938f
C637 VDPWR.n20 VGND 0.03643f
C638 VDPWR.n22 VGND 0.043938f
C639 VDPWR.n23 VGND 0.036559f
C640 VDPWR.n25 VGND 0.022922f
C641 VDPWR.t167 VGND 0.047373f
C642 VDPWR.t371 VGND 0.045479f
C643 VDPWR.t209 VGND 0.027287f
C644 VDPWR.t72 VGND 0.027287f
C645 VDPWR.t216 VGND 0.023876f
C646 VDPWR.t407 VGND 0.034109f
C647 VDPWR.t61 VGND 0.034109f
C648 VDPWR.t182 VGND 0.027287f
C649 VDPWR.t409 VGND 0.027287f
C650 VDPWR.t395 VGND 0.043963f
C651 VDPWR.t351 VGND 0.043963f
C652 VDPWR.t36 VGND 0.033351f
C653 VDPWR.t169 VGND 0.033351f
C654 VDPWR.t384 VGND 0.046994f
C655 VDPWR.t161 VGND 0.048889f
C656 VDPWR.n26 VGND 0.022922f
C657 VDPWR.n28 VGND 0.037136f
C658 VDPWR.n30 VGND 0.046825f
C659 VDPWR.n32 VGND 0.042494f
C660 VDPWR.n33 VGND 0.03669f
C661 VDPWR.n34 VGND 0.030337f
C662 VDPWR.n36 VGND 0.036141f
C663 VDPWR.n38 VGND 0.041339f
C664 VDPWR.n40 VGND 0.052023f
C665 VDPWR.n42 VGND 0.053694f
C666 VDPWR.n43 VGND 0.042334f
C667 VDPWR.n45 VGND 0.028986f
C668 VDPWR.t125 VGND 0.057227f
C669 VDPWR.t74 VGND 0.055332f
C670 VDPWR.t149 VGND 0.016675f
C671 VDPWR.t71 VGND 0.033351f
C672 VDPWR.t14 VGND 0.033351f
C673 VDPWR.t89 VGND 0.050784f
C674 VDPWR.t153 VGND 0.050784f
C675 VDPWR.t369 VGND 0.02994f
C676 VDPWR.t244 VGND 0.065565f
C677 VDPWR.n46 VGND 0.028986f
C678 VDPWR.n48 VGND 0.591495f
C679 VDPWR.n49 VGND 0.016597f
C680 VDPWR.n50 VGND 0.074071f
C681 VDPWR.n51 VGND 0.016184f
C682 VDPWR.n52 VGND 0.012994f
C683 VDPWR.n53 VGND 0.021656f
C684 VDPWR.t279 VGND 0.090018f
C685 VDPWR.t278 VGND 0.033953f
C686 VDPWR.t310 VGND 0.033953f
C687 VDPWR.n57 VGND 0.015296f
C688 VDPWR.n58 VGND 0.038146f
C689 VDPWR.n59 VGND 0.021656f
C690 VDPWR.n60 VGND 0.020213f
C691 VDPWR.t313 VGND 0.036285f
C692 VDPWR.n62 VGND 0.022954f
C693 VDPWR.n64 VGND 0.011695f
C694 VDPWR.n66 VGND 0.012994f
C695 VDPWR.n70 VGND 0.016184f
C696 VDPWR.n71 VGND 0.012994f
C697 VDPWR.t361 VGND 0.092112f
C698 VDPWR.t155 VGND 0.092112f
C699 VDPWR.t138 VGND 0.092112f
C700 VDPWR.t117 VGND 0.092112f
C701 VDPWR.t314 VGND 0.090018f
C702 VDPWR.n74 VGND 0.081645f
C703 VDPWR.n76 VGND 0.01178f
C704 VDPWR.n77 VGND 0.021656f
C705 VDPWR.t315 VGND 0.014438f
C706 VDPWR.n78 VGND 0.016597f
C707 VDPWR.n79 VGND 0.082328f
C708 VDPWR.n80 VGND 0.016597f
C709 VDPWR.n81 VGND 0.080424f
C710 VDPWR.n82 VGND 0.016597f
C711 VDPWR.n83 VGND 0.076959f
C712 VDPWR.n86 VGND 0.020213f
C713 VDPWR.n87 VGND 0.020213f
C714 VDPWR.n88 VGND 0.019612f
C715 VDPWR.n89 VGND 0.030929f
C716 VDPWR.n90 VGND 0.019025f
C717 VDPWR.n91 VGND 0.016597f
C718 VDPWR.n92 VGND 0.080424f
C719 VDPWR.n93 VGND 0.076959f
C720 VDPWR.n94 VGND 0.016597f
C721 VDPWR.t312 VGND 0.014438f
C722 VDPWR.n95 VGND 0.021656f
C723 VDPWR.n97 VGND 0.026324f
C724 VDPWR.n99 VGND 0.087925f
C725 VDPWR.t311 VGND 0.090018f
C726 VDPWR.t382 VGND 0.092112f
C727 VDPWR.t339 VGND 0.092112f
C728 VDPWR.t341 VGND 0.092112f
C729 VDPWR.t123 VGND 0.092112f
C730 VDPWR.t290 VGND 0.090018f
C731 VDPWR.n102 VGND 0.012994f
C732 VDPWR.n104 VGND 0.013201f
C733 VDPWR.n106 VGND 0.081645f
C734 VDPWR.n108 VGND 0.013115f
C735 VDPWR.t289 VGND 0.036285f
C736 VDPWR.n110 VGND 0.022347f
C737 VDPWR.n111 VGND 0.027666f
C738 VDPWR.n112 VGND 0.030205f
C739 VDPWR.n117 VGND 0.091702f
C740 VDPWR.t331 VGND 0.015198f
C741 VDPWR.n122 VGND 0.023176f
C742 VDPWR.n123 VGND 0.030431f
C743 VDPWR.t199 VGND 0.015198f
C744 VDPWR.n133 VGND 0.091702f
C745 VDPWR.t329 VGND 0.015198f
C746 VDPWR.n138 VGND 0.023176f
C747 VDPWR.n139 VGND 0.030431f
C748 VDPWR.t235 VGND 0.015198f
C749 VDPWR.n145 VGND 0.011394f
C750 VDPWR.n146 VGND 0.010251f
C751 VDPWR.n147 VGND 0.063671f
C752 VDPWR.n148 VGND 0.03861f
C753 VDPWR.n149 VGND 0.063671f
C754 VDPWR.n150 VGND 0.138944f
C755 VDPWR.n151 VGND 0.042224f
C756 VDPWR.n153 VGND 0.016854f
C757 VDPWR.n158 VGND 0.091702f
C758 VDPWR.t327 VGND 0.015198f
C759 VDPWR.n163 VGND 0.023176f
C760 VDPWR.n164 VGND 0.030431f
C761 VDPWR.t250 VGND 0.015198f
C762 VDPWR.n170 VGND 0.011394f
C763 VDPWR.n171 VGND 0.045104f
C764 VDPWR.t23 VGND 0.015561f
C765 VDPWR.n172 VGND 0.055444f
C766 VDPWR.n174 VGND 0.012135f
C767 VDPWR.n175 VGND 0.0251f
C768 VDPWR.n176 VGND 0.249108f
C769 VDPWR.t22 VGND 0.49577f
C770 VDPWR.t249 VGND 0.43737f
C771 VDPWR.t238 VGND 0.186967f
C772 VDPWR.n177 VGND 0.25708f
C773 VDPWR.t234 VGND 0.250402f
C774 VDPWR.t328 VGND 0.347225f
C775 VDPWR.t198 VGND 0.347225f
C776 VDPWR.t330 VGND 0.264449f
C777 VDPWR.n178 VGND 0.195486f
C778 VDPWR.n179 VGND 0.047337f
C779 VDPWR.n180 VGND 0.026219f
C780 VDPWR.n181 VGND 0.011394f
C781 VDPWR.n182 VGND 0.118274f
C782 VDPWR.n183 VGND 2.33098f
C783 VDPWR.n184 VGND 0.029101f
C784 VDPWR.n185 VGND 0.014367f
C785 VDPWR.t377 VGND 0.109654f
C786 VDPWR.n193 VGND 0.015881f
C787 VDPWR.n196 VGND 0.015881f
C788 VDPWR.n197 VGND 0.019008f
C789 VDPWR.n201 VGND 0.015881f
C790 VDPWR.t378 VGND 0.015233f
C791 VDPWR.n204 VGND 0.015832f
C792 VDPWR.n206 VGND 0.022436f
C793 VDPWR.n207 VGND 0.014367f
C794 VDPWR.n210 VGND 0.087275f
C795 VDPWR.n213 VGND 0.010106f
C796 VDPWR.t406 VGND 0.021451f
C797 VDPWR.n214 VGND 0.027059f
C798 VDPWR.n216 VGND 0.025347f
C799 VDPWR.t388 VGND 0.060421f
C800 VDPWR.t109 VGND 0.174551f
C801 VDPWR.n227 VGND 0.021656f
C802 VDPWR.n228 VGND 0.021656f
C803 VDPWR.n230 VGND 0.013115f
C804 VDPWR.n231 VGND 0.012994f
C805 VDPWR.n234 VGND 0.012994f
C806 VDPWR.n235 VGND 0.015415f
C807 VDPWR.n236 VGND 0.056644f
C808 VDPWR.n237 VGND 0.021656f
C809 VDPWR.n238 VGND 0.012994f
C810 VDPWR.t16 VGND 0.203643f
C811 VDPWR.n244 VGND 0.021656f
C812 VDPWR.n245 VGND 0.021656f
C813 VDPWR.n247 VGND 0.013115f
C814 VDPWR.n248 VGND 0.012994f
C815 VDPWR.n251 VGND 0.012994f
C816 VDPWR.n252 VGND 0.015415f
C817 VDPWR.n253 VGND 0.021656f
C818 VDPWR.n254 VGND 0.012994f
C819 VDPWR.t230 VGND 0.212594f
C820 VDPWR.n259 VGND 0.012994f
C821 VDPWR.n260 VGND 0.011695f
C822 VDPWR.t200 VGND 0.230497f
C823 VDPWR.n262 VGND 0.174551f
C824 VDPWR.n264 VGND 0.016045f
C825 VDPWR.n265 VGND 0.059112f
C826 VDPWR.n266 VGND 0.010189f
C827 VDPWR.n267 VGND 0.015415f
C828 VDPWR.n269 VGND 0.012994f
C829 VDPWR.n271 VGND 0.012994f
C830 VDPWR.n272 VGND 0.013115f
C831 VDPWR.n274 VGND 0.174551f
C832 VDPWR.t190 VGND 0.174551f
C833 VDPWR.n275 VGND 0.013115f
C834 VDPWR.n277 VGND 0.012994f
C835 VDPWR.n280 VGND 0.174551f
C836 VDPWR.n282 VGND 0.016999f
C837 VDPWR.n283 VGND 0.027012f
C838 VDPWR.n284 VGND 0.02708f
C839 VDPWR.n285 VGND 0.010189f
C840 VDPWR.n286 VGND 0.015415f
C841 VDPWR.n288 VGND 0.012994f
C842 VDPWR.n290 VGND 0.012994f
C843 VDPWR.n291 VGND 0.013115f
C844 VDPWR.n293 VGND 0.190216f
C845 VDPWR.t246 VGND 0.060421f
C846 VDPWR.n295 VGND 0.010106f
C847 VDPWR.n296 VGND 0.010106f
C848 VDPWR.t389 VGND 0.015226f
C849 VDPWR.n297 VGND 0.014061f
C850 VDPWR.n299 VGND 0.123081f
C851 VDPWR.n301 VGND 0.014367f
C852 VDPWR.n302 VGND 0.010253f
C853 VDPWR.n303 VGND 0.010106f
C854 VDPWR.n305 VGND 0.010106f
C855 VDPWR.n306 VGND 0.014061f
C856 VDPWR.t247 VGND 0.015226f
C857 VDPWR.n308 VGND 0.014367f
C858 VDPWR.n310 VGND 0.087275f
C859 VDPWR.t115 VGND 0.060421f
C860 VDPWR.t24 VGND 0.060421f
C861 VDPWR.n312 VGND 0.010106f
C862 VDPWR.n313 VGND 0.010106f
C863 VDPWR.t116 VGND 0.015226f
C864 VDPWR.n314 VGND 0.014061f
C865 VDPWR.n316 VGND 0.087275f
C866 VDPWR.n318 VGND 0.014367f
C867 VDPWR.t25 VGND 0.015226f
C868 VDPWR.n322 VGND 0.014061f
C869 VDPWR.n323 VGND 0.010106f
C870 VDPWR.n324 VGND 0.010106f
C871 VDPWR.n327 VGND 0.014367f
C872 VDPWR.n328 VGND 0.010253f
C873 VDPWR.n329 VGND 0.018706f
C874 VDPWR.n334 VGND 0.014213f
C875 VDPWR.n336 VGND 0.010106f
C876 VDPWR.t130 VGND 0.015226f
C877 VDPWR.n338 VGND 0.014061f
C878 VDPWR.n340 VGND 0.087275f
C879 VDPWR.t405 VGND 0.055946f
C880 VDPWR.t334 VGND 0.053708f
C881 VDPWR.t129 VGND 0.060421f
C882 VDPWR.n343 VGND 0.010106f
C883 VDPWR.n345 VGND 0.010106f
C884 VDPWR.n346 VGND 0.014061f
C885 VDPWR.t335 VGND 0.015151f
C886 VDPWR.n348 VGND 0.015671f
C887 VDPWR.n350 VGND 0.118605f
C888 VDPWR.t175 VGND 0.232734f
C889 VDPWR.t2 VGND 0.232734f
C890 VDPWR.t34 VGND 0.109654f
C891 VDPWR.t35 VGND 0.015226f
C892 VDPWR.n352 VGND 0.014061f
C893 VDPWR.n353 VGND 0.010106f
C894 VDPWR.n354 VGND 0.010106f
C895 VDPWR.n358 VGND 0.010106f
C896 VDPWR.n360 VGND 0.010106f
C897 VDPWR.t394 VGND 0.015226f
C898 VDPWR.n362 VGND 0.014061f
C899 VDPWR.n364 VGND 0.123081f
C900 VDPWR.n366 VGND 0.014367f
C901 VDPWR.n367 VGND 0.010253f
C902 VDPWR.n368 VGND 0.0317f
C903 VDPWR.n369 VGND 0.029101f
C904 VDPWR.n372 VGND 0.015832f
C905 VDPWR.n375 VGND 0.015881f
C906 VDPWR.t411 VGND 0.015233f
C907 VDPWR.n378 VGND 0.019008f
C908 VDPWR.n380 VGND 0.120843f
C909 VDPWR.t151 VGND 0.109654f
C910 VDPWR.t379 VGND 0.232734f
C911 VDPWR.t55 VGND 0.232734f
C912 VDPWR.t69 VGND 0.109654f
C913 VDPWR.t140 VGND 0.015226f
C914 VDPWR.n382 VGND 0.014061f
C915 VDPWR.n383 VGND 0.010106f
C916 VDPWR.n384 VGND 0.010106f
C917 VDPWR.n388 VGND 0.010106f
C918 VDPWR.n390 VGND 0.010106f
C919 VDPWR.t70 VGND 0.015226f
C920 VDPWR.n392 VGND 0.014061f
C921 VDPWR.n394 VGND 0.132032f
C922 VDPWR.n396 VGND 0.014367f
C923 VDPWR.n397 VGND 0.010253f
C924 VDPWR.n398 VGND 0.660617f
C925 VDPWR.t88 VGND 0.161413f
C926 VDPWR.t211 VGND 0.170075f
C927 VDPWR.t207 VGND 0.170075f
C928 VDPWR.t360 VGND 0.170075f
C929 VDPWR.t392 VGND 0.170075f
C930 VDPWR.t79 VGND 0.170075f
C931 VDPWR.t359 VGND 0.170075f
C932 VDPWR.t241 VGND 0.170075f
C933 VDPWR.t107 VGND 0.161998f
C934 VDPWR.t47 VGND 0.078035f
C935 VDPWR.n399 VGND 0.100654f
C936 VDPWR.t78 VGND 0.176936f
C937 VDPWR.t48 VGND 0.162678f
C938 VDPWR.t108 VGND 0.170075f
C939 VDPWR.t46 VGND 0.170075f
C940 VDPWR.t373 VGND 0.170075f
C941 VDPWR.t414 VGND 0.170075f
C942 VDPWR.t393 VGND 0.170075f
C943 VDPWR.t374 VGND 0.170075f
C944 VDPWR.t208 VGND 0.170075f
C945 VDPWR.t133 VGND 0.273581f
C946 VDPWR.t423 VGND 0.34111f
C947 VDPWR.t424 VGND 0.34111f
C948 VDPWR.t425 VGND 0.324071f
C949 VDPWR.n400 VGND 0.627227f
C950 VDPWR.n401 VGND 0.331175f
C951 VDPWR.t429 VGND 0.320121f
C952 VDPWR.n402 VGND 0.485349f
C953 VDPWR.n403 VGND 0.451194f
C954 VDPWR.n404 VGND 0.021362f
C955 VDPWR.n405 VGND 0.085621f
C956 VDPWR.n406 VGND 0.010887f
C957 VDPWR.t99 VGND 0.078017f
C958 VDPWR.n413 VGND 0.090075f
C959 VDPWR.n417 VGND 0.02707f
C960 VDPWR.n418 VGND 0.012994f
C961 VDPWR.t283 VGND 0.139485f
C962 VDPWR.t390 VGND 0.122936f
C963 VDPWR.t159 VGND 0.122936f
C964 VDPWR.t6 VGND 0.122936f
C965 VDPWR.t49 VGND 0.122936f
C966 VDPWR.t273 VGND 0.243002f
C967 VDPWR.t274 VGND 0.016553f
C968 VDPWR.n423 VGND 0.099215f
C969 VDPWR.n425 VGND 0.01561f
C970 VDPWR.t285 VGND 0.012937f
C971 VDPWR.n427 VGND 0.027153f
C972 VDPWR.n429 VGND 0.01561f
C973 VDPWR.n430 VGND 0.022592f
C974 VDPWR.n431 VGND 0.021362f
C975 VDPWR.n432 VGND 0.091396f
C976 VDPWR.n433 VGND 0.021362f
C977 VDPWR.n434 VGND 0.091396f
C978 VDPWR.n435 VGND 0.018754f
C979 VDPWR.n436 VGND 0.070903f
C980 VDPWR.n437 VGND 0.01386f
C981 VDPWR.n438 VGND 0.01155f
C982 VDPWR.t259 VGND 0.018047f
C983 VDPWR.n439 VGND 0.021362f
C984 VDPWR.n440 VGND 0.083311f
C985 VDPWR.n441 VGND 0.05122f
C986 VDPWR.t257 VGND 0.036065f
C987 VDPWR.n442 VGND 0.026302f
C988 VDPWR.n444 VGND 0.013115f
C989 VDPWR.n446 VGND 0.012994f
C990 VDPWR.n449 VGND 0.012994f
C991 VDPWR.n450 VGND 0.016184f
C992 VDPWR.n452 VGND 0.01178f
C993 VDPWR.n454 VGND 0.075653f
C994 VDPWR.t307 VGND 0.078017f
C995 VDPWR.t218 VGND 0.078017f
C996 VDPWR.t103 VGND 0.061468f
C997 VDPWR.t232 VGND 0.094566f
C998 VDPWR.t91 VGND 0.061468f
C999 VDPWR.t386 VGND 0.073289f
C1000 VDPWR.t67 VGND 0.082746f
C1001 VDPWR.t95 VGND 0.061468f
C1002 VDPWR.t267 VGND 0.094566f
C1003 VDPWR.t258 VGND 0.078017f
C1004 VDPWR.n455 VGND 0.101911f
C1005 VDPWR.t268 VGND 0.016555f
C1006 VDPWR.n456 VGND 0.042644f
C1007 VDPWR.n458 VGND 0.025354f
C1008 VDPWR.n459 VGND 0.031106f
C1009 VDPWR.n460 VGND 0.025354f
C1010 VDPWR.t309 VGND 0.012941f
C1011 VDPWR.n462 VGND 0.037508f
C1012 VDPWR.n463 VGND 0.101902f
C1013 VDPWR.t97 VGND 0.127665f
C1014 VDPWR.t93 VGND 0.120572f
C1015 VDPWR.t82 VGND 0.087474f
C1016 VDPWR.t248 VGND 0.068561f
C1017 VDPWR.t105 VGND 0.061468f
C1018 VDPWR.t5 VGND 0.094566f
C1019 VDPWR.t101 VGND 0.061468f
C1020 VDPWR.t332 VGND 0.082746f
C1021 VDPWR.t333 VGND 0.073289f
C1022 VDPWR.t303 VGND 0.061468f
C1023 VDPWR.t83 VGND 0.094566f
C1024 VDPWR.n467 VGND 0.012994f
C1025 VDPWR.n468 VGND 0.016184f
C1026 VDPWR.n469 VGND 0.012994f
C1027 VDPWR.n470 VGND 0.012994f
C1028 VDPWR.n472 VGND 0.02707f
C1029 VDPWR.n473 VGND 0.013201f
C1030 VDPWR.n475 VGND 0.196225f
C1031 VDPWR.n477 VGND 0.014618f
C1032 VDPWR.t302 VGND 0.035758f
C1033 VDPWR.n478 VGND 0.017414f
C1034 VDPWR.n479 VGND 0.08701f
C1035 VDPWR.n480 VGND 0.18141f
C1036 VDPWR.n482 VGND 0.077192f
C1037 VDPWR.n483 VGND 0.011227f
C1038 VDPWR.n484 VGND 0.011142f
C1039 VDPWR.n486 VGND 0.077192f
C1040 VDPWR.n488 VGND 0.077192f
C1041 VDPWR.n490 VGND 0.077192f
C1042 VDPWR.n492 VGND 0.077192f
C1043 VDPWR.n494 VGND 0.077192f
C1044 VDPWR.n496 VGND 0.077192f
C1045 VDPWR.n498 VGND 0.077192f
C1046 VDPWR.n500 VGND 0.077192f
C1047 VDPWR.n502 VGND 0.077192f
C1048 VDPWR.n503 VGND 0.011227f
C1049 VDPWR.n504 VGND 0.011142f
C1050 VDPWR.n506 VGND 0.077192f
C1051 VDPWR.n508 VGND 0.077192f
C1052 VDPWR.n510 VGND 0.077192f
C1053 VDPWR.n512 VGND 0.077192f
C1054 VDPWR.n514 VGND 0.077192f
C1055 VDPWR.n516 VGND 0.077192f
C1056 VDPWR.n518 VGND 0.077192f
C1057 VDPWR.n520 VGND 0.105185f
C1058 VDPWR.n521 VGND 0.033758f
C1059 VDPWR.t277 VGND 0.010044f
C1060 VDPWR.n523 VGND 0.011227f
C1061 VDPWR.n524 VGND 0.035593f
C1062 VDPWR.t276 VGND 0.029966f
C1063 VDPWR.t180 VGND 0.024255f
C1064 VDPWR.t59 VGND 0.024255f
C1065 VDPWR.t127 VGND 0.024255f
C1066 VDPWR.t205 VGND 0.024255f
C1067 VDPWR.t12 VGND 0.024255f
C1068 VDPWR.t220 VGND 0.024255f
C1069 VDPWR.t343 VGND 0.024255f
C1070 VDPWR.t147 VGND 0.024255f
C1071 VDPWR.t178 VGND 0.024255f
C1072 VDPWR.t76 VGND 0.024255f
C1073 VDPWR.t357 VGND 0.024255f
C1074 VDPWR.t325 VGND 0.024255f
C1075 VDPWR.t10 VGND 0.024255f
C1076 VDPWR.t192 VGND 0.024255f
C1077 VDPWR.t403 VGND 0.024255f
C1078 VDPWR.t20 VGND 0.024255f
C1079 VDPWR.t196 VGND 0.024255f
C1080 VDPWR.t345 VGND 0.024255f
C1081 VDPWR.t320 VGND 0.036856f
C1082 VDPWR.n525 VGND 0.030725f
C1083 VDPWR.t321 VGND 0.010044f
C1084 VDPWR.n526 VGND 0.011142f
C1085 VDPWR.n528 VGND 0.02384f
C1086 VDPWR.n529 VGND 0.078471f
C1087 VDPWR.n530 VGND 0.078471f
C1088 VDPWR.n531 VGND 0.031789f
C1089 VDPWR.t262 VGND 0.010044f
C1090 VDPWR.n533 VGND 0.011227f
C1091 VDPWR.n534 VGND 0.037369f
C1092 VDPWR.t261 VGND 0.030212f
C1093 VDPWR.t421 VGND 0.024255f
C1094 VDPWR.t57 VGND 0.024255f
C1095 VDPWR.t236 VGND 0.024255f
C1096 VDPWR.t145 VGND 0.024255f
C1097 VDPWR.t3 VGND 0.024255f
C1098 VDPWR.t84 VGND 0.024255f
C1099 VDPWR.t184 VGND 0.024255f
C1100 VDPWR.t375 VGND 0.024255f
C1101 VDPWR.t111 VGND 0.024255f
C1102 VDPWR.t18 VGND 0.024255f
C1103 VDPWR.t188 VGND 0.024255f
C1104 VDPWR.t42 VGND 0.024255f
C1105 VDPWR.t186 VGND 0.024255f
C1106 VDPWR.t194 VGND 0.024255f
C1107 VDPWR.t412 VGND 0.024255f
C1108 VDPWR.t203 VGND 0.024255f
C1109 VDPWR.t401 VGND 0.024255f
C1110 VDPWR.t8 VGND 0.024255f
C1111 VDPWR.t252 VGND 0.036294f
C1112 VDPWR.n535 VGND 0.029265f
C1113 VDPWR.t253 VGND 0.010044f
C1114 VDPWR.n536 VGND 0.011142f
C1115 VDPWR.n538 VGND 0.02384f
C1116 VDPWR.n539 VGND 0.205043f
C1117 VDPWR.n540 VGND 0.234087f
C1118 VDPWR.t269 VGND 0.041307f
C1119 VDPWR.n541 VGND 0.015834f
C1120 VDPWR.n542 VGND 0.033705f
C1121 VDPWR.n543 VGND 0.033705f
C1122 VDPWR.n544 VGND 0.033705f
C1123 VDPWR.n545 VGND 0.033705f
C1124 VDPWR.n546 VGND 0.033705f
C1125 VDPWR.n547 VGND 0.033705f
C1126 VDPWR.n548 VGND 0.033705f
C1127 VDPWR.n549 VGND 0.033705f
C1128 VDPWR.n559 VGND 0.010046f
C1129 VDPWR.n560 VGND 0.010046f
C1130 VDPWR.n562 VGND 0.010106f
C1131 VDPWR.n564 VGND 0.011539f
C1132 VDPWR.n567 VGND 0.010106f
C1133 VDPWR.n570 VGND 0.010106f
C1134 VDPWR.n571 VGND 0.010106f
C1135 VDPWR.n573 VGND 0.010892f
C1136 VDPWR.n575 VGND 0.080995f
C1137 VDPWR.t270 VGND 0.085904f
C1138 VDPWR.t347 VGND 0.088358f
C1139 VDPWR.t131 VGND 0.088358f
C1140 VDPWR.t28 VGND 0.088358f
C1141 VDPWR.t32 VGND 0.088358f
C1142 VDPWR.t415 VGND 0.088358f
C1143 VDPWR.t239 VGND 0.088358f
C1144 VDPWR.t26 VGND 0.088358f
C1145 VDPWR.t30 VGND 0.088358f
C1146 VDPWR.t228 VGND 0.088358f
C1147 VDPWR.t121 VGND 0.088358f
C1148 VDPWR.t349 VGND 0.088358f
C1149 VDPWR.t86 VGND 0.088358f
C1150 VDPWR.t226 VGND 0.088358f
C1151 VDPWR.t119 VGND 0.088358f
C1152 VDPWR.t44 VGND 0.088358f
C1153 VDPWR.t212 VGND 0.088358f
C1154 VDPWR.t264 VGND 0.085904f
C1155 VDPWR.n580 VGND 0.010106f
C1156 VDPWR.n583 VGND 0.010106f
C1157 VDPWR.n584 VGND 0.010046f
C1158 VDPWR.n586 VGND 0.010106f
C1159 VDPWR.n587 VGND 0.010106f
C1160 VDPWR.n588 VGND 0.010046f
C1161 VDPWR.n590 VGND 0.012185f
C1162 VDPWR.n592 VGND 0.080995f
C1163 VDPWR.n594 VGND 0.011539f
C1164 VDPWR.t263 VGND 0.041307f
C1165 VDPWR.n595 VGND 0.016683f
C1166 VDPWR.n596 VGND 0.165081f
C1167 VDPWR.n597 VGND 0.115868f
C1168 VDPWR.n598 VGND 0.115868f
C1169 VDPWR.n599 VGND 0.115868f
C1170 VDPWR.n600 VGND 0.115868f
C1171 VDPWR.n601 VGND 0.115868f
C1172 VDPWR.n602 VGND 0.115868f
C1173 VDPWR.n603 VGND 0.115868f
C1174 VDPWR.n604 VGND 0.097705f
C1175 VDPWR.n605 VGND 0.096351f
C1176 VDPWR.n606 VGND 0.011227f
C1177 VDPWR.n607 VGND 0.011806f
C1178 VDPWR.n608 VGND 0.036746f
C1179 VDPWR.t256 VGND 0.011458f
C1180 VDPWR.n610 VGND 0.011892f
C1181 VDPWR.n611 VGND 0.036151f
C1182 VDPWR.t255 VGND 0.029408f
C1183 VDPWR.t397 VGND 0.022234f
C1184 VDPWR.t398 VGND 0.022234f
C1185 VDPWR.t297 VGND 0.034899f
C1186 VDPWR.n612 VGND 0.028639f
C1187 VDPWR.t298 VGND 0.010044f
C1188 VDPWR.n613 VGND 0.011142f
C1189 VDPWR.n615 VGND 0.02768f
C1190 VDPWR.n616 VGND 0.227073f
C1191 VDPWR.n617 VGND 0.229015f
C1192 VDPWR.n619 VGND 0.034188f
C1193 VDPWR.n620 VGND 0.011313f
C1194 VDPWR.n621 VGND 0.011142f
C1195 VDPWR.t318 VGND 0.010044f
C1196 VDPWR.n624 VGND 0.034188f
C1197 VDPWR.n626 VGND 0.034188f
C1198 VDPWR.n628 VGND 0.034188f
C1199 VDPWR.n630 VGND 0.034188f
C1200 VDPWR.n632 VGND 0.034188f
C1201 VDPWR.n633 VGND 0.011313f
C1202 VDPWR.n634 VGND 0.011142f
C1203 VDPWR.t301 VGND 0.010044f
C1204 VDPWR.n637 VGND 0.034188f
C1205 VDPWR.n639 VGND 0.034188f
C1206 VDPWR.n641 VGND 0.034188f
C1207 VDPWR.n643 VGND 0.042236f
C1208 VDPWR.n644 VGND 0.014318f
C1209 VDPWR.n645 VGND 0.019014f
C1210 VDPWR.n646 VGND 0.011313f
C1211 VDPWR.n647 VGND 0.035032f
C1212 VDPWR.t300 VGND 0.028506f
C1213 VDPWR.t419 VGND 0.022234f
C1214 VDPWR.t141 VGND 0.022234f
C1215 VDPWR.t222 VGND 0.022234f
C1216 VDPWR.t134 VGND 0.022234f
C1217 VDPWR.t38 VGND 0.022234f
C1218 VDPWR.t171 VGND 0.022234f
C1219 VDPWR.t163 VGND 0.022234f
C1220 VDPWR.t224 VGND 0.022234f
C1221 VDPWR.t365 VGND 0.022234f
C1222 VDPWR.t51 VGND 0.022234f
C1223 VDPWR.t294 VGND 0.034899f
C1224 VDPWR.n648 VGND 0.028639f
C1225 VDPWR.t295 VGND 0.010044f
C1226 VDPWR.n649 VGND 0.011142f
C1227 VDPWR.n650 VGND 0.019014f
C1228 VDPWR.n651 VGND 0.013703f
C1229 VDPWR.n652 VGND 0.0231f
C1230 VDPWR.n653 VGND 0.0231f
C1231 VDPWR.n654 VGND 0.013703f
C1232 VDPWR.n655 VGND 0.019014f
C1233 VDPWR.n656 VGND 0.011313f
C1234 VDPWR.n657 VGND 0.035032f
C1235 VDPWR.t317 VGND 0.028506f
C1236 VDPWR.t355 VGND 0.022234f
C1237 VDPWR.t165 VGND 0.022234f
C1238 VDPWR.t417 VGND 0.022234f
C1239 VDPWR.t136 VGND 0.022234f
C1240 VDPWR.t40 VGND 0.022234f
C1241 VDPWR.t173 VGND 0.022234f
C1242 VDPWR.t363 VGND 0.022234f
C1243 VDPWR.t353 VGND 0.022234f
C1244 VDPWR.t143 VGND 0.022234f
C1245 VDPWR.t53 VGND 0.022234f
C1246 VDPWR.t287 VGND 0.034899f
C1247 VDPWR.n658 VGND 0.028639f
C1248 VDPWR.t288 VGND 0.010044f
C1249 VDPWR.n659 VGND 0.011142f
C1250 VDPWR.n660 VGND 0.019014f
C1251 VDPWR.n661 VGND 0.013703f
C1252 VDPWR.n662 VGND 0.099092f
C1253 VDPWR.n663 VGND 2.38946f
C1254 VDPWR.n664 VGND 13.061701f
C1255 VDPWR.n665 VGND 1.8068f
C1256 VDPWR.n666 VGND 1.8741f
C1257 a_18160_10940.t11 VGND 0.021157f
C1258 a_18160_10940.t4 VGND 0.021157f
C1259 a_18160_10940.n0 VGND 0.0506f
C1260 a_18160_10940.t0 VGND 0.021157f
C1261 a_18160_10940.t12 VGND 0.021157f
C1262 a_18160_10940.n1 VGND 0.0506f
C1263 a_18160_10940.t10 VGND 0.021157f
C1264 a_18160_10940.n2 VGND 0.050792f
C1265 a_18160_10940.t2 VGND 0.109026f
C1266 a_18160_10940.t1 VGND 0.032027f
C1267 a_18160_10940.n3 VGND 0.178496f
C1268 a_18160_10940.n4 VGND 0.147792f
C1269 a_18160_10940.t6 VGND 0.052891f
C1270 a_18160_10940.t7 VGND 0.052891f
C1271 a_18160_10940.n5 VGND 0.109442f
C1272 a_18160_10940.t8 VGND 0.052891f
C1273 a_18160_10940.t9 VGND 0.052891f
C1274 a_18160_10940.n6 VGND 0.158354f
C1275 a_18160_10940.n7 VGND 1.17815f
C1276 a_18160_10940.n8 VGND 0.051715f
C1277 a_18160_10940.n9 VGND 0.149118f
C1278 a_18160_10940.n10 VGND 0.14861f
C1279 a_18160_10940.t3 VGND 0.032027f
C1280 a_18160_10940.n11 VGND 0.150205f
C1281 a_18160_10940.t5 VGND 0.085694f
C1282 a_17714_9374.t7 VGND 0.035769f
C1283 a_17714_9374.t8 VGND 0.070362f
C1284 a_17714_9374.n0 VGND 1.12772f
C1285 a_17714_9374.t0 VGND 0.098723f
C1286 a_17714_9374.t4 VGND 0.098723f
C1287 a_17714_9374.t2 VGND 0.098723f
C1288 a_17714_9374.t12 VGND 0.098723f
C1289 a_17714_9374.t11 VGND 0.135741f
C1290 a_17714_9374.n1 VGND 0.076013f
C1291 a_17714_9374.n2 VGND 0.05394f
C1292 a_17714_9374.t3 VGND 0.035769f
C1293 a_17714_9374.t5 VGND 0.035769f
C1294 a_17714_9374.n3 VGND 0.073951f
C1295 a_17714_9374.n4 VGND 0.268783f
C1296 a_17714_9374.n5 VGND 0.024234f
C1297 a_17714_9374.n6 VGND 0.05394f
C1298 a_17714_9374.n7 VGND 0.05394f
C1299 a_17714_9374.t6 VGND 0.098723f
C1300 a_17714_9374.t9 VGND 0.098723f
C1301 a_17714_9374.t10 VGND 0.135741f
C1302 a_17714_9374.n8 VGND 0.076013f
C1303 a_17714_9374.n9 VGND 0.05394f
C1304 a_17714_9374.n10 VGND 0.024234f
C1305 a_17714_9374.n11 VGND 0.262083f
C1306 a_17714_9374.n12 VGND 0.073951f
C1307 a_17714_9374.t1 VGND 0.035769f
C1308 a_11860_6640.t7 VGND 0.028262f
C1309 a_11860_6640.t8 VGND 0.064454f
C1310 a_11860_6640.n0 VGND 0.162805f
C1311 a_11860_6640.t3 VGND 0.029978f
C1312 a_11860_6640.t4 VGND 0.063823f
C1313 a_11860_6640.n1 VGND 0.09612f
C1314 a_11860_6640.t6 VGND 0.063823f
C1315 a_11860_6640.t5 VGND 0.092852f
C1316 a_11860_6640.n2 VGND 1.17335f
C1317 a_11860_6640.n3 VGND 0.254916f
C1318 a_11860_6640.t0 VGND 0.025787f
C1319 a_11860_6640.t2 VGND 0.025787f
C1320 a_11860_6640.n4 VGND 0.137692f
C1321 a_11860_6640.n5 VGND 0.244629f
C1322 a_11860_6640.t1 VGND 0.135725f
C1323 V_CONT.t5 VGND 7.3922f
C1324 V_CONT.t4 VGND 0.01223f
C1325 V_CONT.n7 VGND 0.625987f
C1326 V_CONT.n13 VGND 0.087506f
C1327 V_CONT.n14 VGND 0.348177f
C1328 V_CONT.n16 VGND 0.658859f
C1329 V_CONT.n18 VGND 0.071511f
C1330 V_CONT.n22 VGND 0.039942f
C1331 V_CONT.n23 VGND 0.045404f
C1332 V_CONT.n24 VGND 0.345356f
C1333 V_CONT.n25 VGND 0.017231f
C1334 V_CONT.n26 VGND 0.010717f
C1335 V_CONT.n27 VGND 0.01887f
.ends

