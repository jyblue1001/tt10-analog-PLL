magic
tech sky130A
timestamp 1756757267
<< metal1 >>
rect 5210 15755 5250 15760
rect 5210 15725 5215 15755
rect 5245 15725 5250 15755
rect 5210 13735 5250 15725
rect 5210 13705 5215 13735
rect 5245 13705 5250 13735
rect 5210 13700 5250 13705
rect 12150 15380 12350 15385
rect 12150 15350 12155 15380
rect 12185 15350 12195 15380
rect 12225 15350 12235 15380
rect 12265 15350 12275 15380
rect 12305 15350 12315 15380
rect 12345 15350 12350 15380
rect 12150 13465 12350 15350
rect 12110 13425 12350 13465
rect 12150 13290 12350 13425
rect 12150 13260 12155 13290
rect 12185 13260 12195 13290
rect 12225 13260 12235 13290
rect 12265 13260 12275 13290
rect 12305 13260 12315 13290
rect 12345 13260 12350 13290
rect 12150 12645 12350 13260
rect 12150 12615 12155 12645
rect 12185 12615 12195 12645
rect 12225 12615 12235 12645
rect 12265 12615 12275 12645
rect 12305 12615 12315 12645
rect 12345 12615 12350 12645
rect 12150 12605 12350 12615
rect 12150 12575 12155 12605
rect 12185 12575 12195 12605
rect 12225 12575 12235 12605
rect 12265 12575 12275 12605
rect 12305 12575 12315 12605
rect 12345 12575 12350 12605
rect 12150 12565 12350 12575
rect 12150 12535 12155 12565
rect 12185 12535 12195 12565
rect 12225 12535 12235 12565
rect 12265 12535 12275 12565
rect 12305 12535 12315 12565
rect 12345 12535 12350 12565
rect 12150 7300 12350 12535
rect 12150 7270 12155 7300
rect 12185 7270 12195 7300
rect 12225 7270 12235 7300
rect 12265 7270 12275 7300
rect 12305 7270 12315 7300
rect 12345 7270 12350 7300
rect 12150 7265 12350 7270
<< via1 >>
rect 5215 15725 5245 15755
rect 5215 13705 5245 13735
rect 12155 15350 12185 15380
rect 12195 15350 12225 15380
rect 12235 15350 12265 15380
rect 12275 15350 12305 15380
rect 12315 15350 12345 15380
rect 12155 13260 12185 13290
rect 12195 13260 12225 13290
rect 12235 13260 12265 13290
rect 12275 13260 12305 13290
rect 12315 13260 12345 13290
rect 12155 12615 12185 12645
rect 12195 12615 12225 12645
rect 12235 12615 12265 12645
rect 12275 12615 12305 12645
rect 12315 12615 12345 12645
rect 12155 12575 12185 12605
rect 12195 12575 12225 12605
rect 12235 12575 12265 12605
rect 12275 12575 12305 12605
rect 12315 12575 12345 12605
rect 12155 12535 12185 12565
rect 12195 12535 12225 12565
rect 12235 12535 12265 12565
rect 12275 12535 12305 12565
rect 12315 12535 12345 12565
rect 12155 7270 12185 7300
rect 12195 7270 12225 7300
rect 12235 7270 12265 7300
rect 12275 7270 12305 7300
rect 12315 7270 12345 7300
<< metal2 >>
rect 5210 15755 15265 15760
rect 5210 15725 5215 15755
rect 5245 15740 15265 15755
rect 5245 15725 15205 15740
rect 5210 15720 15205 15725
rect 15185 15700 15205 15720
rect 15245 15700 15265 15740
rect 15185 15680 15265 15700
rect 12150 15380 12350 15385
rect 12150 15350 12155 15380
rect 12185 15350 12195 15380
rect 12225 15350 12235 15380
rect 12265 15350 12275 15380
rect 12305 15350 12315 15380
rect 12345 15350 12350 15380
rect 11830 14980 13335 15000
rect 11830 14960 13275 14980
rect 13255 14940 13275 14960
rect 13315 14940 13335 14980
rect 13255 14920 13335 14940
rect 12150 13290 12350 13295
rect 12150 13260 12155 13290
rect 12185 13260 12195 13290
rect 12225 13260 12235 13290
rect 12265 13260 12275 13290
rect 12305 13260 12315 13290
rect 12345 13260 12350 13290
rect 12150 13255 12350 13260
rect 12150 12645 12350 12650
rect 12150 12615 12155 12645
rect 12185 12615 12195 12645
rect 12225 12615 12235 12645
rect 12265 12615 12275 12645
rect 12305 12615 12315 12645
rect 12345 12615 12350 12645
rect 12150 12605 12350 12615
rect 12150 12575 12155 12605
rect 12185 12575 12195 12605
rect 12225 12575 12235 12605
rect 12265 12575 12275 12605
rect 12305 12575 12315 12605
rect 12345 12575 12350 12605
rect 12150 12565 12350 12575
rect 12150 12535 12155 12565
rect 12185 12535 12195 12565
rect 12225 12535 12235 12565
rect 12265 12535 12275 12565
rect 12305 12535 12315 12565
rect 12345 12535 12350 12565
rect 12150 12530 12350 12535
rect 3890 7475 4905 7495
rect 3890 7445 3895 7475
rect 3925 7445 3940 7475
rect 3970 7445 3985 7475
rect 4015 7445 4905 7475
rect 3890 7425 4905 7445
rect 3890 7395 3895 7425
rect 3925 7395 3940 7425
rect 3970 7395 3985 7425
rect 4015 7395 4905 7425
rect 3890 7375 4905 7395
rect 12150 7300 12350 7305
rect 12150 7270 12155 7300
rect 12185 7270 12195 7300
rect 12225 7270 12235 7300
rect 12265 7270 12275 7300
rect 12305 7270 12315 7300
rect 12345 7270 12350 7300
rect 12150 7265 12350 7270
rect 3890 7150 4020 7155
rect 3890 7120 3895 7150
rect 3925 7120 3940 7150
rect 3970 7120 3985 7150
rect 4015 7120 4020 7150
rect 3890 7105 4020 7120
rect 3890 7075 3895 7105
rect 3925 7075 3940 7105
rect 3970 7075 3985 7105
rect 4015 7075 4020 7105
rect 3890 7060 4020 7075
rect 3890 7030 3895 7060
rect 3925 7030 3940 7060
rect 3970 7030 3985 7060
rect 4015 7030 4020 7060
rect 3890 7025 4020 7030
<< via2 >>
rect 15205 15700 15245 15740
rect 13275 14940 13315 14980
rect 3895 7445 3925 7475
rect 3940 7445 3970 7475
rect 3985 7445 4015 7475
rect 3895 7395 3925 7425
rect 3940 7395 3970 7425
rect 3985 7395 4015 7425
rect 3895 7120 3925 7150
rect 3940 7120 3970 7150
rect 3985 7120 4015 7150
rect 3895 7075 3925 7105
rect 3940 7075 3970 7105
rect 3985 7075 4015 7105
rect 3895 7030 3925 7060
rect 3940 7030 3970 7060
rect 3985 7030 4015 7060
<< metal3 >>
rect 15185 15740 15265 15760
rect 400 15690 4020 15705
rect 400 15650 405 15690
rect 445 15650 455 15690
rect 495 15650 505 15690
rect 545 15650 555 15690
rect 595 15650 4020 15690
rect 15185 15700 15205 15740
rect 15245 15700 15265 15740
rect 15185 15680 15265 15700
rect 400 15640 4020 15650
rect 400 15600 405 15640
rect 445 15600 455 15640
rect 495 15600 505 15640
rect 545 15600 555 15640
rect 595 15600 4020 15640
rect 400 15585 4020 15600
rect 400 15210 4020 15225
rect 400 15170 405 15210
rect 445 15170 455 15210
rect 495 15170 505 15210
rect 545 15170 555 15210
rect 595 15170 4020 15210
rect 400 15160 4020 15170
rect 400 15120 405 15160
rect 445 15120 455 15160
rect 495 15120 505 15160
rect 545 15120 555 15160
rect 595 15120 4020 15160
rect 400 15105 4020 15120
rect 13255 14980 13335 15000
rect 13255 14940 13275 14980
rect 13315 14940 13335 14980
rect 13255 14920 13335 14940
rect 100 14820 4020 14835
rect 100 14780 105 14820
rect 145 14780 155 14820
rect 195 14780 205 14820
rect 245 14780 255 14820
rect 295 14780 4020 14820
rect 100 14770 4020 14780
rect 100 14730 105 14770
rect 145 14730 155 14770
rect 195 14730 205 14770
rect 245 14730 255 14770
rect 295 14730 4020 14770
rect 100 14715 4020 14730
rect 100 14160 4020 14175
rect 100 14120 105 14160
rect 145 14120 155 14160
rect 195 14120 205 14160
rect 245 14120 255 14160
rect 295 14120 4020 14160
rect 100 14110 4020 14120
rect 100 14070 105 14110
rect 145 14070 155 14110
rect 195 14070 205 14110
rect 245 14070 255 14110
rect 295 14070 4020 14110
rect 100 14055 4020 14070
rect 400 14010 4020 14025
rect 400 13970 405 14010
rect 445 13970 455 14010
rect 495 13970 505 14010
rect 545 13970 555 14010
rect 595 13970 4020 14010
rect 400 13960 4020 13970
rect 400 13920 405 13960
rect 445 13920 455 13960
rect 495 13920 505 13960
rect 545 13920 555 13960
rect 595 13920 4020 13960
rect 400 13905 4020 13920
rect 100 13420 4020 13435
rect 100 13380 105 13420
rect 145 13380 155 13420
rect 195 13380 205 13420
rect 245 13380 255 13420
rect 295 13380 4020 13420
rect 100 13370 4020 13380
rect 100 13330 105 13370
rect 145 13330 155 13370
rect 195 13330 205 13370
rect 245 13330 255 13370
rect 295 13330 4020 13370
rect 100 13315 4020 13330
rect 400 12830 4020 12845
rect 400 12790 405 12830
rect 445 12790 455 12830
rect 495 12790 505 12830
rect 545 12790 555 12830
rect 595 12790 4020 12830
rect 400 12780 4020 12790
rect 400 12740 405 12780
rect 445 12740 455 12780
rect 495 12740 505 12780
rect 545 12740 555 12780
rect 595 12740 4020 12780
rect 400 12725 4020 12740
rect 400 12655 4020 12670
rect 400 12615 405 12655
rect 445 12615 455 12655
rect 495 12615 505 12655
rect 545 12615 555 12655
rect 595 12615 4020 12655
rect 400 12605 4020 12615
rect 400 12565 405 12605
rect 445 12565 455 12605
rect 495 12565 505 12605
rect 545 12565 555 12605
rect 595 12565 4020 12605
rect 400 12550 4020 12565
rect 100 12505 4020 12520
rect 100 12465 105 12505
rect 145 12465 155 12505
rect 195 12465 205 12505
rect 245 12465 255 12505
rect 295 12465 4020 12505
rect 100 12455 4020 12465
rect 100 12415 105 12455
rect 145 12415 155 12455
rect 195 12415 205 12455
rect 245 12415 255 12455
rect 295 12415 4020 12455
rect 100 12400 4020 12415
rect 400 7480 4020 7495
rect 400 7440 405 7480
rect 445 7440 455 7480
rect 495 7440 505 7480
rect 545 7440 555 7480
rect 595 7475 4020 7480
rect 595 7445 3895 7475
rect 3925 7445 3940 7475
rect 3970 7445 3985 7475
rect 4015 7445 4020 7475
rect 595 7440 4020 7445
rect 400 7430 4020 7440
rect 400 7390 405 7430
rect 445 7390 455 7430
rect 495 7390 505 7430
rect 545 7390 555 7430
rect 595 7425 4020 7430
rect 595 7395 3895 7425
rect 3925 7395 3940 7425
rect 3970 7395 3985 7425
rect 4015 7395 4020 7425
rect 595 7390 4020 7395
rect 400 7375 4020 7390
rect 400 7150 4020 7155
rect 400 7140 3895 7150
rect 400 7100 405 7140
rect 445 7100 455 7140
rect 495 7100 505 7140
rect 545 7100 555 7140
rect 595 7120 3895 7140
rect 3925 7120 3940 7150
rect 3970 7120 3985 7150
rect 4015 7120 4020 7150
rect 595 7105 4020 7120
rect 595 7100 3895 7105
rect 400 7080 3895 7100
rect 400 7040 405 7080
rect 445 7040 455 7080
rect 495 7040 505 7080
rect 545 7040 555 7080
rect 595 7075 3895 7080
rect 3925 7075 3940 7105
rect 3970 7075 3985 7105
rect 4015 7075 4020 7105
rect 595 7060 4020 7075
rect 595 7040 3895 7060
rect 400 7030 3895 7040
rect 3925 7030 3940 7060
rect 3970 7030 3985 7060
rect 4015 7030 4020 7060
rect 400 7025 4020 7030
<< via3 >>
rect 405 15650 445 15690
rect 455 15650 495 15690
rect 505 15650 545 15690
rect 555 15650 595 15690
rect 15205 15700 15245 15740
rect 405 15600 445 15640
rect 455 15600 495 15640
rect 505 15600 545 15640
rect 555 15600 595 15640
rect 405 15170 445 15210
rect 455 15170 495 15210
rect 505 15170 545 15210
rect 555 15170 595 15210
rect 405 15120 445 15160
rect 455 15120 495 15160
rect 505 15120 545 15160
rect 555 15120 595 15160
rect 13275 14940 13315 14980
rect 105 14780 145 14820
rect 155 14780 195 14820
rect 205 14780 245 14820
rect 255 14780 295 14820
rect 105 14730 145 14770
rect 155 14730 195 14770
rect 205 14730 245 14770
rect 255 14730 295 14770
rect 105 14120 145 14160
rect 155 14120 195 14160
rect 205 14120 245 14160
rect 255 14120 295 14160
rect 105 14070 145 14110
rect 155 14070 195 14110
rect 205 14070 245 14110
rect 255 14070 295 14110
rect 405 13970 445 14010
rect 455 13970 495 14010
rect 505 13970 545 14010
rect 555 13970 595 14010
rect 405 13920 445 13960
rect 455 13920 495 13960
rect 505 13920 545 13960
rect 555 13920 595 13960
rect 105 13380 145 13420
rect 155 13380 195 13420
rect 205 13380 245 13420
rect 255 13380 295 13420
rect 105 13330 145 13370
rect 155 13330 195 13370
rect 205 13330 245 13370
rect 255 13330 295 13370
rect 405 12790 445 12830
rect 455 12790 495 12830
rect 505 12790 545 12830
rect 555 12790 595 12830
rect 405 12740 445 12780
rect 455 12740 495 12780
rect 505 12740 545 12780
rect 555 12740 595 12780
rect 405 12615 445 12655
rect 455 12615 495 12655
rect 505 12615 545 12655
rect 555 12615 595 12655
rect 405 12565 445 12605
rect 455 12565 495 12605
rect 505 12565 545 12605
rect 555 12565 595 12605
rect 105 12465 145 12505
rect 155 12465 195 12505
rect 205 12465 245 12505
rect 255 12465 295 12505
rect 105 12415 145 12455
rect 155 12415 195 12455
rect 205 12415 245 12455
rect 255 12415 295 12455
rect 405 7440 445 7480
rect 455 7440 495 7480
rect 505 7440 545 7480
rect 555 7440 595 7480
rect 405 7390 445 7430
rect 455 7390 495 7430
rect 505 7390 545 7430
rect 555 7390 595 7430
rect 405 7100 445 7140
rect 455 7100 495 7140
rect 505 7100 545 7140
rect 555 7100 595 7140
rect 405 7040 445 7080
rect 455 7040 495 7080
rect 505 7040 545 7080
rect 555 7040 595 7080
<< metal4 >>
rect 100 14820 300 22076
rect 100 14780 105 14820
rect 145 14780 155 14820
rect 195 14780 205 14820
rect 245 14780 255 14820
rect 295 14780 300 14820
rect 100 14770 300 14780
rect 100 14730 105 14770
rect 145 14730 155 14770
rect 195 14730 205 14770
rect 245 14730 255 14770
rect 295 14730 300 14770
rect 100 14160 300 14730
rect 100 14120 105 14160
rect 145 14120 155 14160
rect 195 14120 205 14160
rect 245 14120 255 14160
rect 295 14120 300 14160
rect 100 14110 300 14120
rect 100 14070 105 14110
rect 145 14070 155 14110
rect 195 14070 205 14110
rect 245 14070 255 14110
rect 295 14070 300 14110
rect 100 13420 300 14070
rect 100 13380 105 13420
rect 145 13380 155 13420
rect 195 13380 205 13420
rect 245 13380 255 13420
rect 295 13380 300 13420
rect 100 13370 300 13380
rect 100 13330 105 13370
rect 145 13330 155 13370
rect 195 13330 205 13370
rect 245 13330 255 13370
rect 295 13330 300 13370
rect 100 12505 300 13330
rect 100 12465 105 12505
rect 145 12465 155 12505
rect 195 12465 205 12505
rect 245 12465 255 12505
rect 295 12465 300 12505
rect 100 12455 300 12465
rect 100 12415 105 12455
rect 145 12415 155 12455
rect 195 12415 205 12455
rect 245 12415 255 12455
rect 295 12415 300 12455
rect 100 500 300 12415
rect 400 15690 600 22076
rect 400 15650 405 15690
rect 445 15650 455 15690
rect 495 15650 505 15690
rect 545 15650 555 15690
rect 595 15650 600 15690
rect 400 15640 600 15650
rect 400 15600 405 15640
rect 445 15600 455 15640
rect 495 15600 505 15640
rect 545 15600 555 15640
rect 595 15600 600 15640
rect 400 15210 600 15600
rect 400 15170 405 15210
rect 445 15170 455 15210
rect 495 15170 505 15210
rect 545 15170 555 15210
rect 595 15170 600 15210
rect 400 15160 600 15170
rect 400 15120 405 15160
rect 445 15120 455 15160
rect 495 15120 505 15160
rect 545 15120 555 15160
rect 595 15120 600 15160
rect 400 14010 600 15120
rect 15185 15740 15265 15760
rect 15185 15700 15205 15740
rect 15245 15700 15265 15740
rect 400 13970 405 14010
rect 445 13970 455 14010
rect 495 13970 505 14010
rect 545 13970 555 14010
rect 595 13970 600 14010
rect 400 13960 600 13970
rect 400 13920 405 13960
rect 445 13920 455 13960
rect 495 13920 505 13960
rect 545 13920 555 13960
rect 595 13920 600 13960
rect 400 12830 600 13920
rect 400 12790 405 12830
rect 445 12790 455 12830
rect 495 12790 505 12830
rect 545 12790 555 12830
rect 595 12790 600 12830
rect 400 12780 600 12790
rect 400 12740 405 12780
rect 445 12740 455 12780
rect 495 12740 505 12780
rect 545 12740 555 12780
rect 595 12740 600 12780
rect 400 12655 600 12740
rect 400 12615 405 12655
rect 445 12615 455 12655
rect 495 12615 505 12655
rect 545 12615 555 12655
rect 595 12615 600 12655
rect 400 12605 600 12615
rect 400 12565 405 12605
rect 445 12565 455 12605
rect 495 12565 505 12605
rect 545 12565 555 12605
rect 595 12565 600 12605
rect 400 7480 600 12565
rect 400 7440 405 7480
rect 445 7440 455 7480
rect 495 7440 505 7480
rect 545 7440 555 7480
rect 595 7440 600 7480
rect 400 7430 600 7440
rect 400 7390 405 7430
rect 445 7390 455 7430
rect 495 7390 505 7430
rect 545 7390 555 7430
rect 595 7390 600 7430
rect 400 7140 600 7390
rect 400 7100 405 7140
rect 445 7100 455 7140
rect 495 7100 505 7140
rect 545 7100 555 7140
rect 595 7100 600 7140
rect 400 7080 600 7100
rect 400 7040 405 7080
rect 445 7040 455 7080
rect 495 7040 505 7080
rect 545 7040 555 7080
rect 595 7040 600 7080
rect 400 500 600 7040
rect 13255 14980 13335 15000
rect 13255 14940 13275 14980
rect 13315 14940 13335 14980
rect 13255 100 13335 14940
rect 15185 100 15265 15700
rect 13249 0 13339 100
rect 15181 0 15271 100
use pll_bgr_magic_3_flat  pll_bgr_magic_3_flat_0
timestamp 1756757103
transform 1 0 6155 0 1 8755
box -2135 -7840 7050 6950
<< labels >>
flabel metal4 s 15181 0 15271 100 0 FreeSans 480 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 13249 0 13339 100 0 FreeSans 480 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 100 500 300 22076 1 FreeSans 200 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 400 500 600 22076 1 FreeSans 200 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal1 12150 13445 12150 13445 3 FreeSans 800 0 400 0 V_CONT
<< properties >>
string FIXED_BBOX 0 0 16100 22576
<< end >>
