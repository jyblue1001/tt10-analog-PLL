magic
tech sky130A
magscale 1 2
timestamp 1756577835
<< nwell >>
rect 390 7590 3120 7870
rect 3420 7590 6150 7870
rect 9960 7400 10710 7420
rect 1490 6030 5050 6710
rect 5350 6230 6120 6510
rect 8110 6090 11550 7400
rect 1500 5430 3140 5710
rect 3400 5430 5040 5710
rect 2020 3110 7000 4350
rect 8000 3820 11220 4400
rect 12360 1240 14640 1260
rect 12150 1160 14640 1240
rect 1720 950 14640 1160
rect 12360 90 14640 950
<< pwell >>
rect 3230 14820 3310 15100
rect 1240 14667 2580 14820
rect 1240 13633 1393 14667
rect 2427 13633 2580 14667
rect 1240 13480 2580 13633
rect 2600 14667 3940 14820
rect 2600 13633 2753 14667
rect 3787 13633 3940 14667
rect 2600 13480 3940 13633
rect 3960 14667 5300 14820
rect 3960 13633 4113 14667
rect 5147 13633 5300 14667
rect 3960 13480 5300 13633
rect 1240 13307 2580 13460
rect 1240 12273 1393 13307
rect 2427 12273 2580 13307
rect 1240 12120 2580 12273
rect 2600 13307 3940 13460
rect 2600 12273 2753 13307
rect 3787 12273 3940 13307
rect 2600 12120 3940 12273
rect 3960 13307 5300 13460
rect 3960 12273 4113 13307
rect 5147 12273 5300 13307
rect 3960 12120 5300 12273
rect 1240 11947 2580 12100
rect 1240 10913 1393 11947
rect 2427 10913 2580 11947
rect 1240 10760 2580 10913
rect 2600 11947 3940 12100
rect 2600 10913 2753 11947
rect 3787 10913 3940 11947
rect 2600 10760 3940 10913
rect 3960 11947 5300 12100
rect 3960 10913 4113 11947
rect 5147 10913 5300 11947
rect 3960 10760 5300 10913
<< nbase >>
rect 1393 13633 2427 14667
rect 2753 13633 3787 14667
rect 4113 13633 5147 14667
rect 1393 12273 2427 13307
rect 2753 12273 3787 13307
rect 4113 12273 5147 13307
rect 1393 10913 2427 11947
rect 2753 10913 3787 11947
rect 4113 10913 5147 11947
<< nmos >>
rect 1230 10090 3230 10290
rect 3310 10090 5310 10290
rect 810 9180 1810 9680
rect 2050 9180 3050 9680
rect 3490 9180 4490 9680
rect 4730 9180 5730 9680
rect 1430 8570 1470 8670
rect 1550 8570 1590 8670
rect 1670 8570 1710 8670
rect 1790 8570 1830 8670
rect 1910 8570 1950 8670
rect 2030 8570 2070 8670
rect 2150 8570 2190 8670
rect 2270 8570 2310 8670
rect 2390 8570 2430 8670
rect 2510 8570 2550 8670
rect 3990 8570 4030 8670
rect 4110 8570 4150 8670
rect 4230 8570 4270 8670
rect 4350 8570 4390 8670
rect 4470 8570 4510 8670
rect 4590 8570 4630 8670
rect 4710 8570 4750 8670
rect 4830 8570 4870 8670
rect 4950 8570 4990 8670
rect 5070 8570 5110 8670
rect 8300 8360 8400 8610
rect 8500 8360 8600 8610
rect 8700 8360 8800 8610
rect 8900 8360 9000 8610
rect 9100 8360 9200 8610
rect 9300 8360 9400 8610
rect 9500 8360 9600 8610
rect 9700 8360 9800 8610
rect 9900 8360 10000 8610
rect 10100 8360 10200 8610
rect 8350 7820 8380 7920
rect 8480 7820 8510 7920
rect 8610 7820 8640 7920
rect 8740 7820 8770 7920
rect 8870 7820 8900 7920
rect 9000 7820 9030 7920
rect 9490 7820 9520 7920
rect 9620 7820 9650 7920
rect 9750 7820 9780 7920
rect 9880 7820 9910 7920
rect 10010 7820 10040 7920
rect 10140 7820 10170 7920
rect 10630 7820 10660 7920
rect 10760 7820 10790 7920
rect 10890 7820 10920 7920
rect 11020 7820 11050 7920
rect 11150 7820 11180 7920
rect 11280 7820 11310 7920
rect 2220 4530 2250 4730
rect 2330 4530 2360 4730
rect 2740 4530 2770 4730
rect 2850 4530 2880 4730
rect 3120 4530 3150 4730
rect 3230 4530 3260 4730
rect 3640 4530 3670 4730
rect 3750 4530 3780 4730
rect 4160 4530 4190 4730
rect 4270 4530 4300 4730
rect 4600 4530 4630 4730
rect 4930 4530 4960 4730
rect 5370 4530 5400 4730
rect 5760 4530 5790 4730
rect 6150 4530 6180 4730
rect 6440 4530 6470 4730
rect 8040 2980 8160 3380
rect 8260 2980 8380 3380
rect 8480 2980 8600 3380
rect 8700 2980 8820 3380
rect 9120 2980 9240 3380
rect 9340 2980 9460 3380
rect 9560 2980 9680 3380
rect 9780 2980 9900 3380
rect 10200 2980 10320 3380
rect 10420 2980 10540 3380
rect 10640 2980 10760 3380
rect 10860 2980 10980 3380
rect 2220 2730 2250 2930
rect 2330 2730 2360 2930
rect 2740 2730 2770 2930
rect 2850 2730 2880 2930
rect 3120 2730 3150 2930
rect 3230 2730 3260 2930
rect 3640 2730 3670 2930
rect 3750 2730 3780 2930
rect 4150 2730 4180 2930
rect 4480 2730 4510 2930
rect 4810 2730 4840 2930
rect 5370 2730 5400 2930
rect 5760 2730 5790 2930
rect 6150 2730 6180 2930
rect 6440 2730 6470 2930
rect 6830 2730 6860 2930
rect 12480 1800 12510 2000
rect 13080 1800 13110 2000
rect 13680 1800 13710 2000
rect 13950 1800 13980 2000
rect 12480 1570 12510 1670
rect 13080 1570 13110 1670
rect 13680 1570 13710 1670
rect 1910 1340 1940 1440
rect 2020 1340 2050 1440
rect 2130 1340 2160 1440
rect 2240 1340 2270 1440
rect 2490 1340 2520 1440
rect 2600 1340 2630 1440
rect 2940 1340 2970 1440
rect 3050 1340 3080 1440
rect 3160 1340 3190 1440
rect 3270 1340 3300 1440
rect 3600 1340 3630 1440
rect 3710 1340 3740 1440
rect 3820 1340 3850 1440
rect 3930 1340 3960 1440
rect 4280 1340 4310 1440
rect 4390 1340 4420 1440
rect 4500 1340 4530 1440
rect 4610 1340 4640 1440
rect 4860 1340 4890 1440
rect 4970 1340 5000 1440
rect 5420 1340 5450 1440
rect 5780 1340 5810 1440
rect 6030 1340 6060 1440
rect 6140 1340 6170 1440
rect 6250 1340 6280 1440
rect 6360 1340 6390 1440
rect 6690 1340 6720 1440
rect 6800 1340 6830 1440
rect 6910 1340 6940 1440
rect 7240 1340 7270 1440
rect 7350 1340 7380 1440
rect 7460 1340 7490 1440
rect 7570 1340 7600 1440
rect 7900 1340 7930 1440
rect 8010 1340 8040 1440
rect 8120 1340 8150 1440
rect 8540 1430 8570 1530
rect 8650 1430 8680 1530
rect 8760 1430 8790 1530
rect 8870 1430 8900 1530
rect 9200 1430 9230 1530
rect 9310 1430 9340 1530
rect 9420 1430 9450 1530
rect 9840 1430 9870 1530
rect 9950 1430 9980 1530
rect 10060 1430 10090 1530
rect 10170 1430 10200 1530
rect 10500 1430 10530 1530
rect 10610 1430 10640 1530
rect 10720 1430 10750 1530
rect 11140 1430 11170 1530
rect 11250 1430 11280 1530
rect 11360 1430 11390 1530
rect 11470 1430 11500 1530
rect 11800 1430 11830 1530
rect 11910 1430 11940 1530
rect 12020 1430 12050 1530
rect 12480 1330 12510 1430
rect 13080 1330 13110 1430
rect 13680 1330 13710 1430
<< pmos >>
rect 590 7630 630 7830
rect 710 7630 750 7830
rect 830 7630 870 7830
rect 950 7630 990 7830
rect 1070 7630 1110 7830
rect 1190 7630 1230 7830
rect 1310 7630 1350 7830
rect 1430 7630 1470 7830
rect 1550 7630 1590 7830
rect 1670 7630 1710 7830
rect 1790 7630 1830 7830
rect 1910 7630 1950 7830
rect 2030 7630 2070 7830
rect 2150 7630 2190 7830
rect 2270 7630 2310 7830
rect 2390 7630 2430 7830
rect 2510 7630 2550 7830
rect 2630 7630 2670 7830
rect 2750 7630 2790 7830
rect 2870 7630 2910 7830
rect 3630 7630 3670 7830
rect 3750 7630 3790 7830
rect 3870 7630 3910 7830
rect 3990 7630 4030 7830
rect 4110 7630 4150 7830
rect 4230 7630 4270 7830
rect 4350 7630 4390 7830
rect 4470 7630 4510 7830
rect 4590 7630 4630 7830
rect 4710 7630 4750 7830
rect 4830 7630 4870 7830
rect 4950 7630 4990 7830
rect 5070 7630 5110 7830
rect 5190 7630 5230 7830
rect 5310 7630 5350 7830
rect 5430 7630 5470 7830
rect 5550 7630 5590 7830
rect 5670 7630 5710 7830
rect 5790 7630 5830 7830
rect 5910 7630 5950 7830
rect 8350 7150 8380 7350
rect 8480 7150 8510 7350
rect 8610 7150 8640 7350
rect 8740 7150 8770 7350
rect 8870 7150 8900 7350
rect 9000 7150 9030 7350
rect 9490 7150 9520 7350
rect 9620 7150 9650 7350
rect 9750 7150 9780 7350
rect 9880 7150 9910 7350
rect 10010 7150 10040 7350
rect 10140 7150 10170 7350
rect 10630 7150 10660 7350
rect 10760 7150 10790 7350
rect 10890 7150 10920 7350
rect 11020 7150 11050 7350
rect 11150 7150 11180 7350
rect 11280 7150 11310 7350
rect 1690 6070 1790 6670
rect 1870 6070 1970 6670
rect 2050 6070 2150 6670
rect 2230 6070 2330 6670
rect 2410 6070 2510 6670
rect 2590 6070 2690 6670
rect 2770 6070 2870 6670
rect 2950 6070 3050 6670
rect 3130 6070 3230 6670
rect 3310 6070 3410 6670
rect 3490 6070 3590 6670
rect 3670 6070 3770 6670
rect 3850 6070 3950 6670
rect 4030 6070 4130 6670
rect 4210 6070 4310 6670
rect 4390 6070 4490 6670
rect 4570 6070 4670 6670
rect 4750 6070 4850 6670
rect 5560 6270 5590 6470
rect 5670 6270 5700 6470
rect 5780 6270 5810 6470
rect 5890 6270 5920 6470
rect 8420 6200 8520 6700
rect 8620 6200 8720 6700
rect 8820 6200 8920 6700
rect 9020 6200 9120 6700
rect 9220 6200 9320 6700
rect 9420 6200 9520 6700
rect 9620 6200 9720 6700
rect 9820 6200 9920 6700
rect 10020 6200 10120 6700
rect 10220 6200 10320 6700
rect 1700 5470 1730 5670
rect 1810 5470 1840 5670
rect 1920 5470 1950 5670
rect 2030 5470 2060 5670
rect 2140 5470 2170 5670
rect 2250 5470 2280 5670
rect 2360 5470 2390 5670
rect 2470 5470 2500 5670
rect 2580 5470 2610 5670
rect 2690 5470 2720 5670
rect 2800 5470 2830 5670
rect 2910 5470 2940 5670
rect 3600 5470 3630 5670
rect 3710 5470 3740 5670
rect 3820 5470 3850 5670
rect 3930 5470 3960 5670
rect 4040 5470 4070 5670
rect 4150 5470 4180 5670
rect 4260 5470 4290 5670
rect 4370 5470 4400 5670
rect 4480 5470 4510 5670
rect 4590 5470 4620 5670
rect 4700 5470 4730 5670
rect 4810 5470 4840 5670
rect 2220 3910 2250 4310
rect 2330 3910 2360 4310
rect 2740 3910 2770 4310
rect 2850 3910 2880 4310
rect 3120 3910 3150 4310
rect 3230 3910 3260 4310
rect 3640 3910 3670 4310
rect 3750 3910 3780 4310
rect 4160 3910 4190 4310
rect 4270 3910 4300 4310
rect 4600 3910 4630 4310
rect 4930 3910 4960 4310
rect 5370 3910 5400 4310
rect 5760 3910 5790 4310
rect 6150 3910 6180 4310
rect 6440 3910 6470 4310
rect 6830 3910 6860 4310
rect 8240 3960 8360 4360
rect 8460 3960 8580 4360
rect 8680 3960 8800 4360
rect 8900 3960 9020 4360
rect 9120 3960 9240 4360
rect 9340 3960 9460 4360
rect 9760 3960 9880 4360
rect 9980 3960 10100 4360
rect 10200 3960 10320 4360
rect 10420 3960 10540 4360
rect 10640 3960 10760 4360
rect 10860 3960 10980 4360
rect 2220 3150 2250 3550
rect 2330 3150 2360 3550
rect 2740 3150 2770 3550
rect 2850 3150 2880 3550
rect 3120 3150 3150 3550
rect 3230 3150 3260 3550
rect 3640 3150 3670 3550
rect 3750 3150 3780 3550
rect 4150 3150 4180 3550
rect 4480 3150 4510 3550
rect 4810 3150 4840 3550
rect 5370 3150 5400 3550
rect 5760 3150 5790 3550
rect 6150 3150 6180 3550
rect 6440 3150 6470 3550
rect 2070 1020 2100 1120
rect 2490 1020 2520 1120
rect 2600 1020 2630 1120
rect 3160 1020 3190 1120
rect 3270 1020 3300 1120
rect 3600 1020 3630 1120
rect 3710 1020 3740 1120
rect 3820 1020 3850 1120
rect 4440 1020 4470 1120
rect 4860 1020 4890 1120
rect 4970 1020 5000 1120
rect 5310 1020 5340 1120
rect 5420 1020 5450 1120
rect 5670 1020 5700 1120
rect 5780 1020 5810 1120
rect 6250 1020 6280 1120
rect 6360 1020 6390 1120
rect 6690 1020 6720 1120
rect 6800 1020 6830 1120
rect 7310 1020 7340 1120
rect 7650 1020 7680 1120
rect 7760 1020 7790 1120
rect 8010 1020 8040 1120
rect 8120 1020 8150 1120
rect 8610 1020 8640 1120
rect 8950 1020 8980 1120
rect 9060 1020 9090 1120
rect 9310 1020 9340 1120
rect 9420 1020 9450 1120
rect 9910 1020 9940 1120
rect 10250 1020 10280 1120
rect 10360 1020 10390 1120
rect 10610 1020 10640 1120
rect 10720 1020 10750 1120
rect 11210 1020 11240 1120
rect 11550 1020 11580 1120
rect 11660 1020 11690 1120
rect 11910 1020 11940 1120
rect 12020 1020 12050 1120
rect 12480 1020 12510 1220
rect 13080 1020 13110 1220
rect 13680 1020 13710 1220
rect 12480 680 12510 880
rect 13080 680 13110 880
rect 13680 680 13710 880
rect 12480 130 12780 530
rect 13080 130 13380 530
rect 13680 130 13980 530
rect 14220 130 14520 530
<< ndiff >>
rect 1150 10260 1230 10290
rect 1150 10220 1170 10260
rect 1210 10220 1230 10260
rect 1150 10160 1230 10220
rect 1150 10120 1170 10160
rect 1210 10120 1230 10160
rect 1150 10090 1230 10120
rect 3230 10260 3310 10290
rect 3230 10220 3250 10260
rect 3290 10220 3310 10260
rect 3230 10160 3310 10220
rect 3230 10120 3250 10160
rect 3290 10120 3310 10160
rect 3230 10090 3310 10120
rect 5310 10260 5390 10290
rect 5310 10220 5330 10260
rect 5370 10220 5390 10260
rect 5310 10160 5390 10220
rect 5310 10120 5330 10160
rect 5370 10120 5390 10160
rect 5310 10090 5390 10120
rect 730 9650 810 9680
rect 730 9610 750 9650
rect 790 9610 810 9650
rect 730 9550 810 9610
rect 730 9510 750 9550
rect 790 9510 810 9550
rect 730 9450 810 9510
rect 730 9410 750 9450
rect 790 9410 810 9450
rect 730 9350 810 9410
rect 730 9310 750 9350
rect 790 9310 810 9350
rect 730 9250 810 9310
rect 730 9210 750 9250
rect 790 9210 810 9250
rect 730 9180 810 9210
rect 1810 9650 1890 9680
rect 1970 9650 2050 9680
rect 1810 9610 1830 9650
rect 1870 9610 1890 9650
rect 1970 9610 1990 9650
rect 2030 9610 2050 9650
rect 1810 9550 1890 9610
rect 1970 9550 2050 9610
rect 1810 9510 1830 9550
rect 1870 9510 1890 9550
rect 1970 9510 1990 9550
rect 2030 9510 2050 9550
rect 1810 9450 1890 9510
rect 1970 9450 2050 9510
rect 1810 9410 1830 9450
rect 1870 9410 1890 9450
rect 1970 9410 1990 9450
rect 2030 9410 2050 9450
rect 1810 9350 1890 9410
rect 1970 9350 2050 9410
rect 1810 9310 1830 9350
rect 1870 9310 1890 9350
rect 1970 9310 1990 9350
rect 2030 9310 2050 9350
rect 1810 9250 1890 9310
rect 1970 9250 2050 9310
rect 1810 9210 1830 9250
rect 1870 9210 1890 9250
rect 1970 9210 1990 9250
rect 2030 9210 2050 9250
rect 1810 9180 1890 9210
rect 1970 9180 2050 9210
rect 3050 9650 3130 9680
rect 3050 9610 3070 9650
rect 3110 9610 3130 9650
rect 3050 9550 3130 9610
rect 3050 9510 3070 9550
rect 3110 9510 3130 9550
rect 3050 9450 3130 9510
rect 3050 9410 3070 9450
rect 3110 9410 3130 9450
rect 3050 9350 3130 9410
rect 3050 9310 3070 9350
rect 3110 9310 3130 9350
rect 3050 9250 3130 9310
rect 3050 9210 3070 9250
rect 3110 9210 3130 9250
rect 3050 9180 3130 9210
rect 3410 9650 3490 9680
rect 3410 9610 3430 9650
rect 3470 9610 3490 9650
rect 3410 9550 3490 9610
rect 3410 9510 3430 9550
rect 3470 9510 3490 9550
rect 3410 9450 3490 9510
rect 3410 9410 3430 9450
rect 3470 9410 3490 9450
rect 3410 9350 3490 9410
rect 3410 9310 3430 9350
rect 3470 9310 3490 9350
rect 3410 9250 3490 9310
rect 3410 9210 3430 9250
rect 3470 9210 3490 9250
rect 3410 9180 3490 9210
rect 4490 9670 4730 9680
rect 4490 9650 4570 9670
rect 4650 9650 4730 9670
rect 4490 9610 4510 9650
rect 4550 9610 4570 9650
rect 4650 9610 4670 9650
rect 4710 9610 4730 9650
rect 4490 9550 4570 9610
rect 4650 9550 4730 9610
rect 4490 9510 4510 9550
rect 4550 9510 4570 9550
rect 4650 9510 4670 9550
rect 4710 9510 4730 9550
rect 4490 9450 4570 9510
rect 4650 9450 4730 9510
rect 4490 9410 4510 9450
rect 4550 9410 4570 9450
rect 4650 9410 4670 9450
rect 4710 9410 4730 9450
rect 4490 9350 4570 9410
rect 4650 9350 4730 9410
rect 4490 9310 4510 9350
rect 4550 9310 4570 9350
rect 4650 9310 4670 9350
rect 4710 9310 4730 9350
rect 4490 9250 4570 9310
rect 4650 9250 4730 9310
rect 4490 9210 4510 9250
rect 4550 9210 4570 9250
rect 4650 9210 4670 9250
rect 4710 9210 4730 9250
rect 4490 9180 4570 9210
rect 4650 9180 4730 9210
rect 5730 9650 5810 9680
rect 5730 9610 5750 9650
rect 5790 9610 5810 9650
rect 5730 9550 5810 9610
rect 5730 9510 5750 9550
rect 5790 9510 5810 9550
rect 5730 9450 5810 9510
rect 5730 9410 5750 9450
rect 5790 9410 5810 9450
rect 5730 9350 5810 9410
rect 5730 9310 5750 9350
rect 5790 9310 5810 9350
rect 5730 9250 5810 9310
rect 5730 9210 5750 9250
rect 5790 9210 5810 9250
rect 5730 9180 5810 9210
rect 1350 8640 1430 8670
rect 1350 8600 1370 8640
rect 1410 8600 1430 8640
rect 1350 8570 1430 8600
rect 1470 8640 1550 8670
rect 1470 8600 1490 8640
rect 1530 8600 1550 8640
rect 1470 8570 1550 8600
rect 1590 8640 1670 8670
rect 1590 8600 1610 8640
rect 1650 8600 1670 8640
rect 1590 8570 1670 8600
rect 1710 8640 1790 8670
rect 1710 8600 1730 8640
rect 1770 8600 1790 8640
rect 1710 8570 1790 8600
rect 1830 8640 1910 8670
rect 1830 8600 1850 8640
rect 1890 8600 1910 8640
rect 1830 8570 1910 8600
rect 1950 8640 2030 8670
rect 1950 8600 1970 8640
rect 2010 8600 2030 8640
rect 1950 8570 2030 8600
rect 2070 8640 2150 8670
rect 2070 8600 2090 8640
rect 2130 8600 2150 8640
rect 2070 8570 2150 8600
rect 2190 8640 2270 8670
rect 2190 8600 2210 8640
rect 2250 8600 2270 8640
rect 2190 8570 2270 8600
rect 2310 8640 2390 8670
rect 2310 8600 2330 8640
rect 2370 8600 2390 8640
rect 2310 8570 2390 8600
rect 2430 8640 2510 8670
rect 2430 8600 2450 8640
rect 2490 8600 2510 8640
rect 2430 8570 2510 8600
rect 2550 8640 2630 8670
rect 2550 8600 2570 8640
rect 2610 8600 2630 8640
rect 2550 8570 2630 8600
rect 3910 8640 3990 8670
rect 3910 8600 3930 8640
rect 3970 8600 3990 8640
rect 3910 8570 3990 8600
rect 4030 8640 4110 8670
rect 4030 8600 4050 8640
rect 4090 8600 4110 8640
rect 4030 8570 4110 8600
rect 4150 8640 4230 8670
rect 4150 8600 4170 8640
rect 4210 8600 4230 8640
rect 4150 8570 4230 8600
rect 4270 8640 4350 8670
rect 4270 8600 4290 8640
rect 4330 8600 4350 8640
rect 4270 8570 4350 8600
rect 4390 8640 4470 8670
rect 4390 8600 4410 8640
rect 4450 8600 4470 8640
rect 4390 8570 4470 8600
rect 4510 8640 4590 8670
rect 4510 8600 4530 8640
rect 4570 8600 4590 8640
rect 4510 8570 4590 8600
rect 4630 8640 4710 8670
rect 4630 8600 4650 8640
rect 4690 8600 4710 8640
rect 4630 8570 4710 8600
rect 4750 8640 4830 8670
rect 4750 8600 4770 8640
rect 4810 8600 4830 8640
rect 4750 8570 4830 8600
rect 4870 8640 4950 8670
rect 4870 8600 4890 8640
rect 4930 8600 4950 8640
rect 4870 8570 4950 8600
rect 4990 8640 5070 8670
rect 4990 8600 5010 8640
rect 5050 8600 5070 8640
rect 4990 8570 5070 8600
rect 5110 8640 5190 8670
rect 5110 8600 5130 8640
rect 5170 8600 5190 8640
rect 5110 8570 5190 8600
rect 8200 8580 8300 8610
rect 8200 8530 8230 8580
rect 8270 8530 8300 8580
rect 8200 8440 8300 8530
rect 8200 8390 8230 8440
rect 8270 8390 8300 8440
rect 8200 8360 8300 8390
rect 8400 8580 8500 8610
rect 8400 8530 8430 8580
rect 8470 8530 8500 8580
rect 8400 8440 8500 8530
rect 8400 8390 8430 8440
rect 8470 8390 8500 8440
rect 8400 8360 8500 8390
rect 8600 8580 8700 8610
rect 8600 8530 8630 8580
rect 8670 8530 8700 8580
rect 8600 8440 8700 8530
rect 8600 8390 8630 8440
rect 8670 8390 8700 8440
rect 8600 8360 8700 8390
rect 8800 8580 8900 8610
rect 8800 8530 8830 8580
rect 8870 8530 8900 8580
rect 8800 8440 8900 8530
rect 8800 8390 8830 8440
rect 8870 8390 8900 8440
rect 8800 8360 8900 8390
rect 9000 8580 9100 8610
rect 9000 8530 9030 8580
rect 9070 8530 9100 8580
rect 9000 8440 9100 8530
rect 9000 8390 9030 8440
rect 9070 8390 9100 8440
rect 9000 8360 9100 8390
rect 9200 8580 9300 8610
rect 9200 8530 9230 8580
rect 9270 8530 9300 8580
rect 9200 8440 9300 8530
rect 9200 8390 9230 8440
rect 9270 8390 9300 8440
rect 9200 8360 9300 8390
rect 9400 8580 9500 8610
rect 9400 8530 9430 8580
rect 9470 8530 9500 8580
rect 9400 8440 9500 8530
rect 9400 8390 9430 8440
rect 9470 8390 9500 8440
rect 9400 8360 9500 8390
rect 9600 8580 9700 8610
rect 9600 8530 9630 8580
rect 9670 8530 9700 8580
rect 9600 8440 9700 8530
rect 9600 8390 9630 8440
rect 9670 8390 9700 8440
rect 9600 8360 9700 8390
rect 9800 8580 9900 8610
rect 9800 8530 9830 8580
rect 9870 8530 9900 8580
rect 9800 8440 9900 8530
rect 9800 8390 9830 8440
rect 9870 8390 9900 8440
rect 9800 8360 9900 8390
rect 10000 8580 10100 8610
rect 10000 8530 10030 8580
rect 10070 8530 10100 8580
rect 10000 8440 10100 8530
rect 10000 8390 10030 8440
rect 10070 8390 10100 8440
rect 10000 8360 10100 8390
rect 10200 8580 10300 8610
rect 10200 8530 10230 8580
rect 10270 8530 10300 8580
rect 10200 8440 10300 8530
rect 10200 8390 10230 8440
rect 10270 8390 10300 8440
rect 10200 8360 10300 8390
rect 8250 7890 8350 7920
rect 8250 7850 8280 7890
rect 8320 7850 8350 7890
rect 8250 7820 8350 7850
rect 8380 7890 8480 7920
rect 8380 7850 8410 7890
rect 8450 7850 8480 7890
rect 8380 7820 8480 7850
rect 8510 7890 8610 7920
rect 8510 7850 8540 7890
rect 8580 7850 8610 7890
rect 8510 7820 8610 7850
rect 8640 7890 8740 7920
rect 8640 7850 8670 7890
rect 8710 7850 8740 7890
rect 8640 7820 8740 7850
rect 8770 7890 8870 7920
rect 8770 7850 8800 7890
rect 8840 7850 8870 7890
rect 8770 7820 8870 7850
rect 8900 7890 9000 7920
rect 8900 7850 8930 7890
rect 8970 7850 9000 7890
rect 8900 7820 9000 7850
rect 9030 7890 9130 7920
rect 9030 7850 9060 7890
rect 9100 7850 9130 7890
rect 9030 7820 9130 7850
rect 9390 7890 9490 7920
rect 9390 7850 9420 7890
rect 9460 7850 9490 7890
rect 9390 7820 9490 7850
rect 9520 7890 9620 7920
rect 9520 7850 9550 7890
rect 9590 7850 9620 7890
rect 9520 7820 9620 7850
rect 9650 7890 9750 7920
rect 9650 7850 9680 7890
rect 9720 7850 9750 7890
rect 9650 7820 9750 7850
rect 9780 7890 9880 7920
rect 9780 7850 9810 7890
rect 9850 7850 9880 7890
rect 9780 7820 9880 7850
rect 9910 7890 10010 7920
rect 9910 7850 9940 7890
rect 9980 7850 10010 7890
rect 9910 7820 10010 7850
rect 10040 7890 10140 7920
rect 10040 7850 10070 7890
rect 10110 7850 10140 7890
rect 10040 7820 10140 7850
rect 10170 7890 10270 7920
rect 10170 7850 10200 7890
rect 10240 7850 10270 7890
rect 10170 7820 10270 7850
rect 10530 7890 10630 7920
rect 10530 7850 10560 7890
rect 10600 7850 10630 7890
rect 10530 7820 10630 7850
rect 10660 7890 10760 7920
rect 10660 7850 10690 7890
rect 10730 7850 10760 7890
rect 10660 7820 10760 7850
rect 10790 7890 10890 7920
rect 10790 7850 10820 7890
rect 10860 7850 10890 7890
rect 10790 7820 10890 7850
rect 10920 7890 11020 7920
rect 10920 7850 10950 7890
rect 10990 7850 11020 7890
rect 10920 7820 11020 7850
rect 11050 7890 11150 7920
rect 11050 7850 11080 7890
rect 11120 7850 11150 7890
rect 11050 7820 11150 7850
rect 11180 7890 11280 7920
rect 11180 7850 11210 7890
rect 11250 7850 11280 7890
rect 11180 7820 11280 7850
rect 11310 7890 11410 7920
rect 11310 7850 11340 7890
rect 11380 7850 11410 7890
rect 11310 7820 11410 7850
rect 2140 4700 2220 4730
rect 2140 4660 2160 4700
rect 2200 4660 2220 4700
rect 2140 4600 2220 4660
rect 2140 4560 2160 4600
rect 2200 4560 2220 4600
rect 2140 4530 2220 4560
rect 2250 4700 2330 4730
rect 2250 4660 2270 4700
rect 2310 4660 2330 4700
rect 2250 4600 2330 4660
rect 2250 4560 2270 4600
rect 2310 4560 2330 4600
rect 2250 4530 2330 4560
rect 2360 4700 2440 4730
rect 2360 4660 2380 4700
rect 2420 4660 2440 4700
rect 2360 4600 2440 4660
rect 2360 4560 2380 4600
rect 2420 4560 2440 4600
rect 2360 4530 2440 4560
rect 2660 4700 2740 4730
rect 2660 4660 2680 4700
rect 2720 4660 2740 4700
rect 2660 4600 2740 4660
rect 2660 4560 2680 4600
rect 2720 4560 2740 4600
rect 2660 4530 2740 4560
rect 2770 4700 2850 4730
rect 2770 4660 2790 4700
rect 2830 4660 2850 4700
rect 2770 4600 2850 4660
rect 2770 4560 2790 4600
rect 2830 4560 2850 4600
rect 2770 4530 2850 4560
rect 2880 4700 2960 4730
rect 3040 4700 3120 4730
rect 2880 4660 2900 4700
rect 2940 4660 2960 4700
rect 3040 4660 3060 4700
rect 3100 4660 3120 4700
rect 2880 4600 2960 4660
rect 3040 4600 3120 4660
rect 2880 4560 2900 4600
rect 2940 4560 2960 4600
rect 3040 4560 3060 4600
rect 3100 4560 3120 4600
rect 2880 4530 2960 4560
rect 3040 4530 3120 4560
rect 3150 4700 3230 4730
rect 3150 4660 3170 4700
rect 3210 4660 3230 4700
rect 3150 4600 3230 4660
rect 3150 4560 3170 4600
rect 3210 4560 3230 4600
rect 3150 4530 3230 4560
rect 3260 4700 3340 4730
rect 3260 4660 3280 4700
rect 3320 4660 3340 4700
rect 3260 4600 3340 4660
rect 3260 4560 3280 4600
rect 3320 4560 3340 4600
rect 3260 4530 3340 4560
rect 3560 4700 3640 4730
rect 3560 4660 3580 4700
rect 3620 4660 3640 4700
rect 3560 4600 3640 4660
rect 3560 4560 3580 4600
rect 3620 4560 3640 4600
rect 3560 4530 3640 4560
rect 3670 4700 3750 4730
rect 3670 4660 3690 4700
rect 3730 4660 3750 4700
rect 3670 4600 3750 4660
rect 3670 4560 3690 4600
rect 3730 4560 3750 4600
rect 3670 4530 3750 4560
rect 3780 4700 3860 4730
rect 3780 4660 3800 4700
rect 3840 4660 3860 4700
rect 3780 4600 3860 4660
rect 3780 4560 3800 4600
rect 3840 4560 3860 4600
rect 3780 4530 3860 4560
rect 4080 4700 4160 4730
rect 4080 4660 4100 4700
rect 4140 4660 4160 4700
rect 4080 4600 4160 4660
rect 4080 4560 4100 4600
rect 4140 4560 4160 4600
rect 4080 4530 4160 4560
rect 4190 4700 4270 4730
rect 4190 4660 4210 4700
rect 4250 4660 4270 4700
rect 4190 4600 4270 4660
rect 4190 4560 4210 4600
rect 4250 4560 4270 4600
rect 4190 4530 4270 4560
rect 4300 4700 4380 4730
rect 4300 4660 4320 4700
rect 4360 4660 4380 4700
rect 4300 4600 4380 4660
rect 4300 4560 4320 4600
rect 4360 4560 4380 4600
rect 4300 4530 4380 4560
rect 4520 4700 4600 4730
rect 4520 4660 4540 4700
rect 4580 4660 4600 4700
rect 4520 4600 4600 4660
rect 4520 4560 4540 4600
rect 4580 4560 4600 4600
rect 4520 4530 4600 4560
rect 4630 4700 4710 4730
rect 4630 4660 4650 4700
rect 4690 4660 4710 4700
rect 4630 4600 4710 4660
rect 4630 4560 4650 4600
rect 4690 4560 4710 4600
rect 4630 4530 4710 4560
rect 4850 4700 4930 4730
rect 4850 4660 4870 4700
rect 4910 4660 4930 4700
rect 4850 4600 4930 4660
rect 4850 4560 4870 4600
rect 4910 4560 4930 4600
rect 4850 4530 4930 4560
rect 4960 4700 5040 4730
rect 4960 4660 4980 4700
rect 5020 4660 5040 4700
rect 4960 4600 5040 4660
rect 4960 4560 4980 4600
rect 5020 4560 5040 4600
rect 4960 4530 5040 4560
rect 5270 4700 5370 4730
rect 5270 4660 5300 4700
rect 5340 4660 5370 4700
rect 5270 4600 5370 4660
rect 5270 4560 5300 4600
rect 5340 4560 5370 4600
rect 5270 4530 5370 4560
rect 5400 4700 5500 4730
rect 5400 4660 5430 4700
rect 5470 4660 5500 4700
rect 5400 4600 5500 4660
rect 5400 4560 5430 4600
rect 5470 4560 5500 4600
rect 5400 4530 5500 4560
rect 5660 4700 5760 4730
rect 5660 4660 5690 4700
rect 5730 4660 5760 4700
rect 5660 4600 5760 4660
rect 5660 4560 5690 4600
rect 5730 4560 5760 4600
rect 5660 4530 5760 4560
rect 5790 4700 5890 4730
rect 5790 4660 5820 4700
rect 5860 4660 5890 4700
rect 5790 4600 5890 4660
rect 5790 4560 5820 4600
rect 5860 4560 5890 4600
rect 5790 4530 5890 4560
rect 6050 4700 6150 4730
rect 6050 4660 6080 4700
rect 6120 4660 6150 4700
rect 6050 4600 6150 4660
rect 6050 4560 6080 4600
rect 6120 4560 6150 4600
rect 6050 4530 6150 4560
rect 6180 4700 6280 4730
rect 6180 4660 6210 4700
rect 6250 4660 6280 4700
rect 6180 4600 6280 4660
rect 6180 4560 6210 4600
rect 6250 4560 6280 4600
rect 6180 4530 6280 4560
rect 6340 4700 6440 4730
rect 6340 4660 6370 4700
rect 6410 4660 6440 4700
rect 6340 4600 6440 4660
rect 6340 4560 6370 4600
rect 6410 4560 6440 4600
rect 6340 4530 6440 4560
rect 6470 4700 6570 4730
rect 6470 4660 6500 4700
rect 6540 4660 6570 4700
rect 6470 4600 6570 4660
rect 6470 4560 6500 4600
rect 6540 4560 6570 4600
rect 6470 4530 6570 4560
rect 7940 3350 8040 3380
rect 7940 3310 7970 3350
rect 8010 3310 8040 3350
rect 7940 3250 8040 3310
rect 7940 3210 7970 3250
rect 8010 3210 8040 3250
rect 7940 3150 8040 3210
rect 7940 3110 7970 3150
rect 8010 3110 8040 3150
rect 7940 3050 8040 3110
rect 7940 3010 7970 3050
rect 8010 3010 8040 3050
rect 7940 2980 8040 3010
rect 8160 3350 8260 3380
rect 8160 3310 8190 3350
rect 8230 3310 8260 3350
rect 8160 3250 8260 3310
rect 8160 3210 8190 3250
rect 8230 3210 8260 3250
rect 8160 3150 8260 3210
rect 8160 3110 8190 3150
rect 8230 3110 8260 3150
rect 8160 3050 8260 3110
rect 8160 3010 8190 3050
rect 8230 3010 8260 3050
rect 8160 2980 8260 3010
rect 8380 3350 8480 3380
rect 8380 3310 8410 3350
rect 8450 3310 8480 3350
rect 8380 3250 8480 3310
rect 8380 3210 8410 3250
rect 8450 3210 8480 3250
rect 8380 3150 8480 3210
rect 8380 3110 8410 3150
rect 8450 3110 8480 3150
rect 8380 3050 8480 3110
rect 8380 3010 8410 3050
rect 8450 3010 8480 3050
rect 8380 2980 8480 3010
rect 8600 3350 8700 3380
rect 8600 3310 8630 3350
rect 8670 3310 8700 3350
rect 8600 3250 8700 3310
rect 8600 3210 8630 3250
rect 8670 3210 8700 3250
rect 8600 3150 8700 3210
rect 8600 3110 8630 3150
rect 8670 3110 8700 3150
rect 8600 3050 8700 3110
rect 8600 3010 8630 3050
rect 8670 3010 8700 3050
rect 8600 2980 8700 3010
rect 8820 3350 8920 3380
rect 9020 3350 9120 3380
rect 8820 3310 8850 3350
rect 8890 3310 8920 3350
rect 9020 3310 9050 3350
rect 9090 3310 9120 3350
rect 8820 3250 8920 3310
rect 9020 3250 9120 3310
rect 8820 3210 8850 3250
rect 8890 3210 8920 3250
rect 9020 3210 9050 3250
rect 9090 3210 9120 3250
rect 8820 3150 8920 3210
rect 9020 3150 9120 3210
rect 8820 3110 8850 3150
rect 8890 3110 8920 3150
rect 9020 3110 9050 3150
rect 9090 3110 9120 3150
rect 8820 3050 8920 3110
rect 9020 3050 9120 3110
rect 8820 3010 8850 3050
rect 8890 3010 8920 3050
rect 9020 3010 9050 3050
rect 9090 3010 9120 3050
rect 8820 2980 8920 3010
rect 9020 2980 9120 3010
rect 9240 3350 9340 3380
rect 9240 3310 9270 3350
rect 9310 3310 9340 3350
rect 9240 3250 9340 3310
rect 9240 3210 9270 3250
rect 9310 3210 9340 3250
rect 9240 3150 9340 3210
rect 9240 3110 9270 3150
rect 9310 3110 9340 3150
rect 9240 3050 9340 3110
rect 9240 3010 9270 3050
rect 9310 3010 9340 3050
rect 9240 2980 9340 3010
rect 9460 3350 9560 3380
rect 9460 3310 9490 3350
rect 9530 3310 9560 3350
rect 9460 3250 9560 3310
rect 9460 3210 9490 3250
rect 9530 3210 9560 3250
rect 9460 3150 9560 3210
rect 9460 3110 9490 3150
rect 9530 3110 9560 3150
rect 9460 3050 9560 3110
rect 9460 3010 9490 3050
rect 9530 3010 9560 3050
rect 9460 2980 9560 3010
rect 9680 3350 9780 3380
rect 9680 3310 9710 3350
rect 9750 3310 9780 3350
rect 9680 3250 9780 3310
rect 9680 3210 9710 3250
rect 9750 3210 9780 3250
rect 9680 3150 9780 3210
rect 9680 3110 9710 3150
rect 9750 3110 9780 3150
rect 9680 3050 9780 3110
rect 9680 3010 9710 3050
rect 9750 3010 9780 3050
rect 9680 2980 9780 3010
rect 9900 3350 10000 3380
rect 10100 3350 10200 3380
rect 9900 3310 9930 3350
rect 9970 3310 10000 3350
rect 10100 3310 10130 3350
rect 10170 3310 10200 3350
rect 9900 3250 10000 3310
rect 10100 3250 10200 3310
rect 9900 3210 9930 3250
rect 9970 3210 10000 3250
rect 10100 3210 10130 3250
rect 10170 3210 10200 3250
rect 9900 3150 10000 3210
rect 10100 3150 10200 3210
rect 9900 3110 9930 3150
rect 9970 3110 10000 3150
rect 10100 3110 10130 3150
rect 10170 3110 10200 3150
rect 9900 3050 10000 3110
rect 10100 3050 10200 3110
rect 9900 3010 9930 3050
rect 9970 3010 10000 3050
rect 10100 3010 10130 3050
rect 10170 3010 10200 3050
rect 9900 2980 10000 3010
rect 10100 2980 10200 3010
rect 10320 3350 10420 3380
rect 10320 3310 10350 3350
rect 10390 3310 10420 3350
rect 10320 3250 10420 3310
rect 10320 3210 10350 3250
rect 10390 3210 10420 3250
rect 10320 3150 10420 3210
rect 10320 3110 10350 3150
rect 10390 3110 10420 3150
rect 10320 3050 10420 3110
rect 10320 3010 10350 3050
rect 10390 3010 10420 3050
rect 10320 2980 10420 3010
rect 10540 3350 10640 3380
rect 10540 3310 10570 3350
rect 10610 3310 10640 3350
rect 10540 3250 10640 3310
rect 10540 3210 10570 3250
rect 10610 3210 10640 3250
rect 10540 3150 10640 3210
rect 10540 3110 10570 3150
rect 10610 3110 10640 3150
rect 10540 3050 10640 3110
rect 10540 3010 10570 3050
rect 10610 3010 10640 3050
rect 10540 2980 10640 3010
rect 10760 3350 10860 3380
rect 10760 3310 10790 3350
rect 10830 3310 10860 3350
rect 10760 3250 10860 3310
rect 10760 3210 10790 3250
rect 10830 3210 10860 3250
rect 10760 3150 10860 3210
rect 10760 3110 10790 3150
rect 10830 3110 10860 3150
rect 10760 3050 10860 3110
rect 10760 3010 10790 3050
rect 10830 3010 10860 3050
rect 10760 2980 10860 3010
rect 10980 3350 11080 3380
rect 10980 3310 11010 3350
rect 11050 3310 11080 3350
rect 10980 3250 11080 3310
rect 10980 3210 11010 3250
rect 11050 3210 11080 3250
rect 10980 3150 11080 3210
rect 10980 3110 11010 3150
rect 11050 3110 11080 3150
rect 10980 3050 11080 3110
rect 10980 3010 11010 3050
rect 11050 3010 11080 3050
rect 10980 2980 11080 3010
rect 2140 2900 2220 2930
rect 2140 2860 2160 2900
rect 2200 2860 2220 2900
rect 2140 2800 2220 2860
rect 2140 2760 2160 2800
rect 2200 2760 2220 2800
rect 2140 2730 2220 2760
rect 2250 2900 2330 2930
rect 2250 2860 2270 2900
rect 2310 2860 2330 2900
rect 2250 2800 2330 2860
rect 2250 2760 2270 2800
rect 2310 2760 2330 2800
rect 2250 2730 2330 2760
rect 2360 2900 2440 2930
rect 2360 2860 2380 2900
rect 2420 2860 2440 2900
rect 2360 2800 2440 2860
rect 2360 2760 2380 2800
rect 2420 2760 2440 2800
rect 2360 2730 2440 2760
rect 2660 2900 2740 2930
rect 2660 2860 2680 2900
rect 2720 2860 2740 2900
rect 2660 2800 2740 2860
rect 2660 2760 2680 2800
rect 2720 2760 2740 2800
rect 2660 2730 2740 2760
rect 2770 2900 2850 2930
rect 2770 2860 2790 2900
rect 2830 2860 2850 2900
rect 2770 2800 2850 2860
rect 2770 2760 2790 2800
rect 2830 2760 2850 2800
rect 2770 2730 2850 2760
rect 2880 2900 2960 2930
rect 3040 2900 3120 2930
rect 2880 2860 2900 2900
rect 2940 2860 2960 2900
rect 3040 2860 3060 2900
rect 3100 2860 3120 2900
rect 2880 2800 2960 2860
rect 3040 2800 3120 2860
rect 2880 2760 2900 2800
rect 2940 2760 2960 2800
rect 3040 2760 3060 2800
rect 3100 2760 3120 2800
rect 2880 2730 2960 2760
rect 3040 2730 3120 2760
rect 3150 2900 3230 2930
rect 3150 2860 3170 2900
rect 3210 2860 3230 2900
rect 3150 2800 3230 2860
rect 3150 2760 3170 2800
rect 3210 2760 3230 2800
rect 3150 2730 3230 2760
rect 3260 2900 3340 2930
rect 3260 2860 3280 2900
rect 3320 2860 3340 2900
rect 3260 2800 3340 2860
rect 3260 2760 3280 2800
rect 3320 2760 3340 2800
rect 3260 2730 3340 2760
rect 3560 2900 3640 2930
rect 3560 2860 3580 2900
rect 3620 2860 3640 2900
rect 3560 2800 3640 2860
rect 3560 2760 3580 2800
rect 3620 2760 3640 2800
rect 3560 2730 3640 2760
rect 3670 2900 3750 2930
rect 3670 2860 3690 2900
rect 3730 2860 3750 2900
rect 3670 2800 3750 2860
rect 3670 2760 3690 2800
rect 3730 2760 3750 2800
rect 3670 2730 3750 2760
rect 3780 2900 3860 2930
rect 3780 2860 3800 2900
rect 3840 2860 3860 2900
rect 3780 2800 3860 2860
rect 3780 2760 3800 2800
rect 3840 2760 3860 2800
rect 3780 2730 3860 2760
rect 4070 2900 4150 2930
rect 4070 2860 4090 2900
rect 4130 2860 4150 2900
rect 4070 2800 4150 2860
rect 4070 2760 4090 2800
rect 4130 2760 4150 2800
rect 4070 2730 4150 2760
rect 4180 2900 4260 2930
rect 4180 2860 4200 2900
rect 4240 2860 4260 2900
rect 4180 2800 4260 2860
rect 4180 2760 4200 2800
rect 4240 2760 4260 2800
rect 4180 2730 4260 2760
rect 4400 2900 4480 2930
rect 4400 2860 4420 2900
rect 4460 2860 4480 2900
rect 4400 2800 4480 2860
rect 4400 2760 4420 2800
rect 4460 2760 4480 2800
rect 4400 2730 4480 2760
rect 4510 2900 4590 2930
rect 4510 2860 4530 2900
rect 4570 2860 4590 2900
rect 4510 2800 4590 2860
rect 4510 2760 4530 2800
rect 4570 2760 4590 2800
rect 4510 2730 4590 2760
rect 4730 2900 4810 2930
rect 4730 2860 4750 2900
rect 4790 2860 4810 2900
rect 4730 2800 4810 2860
rect 4730 2760 4750 2800
rect 4790 2760 4810 2800
rect 4730 2730 4810 2760
rect 4840 2900 4920 2930
rect 4840 2860 4860 2900
rect 4900 2860 4920 2900
rect 4840 2800 4920 2860
rect 4840 2760 4860 2800
rect 4900 2760 4920 2800
rect 4840 2730 4920 2760
rect 5270 2900 5370 2930
rect 5270 2860 5300 2900
rect 5340 2860 5370 2900
rect 5270 2800 5370 2860
rect 5270 2760 5300 2800
rect 5340 2760 5370 2800
rect 5270 2730 5370 2760
rect 5400 2900 5500 2930
rect 5400 2860 5430 2900
rect 5470 2860 5500 2900
rect 5400 2800 5500 2860
rect 5400 2760 5430 2800
rect 5470 2760 5500 2800
rect 5400 2730 5500 2760
rect 5660 2900 5760 2930
rect 5660 2860 5690 2900
rect 5730 2860 5760 2900
rect 5660 2800 5760 2860
rect 5660 2760 5690 2800
rect 5730 2760 5760 2800
rect 5660 2730 5760 2760
rect 5790 2900 5890 2930
rect 5790 2860 5820 2900
rect 5860 2860 5890 2900
rect 5790 2800 5890 2860
rect 5790 2760 5820 2800
rect 5860 2760 5890 2800
rect 5790 2730 5890 2760
rect 6050 2900 6150 2930
rect 6050 2860 6080 2900
rect 6120 2860 6150 2900
rect 6050 2800 6150 2860
rect 6050 2760 6080 2800
rect 6120 2760 6150 2800
rect 6050 2730 6150 2760
rect 6180 2900 6280 2930
rect 6180 2860 6210 2900
rect 6250 2860 6280 2900
rect 6180 2800 6280 2860
rect 6180 2760 6210 2800
rect 6250 2760 6280 2800
rect 6180 2730 6280 2760
rect 6340 2900 6440 2930
rect 6340 2860 6370 2900
rect 6410 2860 6440 2900
rect 6340 2800 6440 2860
rect 6340 2760 6370 2800
rect 6410 2760 6440 2800
rect 6340 2730 6440 2760
rect 6470 2900 6570 2930
rect 6470 2860 6500 2900
rect 6540 2860 6570 2900
rect 6470 2800 6570 2860
rect 6470 2760 6500 2800
rect 6540 2760 6570 2800
rect 6470 2730 6570 2760
rect 6730 2900 6830 2930
rect 6730 2860 6760 2900
rect 6800 2860 6830 2900
rect 6730 2800 6830 2860
rect 6730 2760 6760 2800
rect 6800 2760 6830 2800
rect 6730 2730 6830 2760
rect 6860 2900 6960 2930
rect 6860 2860 6890 2900
rect 6930 2860 6960 2900
rect 6860 2800 6960 2860
rect 6860 2760 6890 2800
rect 6930 2760 6960 2800
rect 6860 2730 6960 2760
rect 12400 1970 12480 2000
rect 12400 1930 12420 1970
rect 12460 1930 12480 1970
rect 12400 1870 12480 1930
rect 12400 1830 12420 1870
rect 12460 1830 12480 1870
rect 12400 1800 12480 1830
rect 12510 1970 12590 2000
rect 12510 1930 12530 1970
rect 12570 1930 12590 1970
rect 12510 1870 12590 1930
rect 12510 1830 12530 1870
rect 12570 1830 12590 1870
rect 12510 1800 12590 1830
rect 13000 1970 13080 2000
rect 13000 1930 13020 1970
rect 13060 1930 13080 1970
rect 13000 1870 13080 1930
rect 13000 1830 13020 1870
rect 13060 1830 13080 1870
rect 13000 1800 13080 1830
rect 13110 1970 13190 2000
rect 13110 1930 13130 1970
rect 13170 1930 13190 1970
rect 13110 1870 13190 1930
rect 13110 1830 13130 1870
rect 13170 1830 13190 1870
rect 13110 1800 13190 1830
rect 13600 1970 13680 2000
rect 13600 1930 13620 1970
rect 13660 1930 13680 1970
rect 13600 1870 13680 1930
rect 13600 1830 13620 1870
rect 13660 1830 13680 1870
rect 13600 1800 13680 1830
rect 13710 1970 13790 2000
rect 13870 1970 13950 2000
rect 13710 1930 13730 1970
rect 13770 1930 13790 1970
rect 13870 1930 13890 1970
rect 13930 1930 13950 1970
rect 13710 1870 13790 1930
rect 13870 1870 13950 1930
rect 13710 1830 13730 1870
rect 13770 1830 13790 1870
rect 13870 1830 13890 1870
rect 13930 1830 13950 1870
rect 13710 1800 13790 1830
rect 13870 1800 13950 1830
rect 13980 1970 14060 2000
rect 13980 1930 14000 1970
rect 14040 1930 14060 1970
rect 13980 1870 14060 1930
rect 13980 1830 14000 1870
rect 14040 1830 14060 1870
rect 13980 1800 14060 1830
rect 12400 1640 12480 1670
rect 12400 1600 12420 1640
rect 12460 1600 12480 1640
rect 12400 1570 12480 1600
rect 12510 1640 12590 1670
rect 12510 1600 12530 1640
rect 12570 1600 12590 1640
rect 12510 1570 12590 1600
rect 13000 1640 13080 1670
rect 13000 1600 13020 1640
rect 13060 1600 13080 1640
rect 13000 1570 13080 1600
rect 13110 1640 13190 1670
rect 13110 1600 13130 1640
rect 13170 1600 13190 1640
rect 13110 1570 13190 1600
rect 13600 1640 13680 1670
rect 13600 1600 13620 1640
rect 13660 1600 13680 1640
rect 13600 1570 13680 1600
rect 13710 1640 13790 1670
rect 13710 1600 13730 1640
rect 13770 1600 13790 1640
rect 13710 1570 13790 1600
rect 1830 1410 1910 1440
rect 1830 1370 1850 1410
rect 1890 1370 1910 1410
rect 1830 1340 1910 1370
rect 1940 1410 2020 1440
rect 1940 1370 1960 1410
rect 2000 1370 2020 1410
rect 1940 1340 2020 1370
rect 2050 1410 2130 1440
rect 2050 1370 2070 1410
rect 2110 1370 2130 1410
rect 2050 1340 2130 1370
rect 2160 1410 2240 1440
rect 2160 1370 2180 1410
rect 2220 1370 2240 1410
rect 2160 1340 2240 1370
rect 2270 1410 2350 1440
rect 2270 1370 2290 1410
rect 2330 1370 2350 1410
rect 2270 1340 2350 1370
rect 2410 1410 2490 1440
rect 2410 1370 2430 1410
rect 2470 1370 2490 1410
rect 2410 1340 2490 1370
rect 2520 1410 2600 1440
rect 2520 1370 2540 1410
rect 2580 1370 2600 1410
rect 2520 1340 2600 1370
rect 2630 1410 2710 1440
rect 2630 1370 2650 1410
rect 2690 1370 2710 1410
rect 2630 1340 2710 1370
rect 2860 1410 2940 1440
rect 2860 1370 2880 1410
rect 2920 1370 2940 1410
rect 2860 1340 2940 1370
rect 2970 1410 3050 1440
rect 2970 1370 2990 1410
rect 3030 1370 3050 1410
rect 2970 1340 3050 1370
rect 3080 1410 3160 1440
rect 3080 1370 3100 1410
rect 3140 1370 3160 1410
rect 3080 1340 3160 1370
rect 3190 1410 3270 1440
rect 3190 1370 3210 1410
rect 3250 1370 3270 1410
rect 3190 1340 3270 1370
rect 3300 1410 3380 1440
rect 3300 1370 3320 1410
rect 3360 1370 3380 1410
rect 3300 1340 3380 1370
rect 3520 1410 3600 1440
rect 3520 1370 3540 1410
rect 3580 1370 3600 1410
rect 3520 1340 3600 1370
rect 3630 1410 3710 1440
rect 3630 1370 3650 1410
rect 3690 1370 3710 1410
rect 3630 1340 3710 1370
rect 3740 1410 3820 1440
rect 3740 1370 3760 1410
rect 3800 1370 3820 1410
rect 3740 1340 3820 1370
rect 3850 1410 3930 1440
rect 3850 1370 3870 1410
rect 3910 1370 3930 1410
rect 3850 1340 3930 1370
rect 3960 1410 4040 1440
rect 3960 1370 3980 1410
rect 4020 1370 4040 1410
rect 3960 1340 4040 1370
rect 4200 1410 4280 1440
rect 4200 1370 4220 1410
rect 4260 1370 4280 1410
rect 4200 1340 4280 1370
rect 4310 1410 4390 1440
rect 4310 1370 4330 1410
rect 4370 1370 4390 1410
rect 4310 1340 4390 1370
rect 4420 1410 4500 1440
rect 4420 1370 4440 1410
rect 4480 1370 4500 1410
rect 4420 1340 4500 1370
rect 4530 1410 4610 1440
rect 4530 1370 4550 1410
rect 4590 1370 4610 1410
rect 4530 1340 4610 1370
rect 4640 1410 4720 1440
rect 4640 1370 4660 1410
rect 4700 1370 4720 1410
rect 4640 1340 4720 1370
rect 4780 1410 4860 1440
rect 4780 1370 4800 1410
rect 4840 1370 4860 1410
rect 4780 1340 4860 1370
rect 4890 1410 4970 1440
rect 4890 1370 4910 1410
rect 4950 1370 4970 1410
rect 4890 1340 4970 1370
rect 5000 1410 5080 1440
rect 5000 1370 5020 1410
rect 5060 1370 5080 1410
rect 5000 1340 5080 1370
rect 5340 1410 5420 1440
rect 5340 1370 5360 1410
rect 5400 1370 5420 1410
rect 5340 1340 5420 1370
rect 5450 1410 5530 1440
rect 5450 1370 5470 1410
rect 5510 1370 5530 1410
rect 5450 1340 5530 1370
rect 5700 1410 5780 1440
rect 5700 1370 5720 1410
rect 5760 1370 5780 1410
rect 5700 1340 5780 1370
rect 5810 1410 5890 1440
rect 5810 1370 5830 1410
rect 5870 1370 5890 1410
rect 5810 1340 5890 1370
rect 5950 1410 6030 1440
rect 5950 1370 5970 1410
rect 6010 1370 6030 1410
rect 5950 1340 6030 1370
rect 6060 1410 6140 1440
rect 6060 1370 6080 1410
rect 6120 1370 6140 1410
rect 6060 1340 6140 1370
rect 6170 1410 6250 1440
rect 6170 1370 6190 1410
rect 6230 1370 6250 1410
rect 6170 1340 6250 1370
rect 6280 1410 6360 1440
rect 6280 1370 6300 1410
rect 6340 1370 6360 1410
rect 6280 1340 6360 1370
rect 6390 1410 6470 1440
rect 6390 1370 6410 1410
rect 6450 1370 6470 1410
rect 6390 1340 6470 1370
rect 6610 1410 6690 1440
rect 6610 1370 6630 1410
rect 6670 1370 6690 1410
rect 6610 1340 6690 1370
rect 6720 1410 6800 1440
rect 6720 1370 6740 1410
rect 6780 1370 6800 1410
rect 6720 1340 6800 1370
rect 6830 1410 6910 1440
rect 6830 1370 6850 1410
rect 6890 1370 6910 1410
rect 6830 1340 6910 1370
rect 6940 1410 7020 1440
rect 6940 1370 6960 1410
rect 7000 1370 7020 1410
rect 6940 1340 7020 1370
rect 7160 1410 7240 1440
rect 7160 1370 7180 1410
rect 7220 1370 7240 1410
rect 7160 1340 7240 1370
rect 7270 1410 7350 1440
rect 7270 1370 7290 1410
rect 7330 1370 7350 1410
rect 7270 1340 7350 1370
rect 7380 1410 7460 1440
rect 7380 1370 7400 1410
rect 7440 1370 7460 1410
rect 7380 1340 7460 1370
rect 7490 1410 7570 1440
rect 7490 1370 7510 1410
rect 7550 1370 7570 1410
rect 7490 1340 7570 1370
rect 7600 1410 7680 1440
rect 7600 1370 7620 1410
rect 7660 1370 7680 1410
rect 7600 1340 7680 1370
rect 7820 1410 7900 1440
rect 7820 1370 7840 1410
rect 7880 1370 7900 1410
rect 7820 1340 7900 1370
rect 7930 1410 8010 1440
rect 7930 1370 7950 1410
rect 7990 1370 8010 1410
rect 7930 1340 8010 1370
rect 8040 1410 8120 1440
rect 8040 1370 8060 1410
rect 8100 1370 8120 1410
rect 8040 1340 8120 1370
rect 8150 1410 8230 1440
rect 8460 1500 8540 1530
rect 8460 1460 8480 1500
rect 8520 1460 8540 1500
rect 8460 1430 8540 1460
rect 8570 1500 8650 1530
rect 8570 1460 8590 1500
rect 8630 1460 8650 1500
rect 8570 1430 8650 1460
rect 8680 1500 8760 1530
rect 8680 1460 8700 1500
rect 8740 1460 8760 1500
rect 8680 1430 8760 1460
rect 8790 1500 8870 1530
rect 8790 1460 8810 1500
rect 8850 1460 8870 1500
rect 8790 1430 8870 1460
rect 8900 1500 8980 1530
rect 8900 1460 8920 1500
rect 8960 1460 8980 1500
rect 8900 1430 8980 1460
rect 9120 1500 9200 1530
rect 9120 1460 9140 1500
rect 9180 1460 9200 1500
rect 9120 1430 9200 1460
rect 9230 1500 9310 1530
rect 9230 1460 9250 1500
rect 9290 1460 9310 1500
rect 9230 1430 9310 1460
rect 9340 1500 9420 1530
rect 9340 1460 9360 1500
rect 9400 1460 9420 1500
rect 9340 1430 9420 1460
rect 9450 1500 9530 1530
rect 9450 1460 9470 1500
rect 9510 1460 9530 1500
rect 9450 1430 9530 1460
rect 9760 1500 9840 1530
rect 9760 1460 9780 1500
rect 9820 1460 9840 1500
rect 9760 1430 9840 1460
rect 9870 1500 9950 1530
rect 9870 1460 9890 1500
rect 9930 1460 9950 1500
rect 9870 1430 9950 1460
rect 9980 1500 10060 1530
rect 9980 1460 10000 1500
rect 10040 1460 10060 1500
rect 9980 1430 10060 1460
rect 10090 1500 10170 1530
rect 10090 1460 10110 1500
rect 10150 1460 10170 1500
rect 10090 1430 10170 1460
rect 10200 1500 10280 1530
rect 10200 1460 10220 1500
rect 10260 1460 10280 1500
rect 10200 1430 10280 1460
rect 10420 1500 10500 1530
rect 10420 1460 10440 1500
rect 10480 1460 10500 1500
rect 10420 1430 10500 1460
rect 10530 1500 10610 1530
rect 10530 1460 10550 1500
rect 10590 1460 10610 1500
rect 10530 1430 10610 1460
rect 10640 1500 10720 1530
rect 10640 1460 10660 1500
rect 10700 1460 10720 1500
rect 10640 1430 10720 1460
rect 10750 1500 10830 1530
rect 10750 1460 10770 1500
rect 10810 1460 10830 1500
rect 10750 1430 10830 1460
rect 11060 1500 11140 1530
rect 11060 1460 11080 1500
rect 11120 1460 11140 1500
rect 11060 1430 11140 1460
rect 11170 1500 11250 1530
rect 11170 1460 11190 1500
rect 11230 1460 11250 1500
rect 11170 1430 11250 1460
rect 11280 1500 11360 1530
rect 11280 1460 11300 1500
rect 11340 1460 11360 1500
rect 11280 1430 11360 1460
rect 11390 1500 11470 1530
rect 11390 1460 11410 1500
rect 11450 1460 11470 1500
rect 11390 1430 11470 1460
rect 11500 1500 11580 1530
rect 11500 1460 11520 1500
rect 11560 1460 11580 1500
rect 11500 1430 11580 1460
rect 11720 1500 11800 1530
rect 11720 1460 11740 1500
rect 11780 1460 11800 1500
rect 11720 1430 11800 1460
rect 11830 1500 11910 1530
rect 11830 1460 11850 1500
rect 11890 1460 11910 1500
rect 11830 1430 11910 1460
rect 11940 1500 12020 1530
rect 11940 1460 11960 1500
rect 12000 1460 12020 1500
rect 11940 1430 12020 1460
rect 12050 1500 12130 1530
rect 12050 1460 12070 1500
rect 12110 1460 12130 1500
rect 12050 1430 12130 1460
rect 8150 1370 8170 1410
rect 8210 1370 8230 1410
rect 8150 1340 8230 1370
rect 12400 1400 12480 1430
rect 12400 1360 12420 1400
rect 12460 1360 12480 1400
rect 12400 1330 12480 1360
rect 12510 1400 12590 1430
rect 12510 1360 12530 1400
rect 12570 1360 12590 1400
rect 12510 1330 12590 1360
rect 13000 1400 13080 1430
rect 13000 1360 13020 1400
rect 13060 1360 13080 1400
rect 13000 1330 13080 1360
rect 13110 1400 13190 1430
rect 13110 1360 13130 1400
rect 13170 1360 13190 1400
rect 13110 1330 13190 1360
rect 13600 1400 13680 1430
rect 13600 1360 13620 1400
rect 13660 1360 13680 1400
rect 13600 1330 13680 1360
rect 13710 1400 13790 1430
rect 13710 1360 13730 1400
rect 13770 1360 13790 1400
rect 13710 1330 13790 1360
<< pdiff >>
rect 1570 14436 2250 14490
rect 1570 14402 1622 14436
rect 1656 14402 1712 14436
rect 1746 14402 1802 14436
rect 1836 14402 1892 14436
rect 1926 14402 1982 14436
rect 2016 14402 2072 14436
rect 2106 14402 2162 14436
rect 2196 14402 2250 14436
rect 1570 14346 2250 14402
rect 1570 14312 1622 14346
rect 1656 14312 1712 14346
rect 1746 14312 1802 14346
rect 1836 14312 1892 14346
rect 1926 14312 1982 14346
rect 2016 14312 2072 14346
rect 2106 14312 2162 14346
rect 2196 14312 2250 14346
rect 1570 14256 2250 14312
rect 1570 14222 1622 14256
rect 1656 14222 1712 14256
rect 1746 14222 1802 14256
rect 1836 14222 1892 14256
rect 1926 14222 1982 14256
rect 2016 14222 2072 14256
rect 2106 14222 2162 14256
rect 2196 14222 2250 14256
rect 1570 14166 2250 14222
rect 1570 14132 1622 14166
rect 1656 14132 1712 14166
rect 1746 14132 1802 14166
rect 1836 14132 1892 14166
rect 1926 14132 1982 14166
rect 2016 14132 2072 14166
rect 2106 14132 2162 14166
rect 2196 14132 2250 14166
rect 1570 14076 2250 14132
rect 1570 14042 1622 14076
rect 1656 14042 1712 14076
rect 1746 14042 1802 14076
rect 1836 14042 1892 14076
rect 1926 14042 1982 14076
rect 2016 14042 2072 14076
rect 2106 14042 2162 14076
rect 2196 14042 2250 14076
rect 1570 13986 2250 14042
rect 1570 13952 1622 13986
rect 1656 13952 1712 13986
rect 1746 13952 1802 13986
rect 1836 13952 1892 13986
rect 1926 13952 1982 13986
rect 2016 13952 2072 13986
rect 2106 13952 2162 13986
rect 2196 13952 2250 13986
rect 1570 13896 2250 13952
rect 1570 13862 1622 13896
rect 1656 13862 1712 13896
rect 1746 13862 1802 13896
rect 1836 13862 1892 13896
rect 1926 13862 1982 13896
rect 2016 13862 2072 13896
rect 2106 13862 2162 13896
rect 2196 13862 2250 13896
rect 1570 13810 2250 13862
rect 2930 14436 3610 14490
rect 2930 14402 2982 14436
rect 3016 14402 3072 14436
rect 3106 14402 3162 14436
rect 3196 14402 3252 14436
rect 3286 14402 3342 14436
rect 3376 14402 3432 14436
rect 3466 14402 3522 14436
rect 3556 14402 3610 14436
rect 2930 14346 3610 14402
rect 2930 14312 2982 14346
rect 3016 14312 3072 14346
rect 3106 14312 3162 14346
rect 3196 14312 3252 14346
rect 3286 14312 3342 14346
rect 3376 14312 3432 14346
rect 3466 14312 3522 14346
rect 3556 14312 3610 14346
rect 2930 14256 3610 14312
rect 2930 14222 2982 14256
rect 3016 14222 3072 14256
rect 3106 14222 3162 14256
rect 3196 14222 3252 14256
rect 3286 14222 3342 14256
rect 3376 14222 3432 14256
rect 3466 14222 3522 14256
rect 3556 14222 3610 14256
rect 2930 14166 3610 14222
rect 2930 14132 2982 14166
rect 3016 14132 3072 14166
rect 3106 14132 3162 14166
rect 3196 14132 3252 14166
rect 3286 14132 3342 14166
rect 3376 14132 3432 14166
rect 3466 14132 3522 14166
rect 3556 14132 3610 14166
rect 2930 14076 3610 14132
rect 2930 14042 2982 14076
rect 3016 14042 3072 14076
rect 3106 14042 3162 14076
rect 3196 14042 3252 14076
rect 3286 14042 3342 14076
rect 3376 14042 3432 14076
rect 3466 14042 3522 14076
rect 3556 14042 3610 14076
rect 2930 13986 3610 14042
rect 2930 13952 2982 13986
rect 3016 13952 3072 13986
rect 3106 13952 3162 13986
rect 3196 13952 3252 13986
rect 3286 13952 3342 13986
rect 3376 13952 3432 13986
rect 3466 13952 3522 13986
rect 3556 13952 3610 13986
rect 2930 13896 3610 13952
rect 2930 13862 2982 13896
rect 3016 13862 3072 13896
rect 3106 13862 3162 13896
rect 3196 13862 3252 13896
rect 3286 13862 3342 13896
rect 3376 13862 3432 13896
rect 3466 13862 3522 13896
rect 3556 13862 3610 13896
rect 2930 13810 3610 13862
rect 4290 14436 4970 14490
rect 4290 14402 4342 14436
rect 4376 14402 4432 14436
rect 4466 14402 4522 14436
rect 4556 14402 4612 14436
rect 4646 14402 4702 14436
rect 4736 14402 4792 14436
rect 4826 14402 4882 14436
rect 4916 14402 4970 14436
rect 4290 14346 4970 14402
rect 4290 14312 4342 14346
rect 4376 14312 4432 14346
rect 4466 14312 4522 14346
rect 4556 14312 4612 14346
rect 4646 14312 4702 14346
rect 4736 14312 4792 14346
rect 4826 14312 4882 14346
rect 4916 14312 4970 14346
rect 4290 14256 4970 14312
rect 4290 14222 4342 14256
rect 4376 14222 4432 14256
rect 4466 14222 4522 14256
rect 4556 14222 4612 14256
rect 4646 14222 4702 14256
rect 4736 14222 4792 14256
rect 4826 14222 4882 14256
rect 4916 14222 4970 14256
rect 4290 14166 4970 14222
rect 4290 14132 4342 14166
rect 4376 14132 4432 14166
rect 4466 14132 4522 14166
rect 4556 14132 4612 14166
rect 4646 14132 4702 14166
rect 4736 14132 4792 14166
rect 4826 14132 4882 14166
rect 4916 14132 4970 14166
rect 4290 14076 4970 14132
rect 4290 14042 4342 14076
rect 4376 14042 4432 14076
rect 4466 14042 4522 14076
rect 4556 14042 4612 14076
rect 4646 14042 4702 14076
rect 4736 14042 4792 14076
rect 4826 14042 4882 14076
rect 4916 14042 4970 14076
rect 4290 13986 4970 14042
rect 4290 13952 4342 13986
rect 4376 13952 4432 13986
rect 4466 13952 4522 13986
rect 4556 13952 4612 13986
rect 4646 13952 4702 13986
rect 4736 13952 4792 13986
rect 4826 13952 4882 13986
rect 4916 13952 4970 13986
rect 4290 13896 4970 13952
rect 4290 13862 4342 13896
rect 4376 13862 4432 13896
rect 4466 13862 4522 13896
rect 4556 13862 4612 13896
rect 4646 13862 4702 13896
rect 4736 13862 4792 13896
rect 4826 13862 4882 13896
rect 4916 13862 4970 13896
rect 4290 13810 4970 13862
rect 1570 13076 2250 13130
rect 1570 13042 1622 13076
rect 1656 13042 1712 13076
rect 1746 13042 1802 13076
rect 1836 13042 1892 13076
rect 1926 13042 1982 13076
rect 2016 13042 2072 13076
rect 2106 13042 2162 13076
rect 2196 13042 2250 13076
rect 1570 12986 2250 13042
rect 1570 12952 1622 12986
rect 1656 12952 1712 12986
rect 1746 12952 1802 12986
rect 1836 12952 1892 12986
rect 1926 12952 1982 12986
rect 2016 12952 2072 12986
rect 2106 12952 2162 12986
rect 2196 12952 2250 12986
rect 1570 12896 2250 12952
rect 1570 12862 1622 12896
rect 1656 12862 1712 12896
rect 1746 12862 1802 12896
rect 1836 12862 1892 12896
rect 1926 12862 1982 12896
rect 2016 12862 2072 12896
rect 2106 12862 2162 12896
rect 2196 12862 2250 12896
rect 1570 12806 2250 12862
rect 1570 12772 1622 12806
rect 1656 12772 1712 12806
rect 1746 12772 1802 12806
rect 1836 12772 1892 12806
rect 1926 12772 1982 12806
rect 2016 12772 2072 12806
rect 2106 12772 2162 12806
rect 2196 12772 2250 12806
rect 1570 12716 2250 12772
rect 1570 12682 1622 12716
rect 1656 12682 1712 12716
rect 1746 12682 1802 12716
rect 1836 12682 1892 12716
rect 1926 12682 1982 12716
rect 2016 12682 2072 12716
rect 2106 12682 2162 12716
rect 2196 12682 2250 12716
rect 1570 12626 2250 12682
rect 1570 12592 1622 12626
rect 1656 12592 1712 12626
rect 1746 12592 1802 12626
rect 1836 12592 1892 12626
rect 1926 12592 1982 12626
rect 2016 12592 2072 12626
rect 2106 12592 2162 12626
rect 2196 12592 2250 12626
rect 1570 12536 2250 12592
rect 1570 12502 1622 12536
rect 1656 12502 1712 12536
rect 1746 12502 1802 12536
rect 1836 12502 1892 12536
rect 1926 12502 1982 12536
rect 2016 12502 2072 12536
rect 2106 12502 2162 12536
rect 2196 12502 2250 12536
rect 1570 12450 2250 12502
rect 2930 13076 3610 13130
rect 2930 13042 2982 13076
rect 3016 13042 3072 13076
rect 3106 13042 3162 13076
rect 3196 13042 3252 13076
rect 3286 13042 3342 13076
rect 3376 13042 3432 13076
rect 3466 13042 3522 13076
rect 3556 13042 3610 13076
rect 2930 12986 3610 13042
rect 2930 12952 2982 12986
rect 3016 12952 3072 12986
rect 3106 12952 3162 12986
rect 3196 12952 3252 12986
rect 3286 12952 3342 12986
rect 3376 12952 3432 12986
rect 3466 12952 3522 12986
rect 3556 12952 3610 12986
rect 2930 12896 3610 12952
rect 2930 12862 2982 12896
rect 3016 12862 3072 12896
rect 3106 12862 3162 12896
rect 3196 12862 3252 12896
rect 3286 12862 3342 12896
rect 3376 12862 3432 12896
rect 3466 12862 3522 12896
rect 3556 12862 3610 12896
rect 2930 12806 3610 12862
rect 2930 12772 2982 12806
rect 3016 12772 3072 12806
rect 3106 12772 3162 12806
rect 3196 12772 3252 12806
rect 3286 12772 3342 12806
rect 3376 12772 3432 12806
rect 3466 12772 3522 12806
rect 3556 12772 3610 12806
rect 2930 12716 3610 12772
rect 2930 12682 2982 12716
rect 3016 12682 3072 12716
rect 3106 12682 3162 12716
rect 3196 12682 3252 12716
rect 3286 12682 3342 12716
rect 3376 12682 3432 12716
rect 3466 12682 3522 12716
rect 3556 12682 3610 12716
rect 2930 12626 3610 12682
rect 2930 12592 2982 12626
rect 3016 12592 3072 12626
rect 3106 12592 3162 12626
rect 3196 12592 3252 12626
rect 3286 12592 3342 12626
rect 3376 12592 3432 12626
rect 3466 12592 3522 12626
rect 3556 12592 3610 12626
rect 2930 12536 3610 12592
rect 2930 12502 2982 12536
rect 3016 12502 3072 12536
rect 3106 12502 3162 12536
rect 3196 12502 3252 12536
rect 3286 12502 3342 12536
rect 3376 12502 3432 12536
rect 3466 12502 3522 12536
rect 3556 12502 3610 12536
rect 2930 12450 3610 12502
rect 4290 13076 4970 13130
rect 4290 13042 4342 13076
rect 4376 13042 4432 13076
rect 4466 13042 4522 13076
rect 4556 13042 4612 13076
rect 4646 13042 4702 13076
rect 4736 13042 4792 13076
rect 4826 13042 4882 13076
rect 4916 13042 4970 13076
rect 4290 12986 4970 13042
rect 4290 12952 4342 12986
rect 4376 12952 4432 12986
rect 4466 12952 4522 12986
rect 4556 12952 4612 12986
rect 4646 12952 4702 12986
rect 4736 12952 4792 12986
rect 4826 12952 4882 12986
rect 4916 12952 4970 12986
rect 4290 12896 4970 12952
rect 4290 12862 4342 12896
rect 4376 12862 4432 12896
rect 4466 12862 4522 12896
rect 4556 12862 4612 12896
rect 4646 12862 4702 12896
rect 4736 12862 4792 12896
rect 4826 12862 4882 12896
rect 4916 12862 4970 12896
rect 4290 12806 4970 12862
rect 4290 12772 4342 12806
rect 4376 12772 4432 12806
rect 4466 12772 4522 12806
rect 4556 12772 4612 12806
rect 4646 12772 4702 12806
rect 4736 12772 4792 12806
rect 4826 12772 4882 12806
rect 4916 12772 4970 12806
rect 4290 12716 4970 12772
rect 4290 12682 4342 12716
rect 4376 12682 4432 12716
rect 4466 12682 4522 12716
rect 4556 12682 4612 12716
rect 4646 12682 4702 12716
rect 4736 12682 4792 12716
rect 4826 12682 4882 12716
rect 4916 12682 4970 12716
rect 4290 12626 4970 12682
rect 4290 12592 4342 12626
rect 4376 12592 4432 12626
rect 4466 12592 4522 12626
rect 4556 12592 4612 12626
rect 4646 12592 4702 12626
rect 4736 12592 4792 12626
rect 4826 12592 4882 12626
rect 4916 12592 4970 12626
rect 4290 12536 4970 12592
rect 4290 12502 4342 12536
rect 4376 12502 4432 12536
rect 4466 12502 4522 12536
rect 4556 12502 4612 12536
rect 4646 12502 4702 12536
rect 4736 12502 4792 12536
rect 4826 12502 4882 12536
rect 4916 12502 4970 12536
rect 4290 12450 4970 12502
rect 1570 11716 2250 11770
rect 1570 11682 1622 11716
rect 1656 11682 1712 11716
rect 1746 11682 1802 11716
rect 1836 11682 1892 11716
rect 1926 11682 1982 11716
rect 2016 11682 2072 11716
rect 2106 11682 2162 11716
rect 2196 11682 2250 11716
rect 1570 11626 2250 11682
rect 1570 11592 1622 11626
rect 1656 11592 1712 11626
rect 1746 11592 1802 11626
rect 1836 11592 1892 11626
rect 1926 11592 1982 11626
rect 2016 11592 2072 11626
rect 2106 11592 2162 11626
rect 2196 11592 2250 11626
rect 1570 11536 2250 11592
rect 1570 11502 1622 11536
rect 1656 11502 1712 11536
rect 1746 11502 1802 11536
rect 1836 11502 1892 11536
rect 1926 11502 1982 11536
rect 2016 11502 2072 11536
rect 2106 11502 2162 11536
rect 2196 11502 2250 11536
rect 1570 11446 2250 11502
rect 1570 11412 1622 11446
rect 1656 11412 1712 11446
rect 1746 11412 1802 11446
rect 1836 11412 1892 11446
rect 1926 11412 1982 11446
rect 2016 11412 2072 11446
rect 2106 11412 2162 11446
rect 2196 11412 2250 11446
rect 1570 11356 2250 11412
rect 1570 11322 1622 11356
rect 1656 11322 1712 11356
rect 1746 11322 1802 11356
rect 1836 11322 1892 11356
rect 1926 11322 1982 11356
rect 2016 11322 2072 11356
rect 2106 11322 2162 11356
rect 2196 11322 2250 11356
rect 1570 11266 2250 11322
rect 1570 11232 1622 11266
rect 1656 11232 1712 11266
rect 1746 11232 1802 11266
rect 1836 11232 1892 11266
rect 1926 11232 1982 11266
rect 2016 11232 2072 11266
rect 2106 11232 2162 11266
rect 2196 11232 2250 11266
rect 1570 11176 2250 11232
rect 1570 11142 1622 11176
rect 1656 11142 1712 11176
rect 1746 11142 1802 11176
rect 1836 11142 1892 11176
rect 1926 11142 1982 11176
rect 2016 11142 2072 11176
rect 2106 11142 2162 11176
rect 2196 11142 2250 11176
rect 1570 11090 2250 11142
rect 2930 11716 3610 11770
rect 2930 11682 2982 11716
rect 3016 11682 3072 11716
rect 3106 11682 3162 11716
rect 3196 11682 3252 11716
rect 3286 11682 3342 11716
rect 3376 11682 3432 11716
rect 3466 11682 3522 11716
rect 3556 11682 3610 11716
rect 2930 11626 3610 11682
rect 2930 11592 2982 11626
rect 3016 11592 3072 11626
rect 3106 11592 3162 11626
rect 3196 11592 3252 11626
rect 3286 11592 3342 11626
rect 3376 11592 3432 11626
rect 3466 11592 3522 11626
rect 3556 11592 3610 11626
rect 2930 11536 3610 11592
rect 2930 11502 2982 11536
rect 3016 11502 3072 11536
rect 3106 11502 3162 11536
rect 3196 11502 3252 11536
rect 3286 11502 3342 11536
rect 3376 11502 3432 11536
rect 3466 11502 3522 11536
rect 3556 11502 3610 11536
rect 2930 11446 3610 11502
rect 2930 11412 2982 11446
rect 3016 11412 3072 11446
rect 3106 11412 3162 11446
rect 3196 11412 3252 11446
rect 3286 11412 3342 11446
rect 3376 11412 3432 11446
rect 3466 11412 3522 11446
rect 3556 11412 3610 11446
rect 2930 11356 3610 11412
rect 2930 11322 2982 11356
rect 3016 11322 3072 11356
rect 3106 11322 3162 11356
rect 3196 11322 3252 11356
rect 3286 11322 3342 11356
rect 3376 11322 3432 11356
rect 3466 11322 3522 11356
rect 3556 11322 3610 11356
rect 2930 11266 3610 11322
rect 2930 11232 2982 11266
rect 3016 11232 3072 11266
rect 3106 11232 3162 11266
rect 3196 11232 3252 11266
rect 3286 11232 3342 11266
rect 3376 11232 3432 11266
rect 3466 11232 3522 11266
rect 3556 11232 3610 11266
rect 2930 11176 3610 11232
rect 2930 11142 2982 11176
rect 3016 11142 3072 11176
rect 3106 11142 3162 11176
rect 3196 11142 3252 11176
rect 3286 11142 3342 11176
rect 3376 11142 3432 11176
rect 3466 11142 3522 11176
rect 3556 11142 3610 11176
rect 2930 11090 3610 11142
rect 4290 11716 4970 11770
rect 4290 11682 4342 11716
rect 4376 11682 4432 11716
rect 4466 11682 4522 11716
rect 4556 11682 4612 11716
rect 4646 11682 4702 11716
rect 4736 11682 4792 11716
rect 4826 11682 4882 11716
rect 4916 11682 4970 11716
rect 4290 11626 4970 11682
rect 4290 11592 4342 11626
rect 4376 11592 4432 11626
rect 4466 11592 4522 11626
rect 4556 11592 4612 11626
rect 4646 11592 4702 11626
rect 4736 11592 4792 11626
rect 4826 11592 4882 11626
rect 4916 11592 4970 11626
rect 4290 11536 4970 11592
rect 4290 11502 4342 11536
rect 4376 11502 4432 11536
rect 4466 11502 4522 11536
rect 4556 11502 4612 11536
rect 4646 11502 4702 11536
rect 4736 11502 4792 11536
rect 4826 11502 4882 11536
rect 4916 11502 4970 11536
rect 4290 11446 4970 11502
rect 4290 11412 4342 11446
rect 4376 11412 4432 11446
rect 4466 11412 4522 11446
rect 4556 11412 4612 11446
rect 4646 11412 4702 11446
rect 4736 11412 4792 11446
rect 4826 11412 4882 11446
rect 4916 11412 4970 11446
rect 4290 11356 4970 11412
rect 4290 11322 4342 11356
rect 4376 11322 4432 11356
rect 4466 11322 4522 11356
rect 4556 11322 4612 11356
rect 4646 11322 4702 11356
rect 4736 11322 4792 11356
rect 4826 11322 4882 11356
rect 4916 11322 4970 11356
rect 4290 11266 4970 11322
rect 4290 11232 4342 11266
rect 4376 11232 4432 11266
rect 4466 11232 4522 11266
rect 4556 11232 4612 11266
rect 4646 11232 4702 11266
rect 4736 11232 4792 11266
rect 4826 11232 4882 11266
rect 4916 11232 4970 11266
rect 4290 11176 4970 11232
rect 4290 11142 4342 11176
rect 4376 11142 4432 11176
rect 4466 11142 4522 11176
rect 4556 11142 4612 11176
rect 4646 11142 4702 11176
rect 4736 11142 4792 11176
rect 4826 11142 4882 11176
rect 4916 11142 4970 11176
rect 4290 11090 4970 11142
rect 510 7800 590 7830
rect 510 7760 530 7800
rect 570 7760 590 7800
rect 510 7700 590 7760
rect 510 7660 530 7700
rect 570 7660 590 7700
rect 510 7630 590 7660
rect 630 7800 710 7830
rect 630 7760 650 7800
rect 690 7760 710 7800
rect 630 7700 710 7760
rect 630 7660 650 7700
rect 690 7660 710 7700
rect 630 7630 710 7660
rect 750 7800 830 7830
rect 750 7760 770 7800
rect 810 7760 830 7800
rect 750 7700 830 7760
rect 750 7660 770 7700
rect 810 7660 830 7700
rect 750 7630 830 7660
rect 870 7800 950 7830
rect 870 7760 890 7800
rect 930 7760 950 7800
rect 870 7700 950 7760
rect 870 7660 890 7700
rect 930 7660 950 7700
rect 870 7630 950 7660
rect 990 7800 1070 7830
rect 990 7760 1010 7800
rect 1050 7760 1070 7800
rect 990 7700 1070 7760
rect 990 7660 1010 7700
rect 1050 7660 1070 7700
rect 990 7630 1070 7660
rect 1110 7800 1190 7830
rect 1110 7760 1130 7800
rect 1170 7760 1190 7800
rect 1110 7700 1190 7760
rect 1110 7660 1130 7700
rect 1170 7660 1190 7700
rect 1110 7630 1190 7660
rect 1230 7800 1310 7830
rect 1230 7760 1250 7800
rect 1290 7760 1310 7800
rect 1230 7700 1310 7760
rect 1230 7660 1250 7700
rect 1290 7660 1310 7700
rect 1230 7630 1310 7660
rect 1350 7800 1430 7830
rect 1350 7760 1370 7800
rect 1410 7760 1430 7800
rect 1350 7700 1430 7760
rect 1350 7660 1370 7700
rect 1410 7660 1430 7700
rect 1350 7630 1430 7660
rect 1470 7800 1550 7830
rect 1470 7760 1490 7800
rect 1530 7760 1550 7800
rect 1470 7700 1550 7760
rect 1470 7660 1490 7700
rect 1530 7660 1550 7700
rect 1470 7630 1550 7660
rect 1590 7800 1670 7830
rect 1590 7760 1610 7800
rect 1650 7760 1670 7800
rect 1590 7700 1670 7760
rect 1590 7660 1610 7700
rect 1650 7660 1670 7700
rect 1590 7630 1670 7660
rect 1710 7800 1790 7830
rect 1710 7760 1730 7800
rect 1770 7760 1790 7800
rect 1710 7700 1790 7760
rect 1710 7660 1730 7700
rect 1770 7660 1790 7700
rect 1710 7630 1790 7660
rect 1830 7800 1910 7830
rect 1830 7760 1850 7800
rect 1890 7760 1910 7800
rect 1830 7700 1910 7760
rect 1830 7660 1850 7700
rect 1890 7660 1910 7700
rect 1830 7630 1910 7660
rect 1950 7800 2030 7830
rect 1950 7760 1970 7800
rect 2010 7760 2030 7800
rect 1950 7700 2030 7760
rect 1950 7660 1970 7700
rect 2010 7660 2030 7700
rect 1950 7630 2030 7660
rect 2070 7800 2150 7830
rect 2070 7760 2090 7800
rect 2130 7760 2150 7800
rect 2070 7700 2150 7760
rect 2070 7660 2090 7700
rect 2130 7660 2150 7700
rect 2070 7630 2150 7660
rect 2190 7800 2270 7830
rect 2190 7760 2210 7800
rect 2250 7760 2270 7800
rect 2190 7700 2270 7760
rect 2190 7660 2210 7700
rect 2250 7660 2270 7700
rect 2190 7630 2270 7660
rect 2310 7800 2390 7830
rect 2310 7760 2330 7800
rect 2370 7760 2390 7800
rect 2310 7700 2390 7760
rect 2310 7660 2330 7700
rect 2370 7660 2390 7700
rect 2310 7630 2390 7660
rect 2430 7800 2510 7830
rect 2430 7760 2450 7800
rect 2490 7760 2510 7800
rect 2430 7700 2510 7760
rect 2430 7660 2450 7700
rect 2490 7660 2510 7700
rect 2430 7630 2510 7660
rect 2550 7800 2630 7830
rect 2550 7760 2570 7800
rect 2610 7760 2630 7800
rect 2550 7700 2630 7760
rect 2550 7660 2570 7700
rect 2610 7660 2630 7700
rect 2550 7630 2630 7660
rect 2670 7800 2750 7830
rect 2670 7760 2690 7800
rect 2730 7760 2750 7800
rect 2670 7700 2750 7760
rect 2670 7660 2690 7700
rect 2730 7660 2750 7700
rect 2670 7630 2750 7660
rect 2790 7800 2870 7830
rect 2790 7760 2810 7800
rect 2850 7760 2870 7800
rect 2790 7700 2870 7760
rect 2790 7660 2810 7700
rect 2850 7660 2870 7700
rect 2790 7630 2870 7660
rect 2910 7800 2990 7830
rect 2910 7760 2930 7800
rect 2970 7760 2990 7800
rect 2910 7700 2990 7760
rect 2910 7660 2930 7700
rect 2970 7660 2990 7700
rect 2910 7630 2990 7660
rect 3550 7800 3630 7830
rect 3550 7760 3570 7800
rect 3610 7760 3630 7800
rect 3550 7700 3630 7760
rect 3550 7660 3570 7700
rect 3610 7660 3630 7700
rect 3550 7630 3630 7660
rect 3670 7800 3750 7830
rect 3670 7760 3690 7800
rect 3730 7760 3750 7800
rect 3670 7700 3750 7760
rect 3670 7660 3690 7700
rect 3730 7660 3750 7700
rect 3670 7630 3750 7660
rect 3790 7800 3870 7830
rect 3790 7760 3810 7800
rect 3850 7760 3870 7800
rect 3790 7700 3870 7760
rect 3790 7660 3810 7700
rect 3850 7660 3870 7700
rect 3790 7630 3870 7660
rect 3910 7800 3990 7830
rect 3910 7760 3930 7800
rect 3970 7760 3990 7800
rect 3910 7700 3990 7760
rect 3910 7660 3930 7700
rect 3970 7660 3990 7700
rect 3910 7630 3990 7660
rect 4030 7800 4110 7830
rect 4030 7760 4050 7800
rect 4090 7760 4110 7800
rect 4030 7700 4110 7760
rect 4030 7660 4050 7700
rect 4090 7660 4110 7700
rect 4030 7630 4110 7660
rect 4150 7800 4230 7830
rect 4150 7760 4170 7800
rect 4210 7760 4230 7800
rect 4150 7700 4230 7760
rect 4150 7660 4170 7700
rect 4210 7660 4230 7700
rect 4150 7630 4230 7660
rect 4270 7800 4350 7830
rect 4270 7760 4290 7800
rect 4330 7760 4350 7800
rect 4270 7700 4350 7760
rect 4270 7660 4290 7700
rect 4330 7660 4350 7700
rect 4270 7630 4350 7660
rect 4390 7800 4470 7830
rect 4390 7760 4410 7800
rect 4450 7760 4470 7800
rect 4390 7700 4470 7760
rect 4390 7660 4410 7700
rect 4450 7660 4470 7700
rect 4390 7630 4470 7660
rect 4510 7800 4590 7830
rect 4510 7760 4530 7800
rect 4570 7760 4590 7800
rect 4510 7700 4590 7760
rect 4510 7660 4530 7700
rect 4570 7660 4590 7700
rect 4510 7630 4590 7660
rect 4630 7800 4710 7830
rect 4630 7760 4650 7800
rect 4690 7760 4710 7800
rect 4630 7700 4710 7760
rect 4630 7660 4650 7700
rect 4690 7660 4710 7700
rect 4630 7630 4710 7660
rect 4750 7800 4830 7830
rect 4750 7760 4770 7800
rect 4810 7760 4830 7800
rect 4750 7700 4830 7760
rect 4750 7660 4770 7700
rect 4810 7660 4830 7700
rect 4750 7630 4830 7660
rect 4870 7800 4950 7830
rect 4870 7760 4890 7800
rect 4930 7760 4950 7800
rect 4870 7700 4950 7760
rect 4870 7660 4890 7700
rect 4930 7660 4950 7700
rect 4870 7630 4950 7660
rect 4990 7800 5070 7830
rect 4990 7760 5010 7800
rect 5050 7760 5070 7800
rect 4990 7700 5070 7760
rect 4990 7660 5010 7700
rect 5050 7660 5070 7700
rect 4990 7630 5070 7660
rect 5110 7800 5190 7830
rect 5110 7760 5130 7800
rect 5170 7760 5190 7800
rect 5110 7700 5190 7760
rect 5110 7660 5130 7700
rect 5170 7660 5190 7700
rect 5110 7630 5190 7660
rect 5230 7800 5310 7830
rect 5230 7760 5250 7800
rect 5290 7760 5310 7800
rect 5230 7700 5310 7760
rect 5230 7660 5250 7700
rect 5290 7660 5310 7700
rect 5230 7630 5310 7660
rect 5350 7800 5430 7830
rect 5350 7760 5370 7800
rect 5410 7760 5430 7800
rect 5350 7700 5430 7760
rect 5350 7660 5370 7700
rect 5410 7660 5430 7700
rect 5350 7630 5430 7660
rect 5470 7800 5550 7830
rect 5470 7760 5490 7800
rect 5530 7760 5550 7800
rect 5470 7700 5550 7760
rect 5470 7660 5490 7700
rect 5530 7660 5550 7700
rect 5470 7630 5550 7660
rect 5590 7800 5670 7830
rect 5590 7760 5610 7800
rect 5650 7760 5670 7800
rect 5590 7700 5670 7760
rect 5590 7660 5610 7700
rect 5650 7660 5670 7700
rect 5590 7630 5670 7660
rect 5710 7800 5790 7830
rect 5710 7760 5730 7800
rect 5770 7760 5790 7800
rect 5710 7700 5790 7760
rect 5710 7660 5730 7700
rect 5770 7660 5790 7700
rect 5710 7630 5790 7660
rect 5830 7800 5910 7830
rect 5830 7760 5850 7800
rect 5890 7760 5910 7800
rect 5830 7700 5910 7760
rect 5830 7660 5850 7700
rect 5890 7660 5910 7700
rect 5830 7630 5910 7660
rect 5950 7800 6030 7830
rect 5950 7760 5970 7800
rect 6010 7760 6030 7800
rect 5950 7700 6030 7760
rect 5950 7660 5970 7700
rect 6010 7660 6030 7700
rect 5950 7630 6030 7660
rect 8250 7320 8350 7350
rect 8250 7280 8280 7320
rect 8320 7280 8350 7320
rect 8250 7220 8350 7280
rect 8250 7180 8280 7220
rect 8320 7180 8350 7220
rect 8250 7150 8350 7180
rect 8380 7320 8480 7350
rect 8380 7280 8410 7320
rect 8450 7280 8480 7320
rect 8380 7220 8480 7280
rect 8380 7180 8410 7220
rect 8450 7180 8480 7220
rect 8380 7150 8480 7180
rect 8510 7320 8610 7350
rect 8510 7280 8540 7320
rect 8580 7280 8610 7320
rect 8510 7220 8610 7280
rect 8510 7180 8540 7220
rect 8580 7180 8610 7220
rect 8510 7150 8610 7180
rect 8640 7320 8740 7350
rect 8640 7280 8670 7320
rect 8710 7280 8740 7320
rect 8640 7220 8740 7280
rect 8640 7180 8670 7220
rect 8710 7180 8740 7220
rect 8640 7150 8740 7180
rect 8770 7320 8870 7350
rect 8770 7280 8800 7320
rect 8840 7280 8870 7320
rect 8770 7220 8870 7280
rect 8770 7180 8800 7220
rect 8840 7180 8870 7220
rect 8770 7150 8870 7180
rect 8900 7320 9000 7350
rect 8900 7280 8930 7320
rect 8970 7280 9000 7320
rect 8900 7220 9000 7280
rect 8900 7180 8930 7220
rect 8970 7180 9000 7220
rect 8900 7150 9000 7180
rect 9030 7320 9130 7350
rect 9030 7280 9060 7320
rect 9100 7280 9130 7320
rect 9030 7220 9130 7280
rect 9030 7180 9060 7220
rect 9100 7180 9130 7220
rect 9030 7150 9130 7180
rect 9390 7320 9490 7350
rect 9390 7280 9420 7320
rect 9460 7280 9490 7320
rect 9390 7220 9490 7280
rect 9390 7180 9420 7220
rect 9460 7180 9490 7220
rect 9390 7150 9490 7180
rect 9520 7320 9620 7350
rect 9520 7280 9550 7320
rect 9590 7280 9620 7320
rect 9520 7220 9620 7280
rect 9520 7180 9550 7220
rect 9590 7180 9620 7220
rect 9520 7150 9620 7180
rect 9650 7320 9750 7350
rect 9650 7280 9680 7320
rect 9720 7280 9750 7320
rect 9650 7220 9750 7280
rect 9650 7180 9680 7220
rect 9720 7180 9750 7220
rect 9650 7150 9750 7180
rect 9780 7320 9880 7350
rect 9780 7280 9810 7320
rect 9850 7280 9880 7320
rect 9780 7220 9880 7280
rect 9780 7180 9810 7220
rect 9850 7180 9880 7220
rect 9780 7150 9880 7180
rect 9910 7320 10010 7350
rect 9910 7280 9940 7320
rect 9980 7280 10010 7320
rect 9910 7220 10010 7280
rect 9910 7180 9940 7220
rect 9980 7180 10010 7220
rect 9910 7150 10010 7180
rect 10040 7320 10140 7350
rect 10040 7280 10070 7320
rect 10110 7280 10140 7320
rect 10040 7220 10140 7280
rect 10040 7180 10070 7220
rect 10110 7180 10140 7220
rect 10040 7150 10140 7180
rect 10170 7320 10270 7350
rect 10170 7280 10200 7320
rect 10240 7280 10270 7320
rect 10170 7220 10270 7280
rect 10170 7180 10200 7220
rect 10240 7180 10270 7220
rect 10170 7150 10270 7180
rect 10530 7320 10630 7350
rect 10530 7280 10560 7320
rect 10600 7280 10630 7320
rect 10530 7220 10630 7280
rect 10530 7180 10560 7220
rect 10600 7180 10630 7220
rect 10530 7150 10630 7180
rect 10660 7320 10760 7350
rect 10660 7280 10690 7320
rect 10730 7280 10760 7320
rect 10660 7220 10760 7280
rect 10660 7180 10690 7220
rect 10730 7180 10760 7220
rect 10660 7150 10760 7180
rect 10790 7320 10890 7350
rect 10790 7280 10820 7320
rect 10860 7280 10890 7320
rect 10790 7220 10890 7280
rect 10790 7180 10820 7220
rect 10860 7180 10890 7220
rect 10790 7150 10890 7180
rect 10920 7320 11020 7350
rect 10920 7280 10950 7320
rect 10990 7280 11020 7320
rect 10920 7220 11020 7280
rect 10920 7180 10950 7220
rect 10990 7180 11020 7220
rect 10920 7150 11020 7180
rect 11050 7320 11150 7350
rect 11050 7280 11080 7320
rect 11120 7280 11150 7320
rect 11050 7220 11150 7280
rect 11050 7180 11080 7220
rect 11120 7180 11150 7220
rect 11050 7150 11150 7180
rect 11180 7320 11280 7350
rect 11180 7280 11210 7320
rect 11250 7280 11280 7320
rect 11180 7220 11280 7280
rect 11180 7180 11210 7220
rect 11250 7180 11280 7220
rect 11180 7150 11280 7180
rect 11310 7320 11410 7350
rect 11310 7280 11340 7320
rect 11380 7280 11410 7320
rect 11310 7220 11410 7280
rect 11310 7180 11340 7220
rect 11380 7180 11410 7220
rect 11310 7150 11410 7180
rect 8320 6670 8420 6700
rect 1610 6640 1690 6670
rect 1610 6600 1630 6640
rect 1670 6600 1690 6640
rect 1610 6540 1690 6600
rect 1610 6500 1630 6540
rect 1670 6500 1690 6540
rect 1610 6440 1690 6500
rect 1610 6400 1630 6440
rect 1670 6400 1690 6440
rect 1610 6340 1690 6400
rect 1610 6300 1630 6340
rect 1670 6300 1690 6340
rect 1610 6240 1690 6300
rect 1610 6200 1630 6240
rect 1670 6200 1690 6240
rect 1610 6140 1690 6200
rect 1610 6100 1630 6140
rect 1670 6100 1690 6140
rect 1610 6070 1690 6100
rect 1790 6640 1870 6670
rect 1790 6600 1810 6640
rect 1850 6600 1870 6640
rect 1790 6540 1870 6600
rect 1790 6500 1810 6540
rect 1850 6500 1870 6540
rect 1790 6440 1870 6500
rect 1790 6400 1810 6440
rect 1850 6400 1870 6440
rect 1790 6340 1870 6400
rect 1790 6300 1810 6340
rect 1850 6300 1870 6340
rect 1790 6240 1870 6300
rect 1790 6200 1810 6240
rect 1850 6200 1870 6240
rect 1790 6140 1870 6200
rect 1790 6100 1810 6140
rect 1850 6100 1870 6140
rect 1790 6070 1870 6100
rect 1970 6640 2050 6670
rect 1970 6600 1990 6640
rect 2030 6600 2050 6640
rect 1970 6540 2050 6600
rect 1970 6500 1990 6540
rect 2030 6500 2050 6540
rect 1970 6440 2050 6500
rect 1970 6400 1990 6440
rect 2030 6400 2050 6440
rect 1970 6340 2050 6400
rect 1970 6300 1990 6340
rect 2030 6300 2050 6340
rect 1970 6240 2050 6300
rect 1970 6200 1990 6240
rect 2030 6200 2050 6240
rect 1970 6140 2050 6200
rect 1970 6100 1990 6140
rect 2030 6100 2050 6140
rect 1970 6070 2050 6100
rect 2150 6640 2230 6670
rect 2150 6600 2170 6640
rect 2210 6600 2230 6640
rect 2150 6540 2230 6600
rect 2150 6500 2170 6540
rect 2210 6500 2230 6540
rect 2150 6440 2230 6500
rect 2150 6400 2170 6440
rect 2210 6400 2230 6440
rect 2150 6340 2230 6400
rect 2150 6300 2170 6340
rect 2210 6300 2230 6340
rect 2150 6240 2230 6300
rect 2150 6200 2170 6240
rect 2210 6200 2230 6240
rect 2150 6140 2230 6200
rect 2150 6100 2170 6140
rect 2210 6100 2230 6140
rect 2150 6070 2230 6100
rect 2330 6640 2410 6670
rect 2330 6600 2350 6640
rect 2390 6600 2410 6640
rect 2330 6540 2410 6600
rect 2330 6500 2350 6540
rect 2390 6500 2410 6540
rect 2330 6440 2410 6500
rect 2330 6400 2350 6440
rect 2390 6400 2410 6440
rect 2330 6340 2410 6400
rect 2330 6300 2350 6340
rect 2390 6300 2410 6340
rect 2330 6240 2410 6300
rect 2330 6200 2350 6240
rect 2390 6200 2410 6240
rect 2330 6140 2410 6200
rect 2330 6100 2350 6140
rect 2390 6100 2410 6140
rect 2330 6070 2410 6100
rect 2510 6640 2590 6670
rect 2510 6600 2530 6640
rect 2570 6600 2590 6640
rect 2510 6540 2590 6600
rect 2510 6500 2530 6540
rect 2570 6500 2590 6540
rect 2510 6440 2590 6500
rect 2510 6400 2530 6440
rect 2570 6400 2590 6440
rect 2510 6340 2590 6400
rect 2510 6300 2530 6340
rect 2570 6300 2590 6340
rect 2510 6240 2590 6300
rect 2510 6200 2530 6240
rect 2570 6200 2590 6240
rect 2510 6140 2590 6200
rect 2510 6100 2530 6140
rect 2570 6100 2590 6140
rect 2510 6070 2590 6100
rect 2690 6640 2770 6670
rect 2690 6600 2710 6640
rect 2750 6600 2770 6640
rect 2690 6540 2770 6600
rect 2690 6500 2710 6540
rect 2750 6500 2770 6540
rect 2690 6440 2770 6500
rect 2690 6400 2710 6440
rect 2750 6400 2770 6440
rect 2690 6340 2770 6400
rect 2690 6300 2710 6340
rect 2750 6300 2770 6340
rect 2690 6240 2770 6300
rect 2690 6200 2710 6240
rect 2750 6200 2770 6240
rect 2690 6140 2770 6200
rect 2690 6100 2710 6140
rect 2750 6100 2770 6140
rect 2690 6070 2770 6100
rect 2870 6640 2950 6670
rect 2870 6600 2890 6640
rect 2930 6600 2950 6640
rect 2870 6540 2950 6600
rect 2870 6500 2890 6540
rect 2930 6500 2950 6540
rect 2870 6440 2950 6500
rect 2870 6400 2890 6440
rect 2930 6400 2950 6440
rect 2870 6340 2950 6400
rect 2870 6300 2890 6340
rect 2930 6300 2950 6340
rect 2870 6240 2950 6300
rect 2870 6200 2890 6240
rect 2930 6200 2950 6240
rect 2870 6140 2950 6200
rect 2870 6100 2890 6140
rect 2930 6100 2950 6140
rect 2870 6070 2950 6100
rect 3050 6640 3130 6670
rect 3050 6600 3070 6640
rect 3110 6600 3130 6640
rect 3050 6540 3130 6600
rect 3050 6500 3070 6540
rect 3110 6500 3130 6540
rect 3050 6440 3130 6500
rect 3050 6400 3070 6440
rect 3110 6400 3130 6440
rect 3050 6340 3130 6400
rect 3050 6300 3070 6340
rect 3110 6300 3130 6340
rect 3050 6240 3130 6300
rect 3050 6200 3070 6240
rect 3110 6200 3130 6240
rect 3050 6140 3130 6200
rect 3050 6100 3070 6140
rect 3110 6100 3130 6140
rect 3050 6070 3130 6100
rect 3230 6640 3310 6670
rect 3230 6600 3250 6640
rect 3290 6600 3310 6640
rect 3230 6540 3310 6600
rect 3230 6500 3250 6540
rect 3290 6500 3310 6540
rect 3230 6440 3310 6500
rect 3230 6400 3250 6440
rect 3290 6400 3310 6440
rect 3230 6340 3310 6400
rect 3230 6300 3250 6340
rect 3290 6300 3310 6340
rect 3230 6240 3310 6300
rect 3230 6200 3250 6240
rect 3290 6200 3310 6240
rect 3230 6140 3310 6200
rect 3230 6100 3250 6140
rect 3290 6100 3310 6140
rect 3230 6070 3310 6100
rect 3410 6640 3490 6670
rect 3410 6600 3430 6640
rect 3470 6600 3490 6640
rect 3410 6540 3490 6600
rect 3410 6500 3430 6540
rect 3470 6500 3490 6540
rect 3410 6440 3490 6500
rect 3410 6400 3430 6440
rect 3470 6400 3490 6440
rect 3410 6340 3490 6400
rect 3410 6300 3430 6340
rect 3470 6300 3490 6340
rect 3410 6240 3490 6300
rect 3410 6200 3430 6240
rect 3470 6200 3490 6240
rect 3410 6140 3490 6200
rect 3410 6100 3430 6140
rect 3470 6100 3490 6140
rect 3410 6070 3490 6100
rect 3590 6640 3670 6670
rect 3590 6600 3610 6640
rect 3650 6600 3670 6640
rect 3590 6540 3670 6600
rect 3590 6500 3610 6540
rect 3650 6500 3670 6540
rect 3590 6440 3670 6500
rect 3590 6400 3610 6440
rect 3650 6400 3670 6440
rect 3590 6340 3670 6400
rect 3590 6300 3610 6340
rect 3650 6300 3670 6340
rect 3590 6240 3670 6300
rect 3590 6200 3610 6240
rect 3650 6200 3670 6240
rect 3590 6140 3670 6200
rect 3590 6100 3610 6140
rect 3650 6100 3670 6140
rect 3590 6070 3670 6100
rect 3770 6640 3850 6670
rect 3770 6600 3790 6640
rect 3830 6600 3850 6640
rect 3770 6540 3850 6600
rect 3770 6500 3790 6540
rect 3830 6500 3850 6540
rect 3770 6440 3850 6500
rect 3770 6400 3790 6440
rect 3830 6400 3850 6440
rect 3770 6340 3850 6400
rect 3770 6300 3790 6340
rect 3830 6300 3850 6340
rect 3770 6240 3850 6300
rect 3770 6200 3790 6240
rect 3830 6200 3850 6240
rect 3770 6140 3850 6200
rect 3770 6100 3790 6140
rect 3830 6100 3850 6140
rect 3770 6070 3850 6100
rect 3950 6640 4030 6670
rect 3950 6600 3970 6640
rect 4010 6600 4030 6640
rect 3950 6540 4030 6600
rect 3950 6500 3970 6540
rect 4010 6500 4030 6540
rect 3950 6440 4030 6500
rect 3950 6400 3970 6440
rect 4010 6400 4030 6440
rect 3950 6340 4030 6400
rect 3950 6300 3970 6340
rect 4010 6300 4030 6340
rect 3950 6240 4030 6300
rect 3950 6200 3970 6240
rect 4010 6200 4030 6240
rect 3950 6140 4030 6200
rect 3950 6100 3970 6140
rect 4010 6100 4030 6140
rect 3950 6070 4030 6100
rect 4130 6640 4210 6670
rect 4130 6600 4150 6640
rect 4190 6600 4210 6640
rect 4130 6540 4210 6600
rect 4130 6500 4150 6540
rect 4190 6500 4210 6540
rect 4130 6440 4210 6500
rect 4130 6400 4150 6440
rect 4190 6400 4210 6440
rect 4130 6340 4210 6400
rect 4130 6300 4150 6340
rect 4190 6300 4210 6340
rect 4130 6240 4210 6300
rect 4130 6200 4150 6240
rect 4190 6200 4210 6240
rect 4130 6140 4210 6200
rect 4130 6100 4150 6140
rect 4190 6100 4210 6140
rect 4130 6070 4210 6100
rect 4310 6640 4390 6670
rect 4310 6600 4330 6640
rect 4370 6600 4390 6640
rect 4310 6540 4390 6600
rect 4310 6500 4330 6540
rect 4370 6500 4390 6540
rect 4310 6440 4390 6500
rect 4310 6400 4330 6440
rect 4370 6400 4390 6440
rect 4310 6340 4390 6400
rect 4310 6300 4330 6340
rect 4370 6300 4390 6340
rect 4310 6240 4390 6300
rect 4310 6200 4330 6240
rect 4370 6200 4390 6240
rect 4310 6140 4390 6200
rect 4310 6100 4330 6140
rect 4370 6100 4390 6140
rect 4310 6070 4390 6100
rect 4490 6640 4570 6670
rect 4490 6600 4510 6640
rect 4550 6600 4570 6640
rect 4490 6540 4570 6600
rect 4490 6500 4510 6540
rect 4550 6500 4570 6540
rect 4490 6440 4570 6500
rect 4490 6400 4510 6440
rect 4550 6400 4570 6440
rect 4490 6340 4570 6400
rect 4490 6300 4510 6340
rect 4550 6300 4570 6340
rect 4490 6240 4570 6300
rect 4490 6200 4510 6240
rect 4550 6200 4570 6240
rect 4490 6140 4570 6200
rect 4490 6100 4510 6140
rect 4550 6100 4570 6140
rect 4490 6070 4570 6100
rect 4670 6640 4750 6670
rect 4670 6600 4690 6640
rect 4730 6600 4750 6640
rect 4670 6540 4750 6600
rect 4670 6500 4690 6540
rect 4730 6500 4750 6540
rect 4670 6440 4750 6500
rect 4670 6400 4690 6440
rect 4730 6400 4750 6440
rect 4670 6340 4750 6400
rect 4670 6300 4690 6340
rect 4730 6300 4750 6340
rect 4670 6240 4750 6300
rect 4670 6200 4690 6240
rect 4730 6200 4750 6240
rect 4670 6140 4750 6200
rect 4670 6100 4690 6140
rect 4730 6100 4750 6140
rect 4670 6070 4750 6100
rect 4850 6640 4930 6670
rect 4850 6600 4870 6640
rect 4910 6600 4930 6640
rect 4850 6540 4930 6600
rect 8320 6630 8350 6670
rect 8390 6630 8420 6670
rect 4850 6500 4870 6540
rect 4910 6500 4930 6540
rect 8320 6570 8420 6630
rect 8320 6530 8350 6570
rect 8390 6530 8420 6570
rect 4850 6440 4930 6500
rect 8320 6470 8420 6530
rect 4850 6400 4870 6440
rect 4910 6400 4930 6440
rect 4850 6340 4930 6400
rect 4850 6300 4870 6340
rect 4910 6300 4930 6340
rect 4850 6240 4930 6300
rect 5470 6440 5560 6470
rect 5470 6400 5500 6440
rect 5540 6400 5560 6440
rect 5470 6340 5560 6400
rect 5470 6300 5500 6340
rect 5540 6300 5560 6340
rect 5470 6270 5560 6300
rect 5590 6440 5670 6470
rect 5590 6400 5610 6440
rect 5650 6400 5670 6440
rect 5590 6340 5670 6400
rect 5590 6300 5610 6340
rect 5650 6300 5670 6340
rect 5590 6270 5670 6300
rect 5700 6440 5780 6470
rect 5700 6400 5720 6440
rect 5760 6400 5780 6440
rect 5700 6340 5780 6400
rect 5700 6300 5720 6340
rect 5760 6300 5780 6340
rect 5700 6270 5780 6300
rect 5810 6440 5890 6470
rect 5810 6400 5830 6440
rect 5870 6400 5890 6440
rect 5810 6340 5890 6400
rect 5810 6300 5830 6340
rect 5870 6300 5890 6340
rect 5810 6270 5890 6300
rect 5920 6440 6000 6470
rect 5920 6400 5940 6440
rect 5980 6400 6000 6440
rect 5920 6340 6000 6400
rect 5920 6300 5940 6340
rect 5980 6300 6000 6340
rect 5920 6270 6000 6300
rect 8320 6430 8350 6470
rect 8390 6430 8420 6470
rect 8320 6370 8420 6430
rect 8320 6330 8350 6370
rect 8390 6330 8420 6370
rect 8320 6270 8420 6330
rect 4850 6200 4870 6240
rect 4910 6200 4930 6240
rect 4850 6140 4930 6200
rect 8320 6230 8350 6270
rect 8390 6230 8420 6270
rect 8320 6200 8420 6230
rect 8520 6670 8620 6700
rect 8520 6630 8550 6670
rect 8590 6630 8620 6670
rect 8520 6570 8620 6630
rect 8520 6530 8550 6570
rect 8590 6530 8620 6570
rect 8520 6470 8620 6530
rect 8520 6430 8550 6470
rect 8590 6430 8620 6470
rect 8520 6370 8620 6430
rect 8520 6330 8550 6370
rect 8590 6330 8620 6370
rect 8520 6270 8620 6330
rect 8520 6230 8550 6270
rect 8590 6230 8620 6270
rect 8520 6200 8620 6230
rect 8720 6670 8820 6700
rect 8720 6630 8750 6670
rect 8790 6630 8820 6670
rect 8720 6570 8820 6630
rect 8720 6530 8750 6570
rect 8790 6530 8820 6570
rect 8720 6470 8820 6530
rect 8720 6430 8750 6470
rect 8790 6430 8820 6470
rect 8720 6370 8820 6430
rect 8720 6330 8750 6370
rect 8790 6330 8820 6370
rect 8720 6270 8820 6330
rect 8720 6230 8750 6270
rect 8790 6230 8820 6270
rect 8720 6200 8820 6230
rect 8920 6670 9020 6700
rect 8920 6630 8950 6670
rect 8990 6630 9020 6670
rect 8920 6570 9020 6630
rect 8920 6530 8950 6570
rect 8990 6530 9020 6570
rect 8920 6470 9020 6530
rect 8920 6430 8950 6470
rect 8990 6430 9020 6470
rect 8920 6370 9020 6430
rect 8920 6330 8950 6370
rect 8990 6330 9020 6370
rect 8920 6270 9020 6330
rect 8920 6230 8950 6270
rect 8990 6230 9020 6270
rect 8920 6200 9020 6230
rect 9120 6670 9220 6700
rect 9120 6630 9150 6670
rect 9190 6630 9220 6670
rect 9120 6570 9220 6630
rect 9120 6530 9150 6570
rect 9190 6530 9220 6570
rect 9120 6470 9220 6530
rect 9120 6430 9150 6470
rect 9190 6430 9220 6470
rect 9120 6370 9220 6430
rect 9120 6330 9150 6370
rect 9190 6330 9220 6370
rect 9120 6270 9220 6330
rect 9120 6230 9150 6270
rect 9190 6230 9220 6270
rect 9120 6200 9220 6230
rect 9320 6670 9420 6700
rect 9320 6630 9350 6670
rect 9390 6630 9420 6670
rect 9320 6570 9420 6630
rect 9320 6530 9350 6570
rect 9390 6530 9420 6570
rect 9320 6470 9420 6530
rect 9320 6430 9350 6470
rect 9390 6430 9420 6470
rect 9320 6370 9420 6430
rect 9320 6330 9350 6370
rect 9390 6330 9420 6370
rect 9320 6270 9420 6330
rect 9320 6230 9350 6270
rect 9390 6230 9420 6270
rect 9320 6200 9420 6230
rect 9520 6670 9620 6700
rect 9520 6630 9550 6670
rect 9590 6630 9620 6670
rect 9520 6570 9620 6630
rect 9520 6530 9550 6570
rect 9590 6530 9620 6570
rect 9520 6470 9620 6530
rect 9520 6430 9550 6470
rect 9590 6430 9620 6470
rect 9520 6370 9620 6430
rect 9520 6330 9550 6370
rect 9590 6330 9620 6370
rect 9520 6270 9620 6330
rect 9520 6230 9550 6270
rect 9590 6230 9620 6270
rect 9520 6200 9620 6230
rect 9720 6670 9820 6700
rect 9720 6630 9750 6670
rect 9790 6630 9820 6670
rect 9720 6570 9820 6630
rect 9720 6530 9750 6570
rect 9790 6530 9820 6570
rect 9720 6470 9820 6530
rect 9720 6430 9750 6470
rect 9790 6430 9820 6470
rect 9720 6370 9820 6430
rect 9720 6330 9750 6370
rect 9790 6330 9820 6370
rect 9720 6270 9820 6330
rect 9720 6230 9750 6270
rect 9790 6230 9820 6270
rect 9720 6200 9820 6230
rect 9920 6670 10020 6700
rect 9920 6630 9950 6670
rect 9990 6630 10020 6670
rect 9920 6570 10020 6630
rect 9920 6530 9950 6570
rect 9990 6530 10020 6570
rect 9920 6470 10020 6530
rect 9920 6430 9950 6470
rect 9990 6430 10020 6470
rect 9920 6370 10020 6430
rect 9920 6330 9950 6370
rect 9990 6330 10020 6370
rect 9920 6270 10020 6330
rect 9920 6230 9950 6270
rect 9990 6230 10020 6270
rect 9920 6200 10020 6230
rect 10120 6670 10220 6700
rect 10120 6630 10150 6670
rect 10190 6630 10220 6670
rect 10120 6570 10220 6630
rect 10120 6530 10150 6570
rect 10190 6530 10220 6570
rect 10120 6470 10220 6530
rect 10120 6430 10150 6470
rect 10190 6430 10220 6470
rect 10120 6370 10220 6430
rect 10120 6330 10150 6370
rect 10190 6330 10220 6370
rect 10120 6270 10220 6330
rect 10120 6230 10150 6270
rect 10190 6230 10220 6270
rect 10120 6200 10220 6230
rect 10320 6670 10420 6700
rect 10320 6630 10350 6670
rect 10390 6630 10420 6670
rect 10320 6570 10420 6630
rect 10320 6530 10350 6570
rect 10390 6530 10420 6570
rect 10320 6470 10420 6530
rect 10320 6430 10350 6470
rect 10390 6430 10420 6470
rect 10320 6370 10420 6430
rect 10320 6330 10350 6370
rect 10390 6330 10420 6370
rect 10320 6270 10420 6330
rect 10320 6230 10350 6270
rect 10390 6230 10420 6270
rect 10320 6200 10420 6230
rect 4850 6100 4870 6140
rect 4910 6100 4930 6140
rect 4850 6070 4930 6100
rect 1620 5640 1700 5670
rect 1620 5600 1640 5640
rect 1680 5600 1700 5640
rect 1620 5540 1700 5600
rect 1620 5500 1640 5540
rect 1680 5500 1700 5540
rect 1620 5470 1700 5500
rect 1730 5640 1810 5670
rect 1730 5600 1750 5640
rect 1790 5600 1810 5640
rect 1730 5540 1810 5600
rect 1730 5500 1750 5540
rect 1790 5500 1810 5540
rect 1730 5470 1810 5500
rect 1840 5640 1920 5670
rect 1840 5600 1860 5640
rect 1900 5600 1920 5640
rect 1840 5540 1920 5600
rect 1840 5500 1860 5540
rect 1900 5500 1920 5540
rect 1840 5470 1920 5500
rect 1950 5640 2030 5670
rect 1950 5600 1970 5640
rect 2010 5600 2030 5640
rect 1950 5540 2030 5600
rect 1950 5500 1970 5540
rect 2010 5500 2030 5540
rect 1950 5470 2030 5500
rect 2060 5640 2140 5670
rect 2060 5600 2080 5640
rect 2120 5600 2140 5640
rect 2060 5540 2140 5600
rect 2060 5500 2080 5540
rect 2120 5500 2140 5540
rect 2060 5470 2140 5500
rect 2170 5640 2250 5670
rect 2170 5600 2190 5640
rect 2230 5600 2250 5640
rect 2170 5540 2250 5600
rect 2170 5500 2190 5540
rect 2230 5500 2250 5540
rect 2170 5470 2250 5500
rect 2280 5640 2360 5670
rect 2280 5600 2300 5640
rect 2340 5600 2360 5640
rect 2280 5540 2360 5600
rect 2280 5500 2300 5540
rect 2340 5500 2360 5540
rect 2280 5470 2360 5500
rect 2390 5640 2470 5670
rect 2390 5600 2410 5640
rect 2450 5600 2470 5640
rect 2390 5540 2470 5600
rect 2390 5500 2410 5540
rect 2450 5500 2470 5540
rect 2390 5470 2470 5500
rect 2500 5640 2580 5670
rect 2500 5600 2520 5640
rect 2560 5600 2580 5640
rect 2500 5540 2580 5600
rect 2500 5500 2520 5540
rect 2560 5500 2580 5540
rect 2500 5470 2580 5500
rect 2610 5640 2690 5670
rect 2610 5600 2630 5640
rect 2670 5600 2690 5640
rect 2610 5540 2690 5600
rect 2610 5500 2630 5540
rect 2670 5500 2690 5540
rect 2610 5470 2690 5500
rect 2720 5640 2800 5670
rect 2720 5600 2740 5640
rect 2780 5600 2800 5640
rect 2720 5540 2800 5600
rect 2720 5500 2740 5540
rect 2780 5500 2800 5540
rect 2720 5470 2800 5500
rect 2830 5640 2910 5670
rect 2830 5600 2850 5640
rect 2890 5600 2910 5640
rect 2830 5540 2910 5600
rect 2830 5500 2850 5540
rect 2890 5500 2910 5540
rect 2830 5470 2910 5500
rect 2940 5640 3020 5670
rect 2940 5600 2960 5640
rect 3000 5600 3020 5640
rect 2940 5540 3020 5600
rect 2940 5500 2960 5540
rect 3000 5500 3020 5540
rect 2940 5470 3020 5500
rect 3520 5640 3600 5670
rect 3520 5600 3540 5640
rect 3580 5600 3600 5640
rect 3520 5540 3600 5600
rect 3520 5500 3540 5540
rect 3580 5500 3600 5540
rect 3520 5470 3600 5500
rect 3630 5640 3710 5670
rect 3630 5600 3650 5640
rect 3690 5600 3710 5640
rect 3630 5540 3710 5600
rect 3630 5500 3650 5540
rect 3690 5500 3710 5540
rect 3630 5470 3710 5500
rect 3740 5640 3820 5670
rect 3740 5600 3760 5640
rect 3800 5600 3820 5640
rect 3740 5540 3820 5600
rect 3740 5500 3760 5540
rect 3800 5500 3820 5540
rect 3740 5470 3820 5500
rect 3850 5640 3930 5670
rect 3850 5600 3870 5640
rect 3910 5600 3930 5640
rect 3850 5540 3930 5600
rect 3850 5500 3870 5540
rect 3910 5500 3930 5540
rect 3850 5470 3930 5500
rect 3960 5640 4040 5670
rect 3960 5600 3980 5640
rect 4020 5600 4040 5640
rect 3960 5540 4040 5600
rect 3960 5500 3980 5540
rect 4020 5500 4040 5540
rect 3960 5470 4040 5500
rect 4070 5640 4150 5670
rect 4070 5600 4090 5640
rect 4130 5600 4150 5640
rect 4070 5540 4150 5600
rect 4070 5500 4090 5540
rect 4130 5500 4150 5540
rect 4070 5470 4150 5500
rect 4180 5640 4260 5670
rect 4180 5600 4200 5640
rect 4240 5600 4260 5640
rect 4180 5540 4260 5600
rect 4180 5500 4200 5540
rect 4240 5500 4260 5540
rect 4180 5470 4260 5500
rect 4290 5640 4370 5670
rect 4290 5600 4310 5640
rect 4350 5600 4370 5640
rect 4290 5540 4370 5600
rect 4290 5500 4310 5540
rect 4350 5500 4370 5540
rect 4290 5470 4370 5500
rect 4400 5640 4480 5670
rect 4400 5600 4420 5640
rect 4460 5600 4480 5640
rect 4400 5540 4480 5600
rect 4400 5500 4420 5540
rect 4460 5500 4480 5540
rect 4400 5470 4480 5500
rect 4510 5640 4590 5670
rect 4510 5600 4530 5640
rect 4570 5600 4590 5640
rect 4510 5540 4590 5600
rect 4510 5500 4530 5540
rect 4570 5500 4590 5540
rect 4510 5470 4590 5500
rect 4620 5640 4700 5670
rect 4620 5600 4640 5640
rect 4680 5600 4700 5640
rect 4620 5540 4700 5600
rect 4620 5500 4640 5540
rect 4680 5500 4700 5540
rect 4620 5470 4700 5500
rect 4730 5640 4810 5670
rect 4730 5600 4750 5640
rect 4790 5600 4810 5640
rect 4730 5540 4810 5600
rect 4730 5500 4750 5540
rect 4790 5500 4810 5540
rect 4730 5470 4810 5500
rect 4840 5640 4920 5670
rect 4840 5600 4860 5640
rect 4900 5600 4920 5640
rect 4840 5540 4920 5600
rect 4840 5500 4860 5540
rect 4900 5500 4920 5540
rect 4840 5470 4920 5500
rect 2140 4280 2220 4310
rect 2140 4240 2160 4280
rect 2200 4240 2220 4280
rect 2140 4180 2220 4240
rect 2140 4140 2160 4180
rect 2200 4140 2220 4180
rect 2140 4080 2220 4140
rect 2140 4040 2160 4080
rect 2200 4040 2220 4080
rect 2140 3980 2220 4040
rect 2140 3940 2160 3980
rect 2200 3940 2220 3980
rect 2140 3910 2220 3940
rect 2250 4280 2330 4310
rect 2250 4240 2270 4280
rect 2310 4240 2330 4280
rect 2250 4180 2330 4240
rect 2250 4140 2270 4180
rect 2310 4140 2330 4180
rect 2250 4080 2330 4140
rect 2250 4040 2270 4080
rect 2310 4040 2330 4080
rect 2250 3980 2330 4040
rect 2250 3940 2270 3980
rect 2310 3940 2330 3980
rect 2250 3910 2330 3940
rect 2360 4280 2440 4310
rect 2360 4240 2380 4280
rect 2420 4240 2440 4280
rect 2360 4180 2440 4240
rect 2360 4140 2380 4180
rect 2420 4140 2440 4180
rect 2360 4080 2440 4140
rect 2360 4040 2380 4080
rect 2420 4040 2440 4080
rect 2360 3980 2440 4040
rect 2360 3940 2380 3980
rect 2420 3940 2440 3980
rect 2360 3910 2440 3940
rect 2660 4280 2740 4310
rect 2660 4240 2680 4280
rect 2720 4240 2740 4280
rect 2660 4180 2740 4240
rect 2660 4140 2680 4180
rect 2720 4140 2740 4180
rect 2660 4080 2740 4140
rect 2660 4040 2680 4080
rect 2720 4040 2740 4080
rect 2660 3980 2740 4040
rect 2660 3940 2680 3980
rect 2720 3940 2740 3980
rect 2660 3910 2740 3940
rect 2770 4280 2850 4310
rect 2770 4240 2790 4280
rect 2830 4240 2850 4280
rect 2770 4180 2850 4240
rect 2770 4140 2790 4180
rect 2830 4140 2850 4180
rect 2770 4080 2850 4140
rect 2770 4040 2790 4080
rect 2830 4040 2850 4080
rect 2770 3980 2850 4040
rect 2770 3940 2790 3980
rect 2830 3940 2850 3980
rect 2770 3910 2850 3940
rect 2880 4280 2960 4310
rect 3040 4280 3120 4310
rect 2880 4240 2900 4280
rect 2940 4240 2960 4280
rect 3040 4240 3060 4280
rect 3100 4240 3120 4280
rect 2880 4180 2960 4240
rect 3040 4180 3120 4240
rect 2880 4140 2900 4180
rect 2940 4140 2960 4180
rect 3040 4140 3060 4180
rect 3100 4140 3120 4180
rect 2880 4080 2960 4140
rect 3040 4080 3120 4140
rect 2880 4040 2900 4080
rect 2940 4040 2960 4080
rect 3040 4040 3060 4080
rect 3100 4040 3120 4080
rect 2880 3980 2960 4040
rect 3040 3980 3120 4040
rect 2880 3940 2900 3980
rect 2940 3940 2960 3980
rect 3040 3940 3060 3980
rect 3100 3940 3120 3980
rect 2880 3910 2960 3940
rect 3040 3910 3120 3940
rect 3150 4280 3230 4310
rect 3150 4240 3170 4280
rect 3210 4240 3230 4280
rect 3150 4180 3230 4240
rect 3150 4140 3170 4180
rect 3210 4140 3230 4180
rect 3150 4080 3230 4140
rect 3150 4040 3170 4080
rect 3210 4040 3230 4080
rect 3150 3980 3230 4040
rect 3150 3940 3170 3980
rect 3210 3940 3230 3980
rect 3150 3910 3230 3940
rect 3260 4280 3340 4310
rect 3260 4240 3280 4280
rect 3320 4240 3340 4280
rect 3260 4180 3340 4240
rect 3260 4140 3280 4180
rect 3320 4140 3340 4180
rect 3260 4080 3340 4140
rect 3260 4040 3280 4080
rect 3320 4040 3340 4080
rect 3260 3980 3340 4040
rect 8140 4330 8240 4360
rect 3260 3940 3280 3980
rect 3320 3940 3340 3980
rect 3260 3910 3340 3940
rect 3560 4280 3640 4310
rect 3560 4240 3580 4280
rect 3620 4240 3640 4280
rect 3560 4180 3640 4240
rect 3560 4140 3580 4180
rect 3620 4140 3640 4180
rect 3560 4080 3640 4140
rect 3560 4040 3580 4080
rect 3620 4040 3640 4080
rect 3560 3980 3640 4040
rect 3560 3940 3580 3980
rect 3620 3940 3640 3980
rect 3560 3910 3640 3940
rect 3670 4280 3750 4310
rect 3670 4240 3690 4280
rect 3730 4240 3750 4280
rect 3670 4180 3750 4240
rect 3670 4140 3690 4180
rect 3730 4140 3750 4180
rect 3670 4080 3750 4140
rect 3670 4040 3690 4080
rect 3730 4040 3750 4080
rect 3670 3980 3750 4040
rect 3670 3940 3690 3980
rect 3730 3940 3750 3980
rect 3670 3910 3750 3940
rect 3780 4280 3860 4310
rect 3780 4240 3800 4280
rect 3840 4240 3860 4280
rect 3780 4180 3860 4240
rect 3780 4140 3800 4180
rect 3840 4140 3860 4180
rect 3780 4080 3860 4140
rect 3780 4040 3800 4080
rect 3840 4040 3860 4080
rect 3780 3980 3860 4040
rect 3780 3940 3800 3980
rect 3840 3940 3860 3980
rect 3780 3910 3860 3940
rect 4080 4280 4160 4310
rect 4080 4240 4100 4280
rect 4140 4240 4160 4280
rect 4080 4180 4160 4240
rect 4080 4140 4100 4180
rect 4140 4140 4160 4180
rect 4080 4080 4160 4140
rect 4080 4040 4100 4080
rect 4140 4040 4160 4080
rect 4080 3980 4160 4040
rect 4080 3940 4100 3980
rect 4140 3940 4160 3980
rect 4080 3920 4160 3940
rect 4060 3910 4160 3920
rect 4190 4280 4270 4310
rect 4190 4240 4210 4280
rect 4250 4240 4270 4280
rect 4190 4180 4270 4240
rect 4190 4140 4210 4180
rect 4250 4140 4270 4180
rect 4190 4080 4270 4140
rect 4190 4040 4210 4080
rect 4250 4040 4270 4080
rect 4190 3980 4270 4040
rect 4190 3940 4210 3980
rect 4250 3940 4270 3980
rect 4190 3910 4270 3940
rect 4300 4280 4380 4310
rect 4300 4240 4320 4280
rect 4360 4240 4380 4280
rect 4300 4180 4380 4240
rect 4300 4140 4320 4180
rect 4360 4140 4380 4180
rect 4300 4080 4380 4140
rect 4300 4040 4320 4080
rect 4360 4040 4380 4080
rect 4300 3980 4380 4040
rect 4300 3940 4320 3980
rect 4360 3940 4380 3980
rect 4300 3910 4380 3940
rect 4520 4280 4600 4310
rect 4520 4240 4540 4280
rect 4580 4240 4600 4280
rect 4520 4180 4600 4240
rect 4520 4140 4540 4180
rect 4580 4140 4600 4180
rect 4520 4080 4600 4140
rect 4520 4040 4540 4080
rect 4580 4040 4600 4080
rect 4520 3980 4600 4040
rect 4520 3940 4540 3980
rect 4580 3940 4600 3980
rect 4520 3910 4600 3940
rect 4630 4280 4710 4310
rect 4630 4240 4650 4280
rect 4690 4240 4710 4280
rect 4630 4180 4710 4240
rect 4630 4140 4650 4180
rect 4690 4140 4710 4180
rect 4630 4080 4710 4140
rect 4630 4040 4650 4080
rect 4690 4040 4710 4080
rect 4630 3980 4710 4040
rect 4630 3940 4650 3980
rect 4690 3940 4710 3980
rect 4630 3910 4710 3940
rect 4850 4280 4930 4310
rect 4850 4240 4870 4280
rect 4910 4240 4930 4280
rect 4850 4180 4930 4240
rect 4850 4140 4870 4180
rect 4910 4140 4930 4180
rect 4850 4080 4930 4140
rect 4850 4040 4870 4080
rect 4910 4040 4930 4080
rect 4850 3980 4930 4040
rect 4850 3940 4870 3980
rect 4910 3940 4930 3980
rect 4850 3910 4930 3940
rect 4960 4280 5040 4310
rect 4960 4240 4980 4280
rect 5020 4240 5040 4280
rect 4960 4180 5040 4240
rect 4960 4140 4980 4180
rect 5020 4140 5040 4180
rect 4960 4080 5040 4140
rect 4960 4040 4980 4080
rect 5020 4040 5040 4080
rect 4960 3980 5040 4040
rect 4960 3940 4980 3980
rect 5020 3940 5040 3980
rect 4960 3910 5040 3940
rect 5270 4280 5370 4310
rect 5270 4240 5300 4280
rect 5340 4240 5370 4280
rect 5270 4180 5370 4240
rect 5270 4140 5300 4180
rect 5340 4140 5370 4180
rect 5270 4080 5370 4140
rect 5270 4040 5300 4080
rect 5340 4040 5370 4080
rect 5270 3980 5370 4040
rect 5270 3940 5300 3980
rect 5340 3940 5370 3980
rect 5270 3910 5370 3940
rect 5400 4280 5500 4310
rect 5400 4240 5430 4280
rect 5470 4240 5500 4280
rect 5400 4180 5500 4240
rect 5400 4140 5430 4180
rect 5470 4140 5500 4180
rect 5400 4080 5500 4140
rect 5400 4040 5430 4080
rect 5470 4040 5500 4080
rect 5400 3980 5500 4040
rect 5400 3940 5430 3980
rect 5470 3940 5500 3980
rect 5400 3910 5500 3940
rect 5660 4280 5760 4310
rect 5660 4240 5690 4280
rect 5730 4240 5760 4280
rect 5660 4180 5760 4240
rect 5660 4140 5690 4180
rect 5730 4140 5760 4180
rect 5660 4080 5760 4140
rect 5660 4040 5690 4080
rect 5730 4040 5760 4080
rect 5660 3980 5760 4040
rect 5660 3940 5690 3980
rect 5730 3940 5760 3980
rect 5660 3910 5760 3940
rect 5790 4280 5890 4310
rect 5790 4240 5820 4280
rect 5860 4240 5890 4280
rect 5790 4180 5890 4240
rect 5790 4140 5820 4180
rect 5860 4140 5890 4180
rect 5790 4080 5890 4140
rect 5790 4040 5820 4080
rect 5860 4040 5890 4080
rect 5790 3980 5890 4040
rect 5790 3940 5820 3980
rect 5860 3940 5890 3980
rect 5790 3910 5890 3940
rect 6050 4280 6150 4310
rect 6050 4240 6080 4280
rect 6120 4240 6150 4280
rect 6050 4180 6150 4240
rect 6050 4140 6080 4180
rect 6120 4140 6150 4180
rect 6050 4080 6150 4140
rect 6050 4040 6080 4080
rect 6120 4040 6150 4080
rect 6050 3980 6150 4040
rect 6050 3940 6080 3980
rect 6120 3940 6150 3980
rect 6050 3910 6150 3940
rect 6180 4280 6280 4310
rect 6180 4240 6210 4280
rect 6250 4240 6280 4280
rect 6180 4180 6280 4240
rect 6180 4140 6210 4180
rect 6250 4140 6280 4180
rect 6180 4080 6280 4140
rect 6180 4040 6210 4080
rect 6250 4040 6280 4080
rect 6180 3980 6280 4040
rect 6180 3940 6210 3980
rect 6250 3940 6280 3980
rect 6180 3910 6280 3940
rect 6340 4280 6440 4310
rect 6340 4240 6370 4280
rect 6410 4240 6440 4280
rect 6340 4180 6440 4240
rect 6340 4140 6370 4180
rect 6410 4140 6440 4180
rect 6340 4080 6440 4140
rect 6340 4040 6370 4080
rect 6410 4040 6440 4080
rect 6340 3980 6440 4040
rect 6340 3940 6370 3980
rect 6410 3940 6440 3980
rect 6340 3910 6440 3940
rect 6470 4280 6570 4310
rect 6470 4240 6500 4280
rect 6540 4240 6570 4280
rect 6470 4180 6570 4240
rect 6470 4140 6500 4180
rect 6540 4140 6570 4180
rect 6470 4080 6570 4140
rect 6470 4040 6500 4080
rect 6540 4040 6570 4080
rect 6470 3980 6570 4040
rect 6470 3940 6500 3980
rect 6540 3940 6570 3980
rect 6470 3910 6570 3940
rect 6730 4280 6830 4310
rect 6730 4240 6760 4280
rect 6800 4240 6830 4280
rect 6730 4180 6830 4240
rect 6730 4140 6760 4180
rect 6800 4140 6830 4180
rect 6730 4080 6830 4140
rect 6730 4040 6760 4080
rect 6800 4040 6830 4080
rect 6730 3980 6830 4040
rect 6730 3940 6760 3980
rect 6800 3940 6830 3980
rect 6730 3910 6830 3940
rect 6860 4280 6960 4310
rect 6860 4240 6890 4280
rect 6930 4240 6960 4280
rect 6860 4180 6960 4240
rect 6860 4140 6890 4180
rect 6930 4140 6960 4180
rect 6860 4080 6960 4140
rect 6860 4040 6890 4080
rect 6930 4040 6960 4080
rect 6860 3980 6960 4040
rect 6860 3940 6890 3980
rect 6930 3940 6960 3980
rect 8140 4290 8170 4330
rect 8210 4290 8240 4330
rect 8140 4230 8240 4290
rect 8140 4190 8170 4230
rect 8210 4190 8240 4230
rect 8140 4130 8240 4190
rect 8140 4090 8170 4130
rect 8210 4090 8240 4130
rect 8140 4030 8240 4090
rect 8140 3990 8170 4030
rect 8210 3990 8240 4030
rect 8140 3960 8240 3990
rect 8360 4330 8460 4360
rect 8360 4290 8390 4330
rect 8430 4290 8460 4330
rect 8360 4230 8460 4290
rect 8360 4190 8390 4230
rect 8430 4190 8460 4230
rect 8360 4130 8460 4190
rect 8360 4090 8390 4130
rect 8430 4090 8460 4130
rect 8360 4030 8460 4090
rect 8360 3990 8390 4030
rect 8430 3990 8460 4030
rect 8360 3960 8460 3990
rect 8580 4330 8680 4360
rect 8580 4290 8610 4330
rect 8650 4290 8680 4330
rect 8580 4230 8680 4290
rect 8580 4190 8610 4230
rect 8650 4190 8680 4230
rect 8580 4130 8680 4190
rect 8580 4090 8610 4130
rect 8650 4090 8680 4130
rect 8580 4030 8680 4090
rect 8580 3990 8610 4030
rect 8650 3990 8680 4030
rect 8580 3960 8680 3990
rect 8800 4330 8900 4360
rect 8800 4290 8830 4330
rect 8870 4290 8900 4330
rect 8800 4230 8900 4290
rect 8800 4190 8830 4230
rect 8870 4190 8900 4230
rect 8800 4130 8900 4190
rect 8800 4090 8830 4130
rect 8870 4090 8900 4130
rect 8800 4030 8900 4090
rect 8800 3990 8830 4030
rect 8870 3990 8900 4030
rect 8800 3960 8900 3990
rect 9020 4330 9120 4360
rect 9020 4290 9050 4330
rect 9090 4290 9120 4330
rect 9020 4230 9120 4290
rect 9020 4190 9050 4230
rect 9090 4190 9120 4230
rect 9020 4130 9120 4190
rect 9020 4090 9050 4130
rect 9090 4090 9120 4130
rect 9020 4030 9120 4090
rect 9020 3990 9050 4030
rect 9090 3990 9120 4030
rect 9020 3960 9120 3990
rect 9240 4330 9340 4360
rect 9240 4290 9270 4330
rect 9310 4290 9340 4330
rect 9240 4230 9340 4290
rect 9240 4190 9270 4230
rect 9310 4190 9340 4230
rect 9240 4130 9340 4190
rect 9240 4090 9270 4130
rect 9310 4090 9340 4130
rect 9240 4030 9340 4090
rect 9240 3990 9270 4030
rect 9310 3990 9340 4030
rect 9240 3960 9340 3990
rect 9460 4330 9560 4360
rect 9660 4330 9760 4360
rect 9460 4290 9490 4330
rect 9530 4290 9560 4330
rect 9660 4290 9690 4330
rect 9730 4290 9760 4330
rect 9460 4230 9560 4290
rect 9660 4230 9760 4290
rect 9460 4190 9490 4230
rect 9530 4190 9560 4230
rect 9660 4190 9690 4230
rect 9730 4190 9760 4230
rect 9460 4130 9560 4190
rect 9660 4130 9760 4190
rect 9460 4090 9490 4130
rect 9530 4090 9560 4130
rect 9660 4090 9690 4130
rect 9730 4090 9760 4130
rect 9460 4030 9560 4090
rect 9660 4030 9760 4090
rect 9460 3990 9490 4030
rect 9530 3990 9560 4030
rect 9660 3990 9690 4030
rect 9730 3990 9760 4030
rect 9460 3960 9560 3990
rect 9660 3960 9760 3990
rect 9880 4330 9980 4360
rect 9880 4290 9910 4330
rect 9950 4290 9980 4330
rect 9880 4230 9980 4290
rect 9880 4190 9910 4230
rect 9950 4190 9980 4230
rect 9880 4130 9980 4190
rect 9880 4090 9910 4130
rect 9950 4090 9980 4130
rect 9880 4030 9980 4090
rect 9880 3990 9910 4030
rect 9950 3990 9980 4030
rect 9880 3960 9980 3990
rect 10100 4330 10200 4360
rect 10100 4290 10130 4330
rect 10170 4290 10200 4330
rect 10100 4230 10200 4290
rect 10100 4190 10130 4230
rect 10170 4190 10200 4230
rect 10100 4130 10200 4190
rect 10100 4090 10130 4130
rect 10170 4090 10200 4130
rect 10100 4030 10200 4090
rect 10100 3990 10130 4030
rect 10170 3990 10200 4030
rect 10100 3960 10200 3990
rect 10320 4330 10420 4360
rect 10320 4290 10350 4330
rect 10390 4290 10420 4330
rect 10320 4230 10420 4290
rect 10320 4190 10350 4230
rect 10390 4190 10420 4230
rect 10320 4130 10420 4190
rect 10320 4090 10350 4130
rect 10390 4090 10420 4130
rect 10320 4030 10420 4090
rect 10320 3990 10350 4030
rect 10390 3990 10420 4030
rect 10320 3960 10420 3990
rect 10540 4330 10640 4360
rect 10540 4290 10570 4330
rect 10610 4290 10640 4330
rect 10540 4230 10640 4290
rect 10540 4190 10570 4230
rect 10610 4190 10640 4230
rect 10540 4130 10640 4190
rect 10540 4090 10570 4130
rect 10610 4090 10640 4130
rect 10540 4030 10640 4090
rect 10540 3990 10570 4030
rect 10610 3990 10640 4030
rect 10540 3960 10640 3990
rect 10760 4330 10860 4360
rect 10760 4290 10790 4330
rect 10830 4290 10860 4330
rect 10760 4230 10860 4290
rect 10760 4190 10790 4230
rect 10830 4190 10860 4230
rect 10760 4130 10860 4190
rect 10760 4090 10790 4130
rect 10830 4090 10860 4130
rect 10760 4030 10860 4090
rect 10760 3990 10790 4030
rect 10830 3990 10860 4030
rect 10760 3960 10860 3990
rect 10980 4330 11080 4360
rect 10980 4290 11010 4330
rect 11050 4290 11080 4330
rect 10980 4230 11080 4290
rect 10980 4190 11010 4230
rect 11050 4190 11080 4230
rect 10980 4130 11080 4190
rect 10980 4090 11010 4130
rect 11050 4090 11080 4130
rect 10980 4030 11080 4090
rect 10980 3990 11010 4030
rect 11050 3990 11080 4030
rect 10980 3960 11080 3990
rect 6860 3910 6960 3940
rect 2140 3520 2220 3550
rect 2140 3480 2160 3520
rect 2200 3480 2220 3520
rect 2140 3420 2220 3480
rect 2140 3380 2160 3420
rect 2200 3380 2220 3420
rect 2140 3320 2220 3380
rect 2140 3280 2160 3320
rect 2200 3280 2220 3320
rect 2140 3220 2220 3280
rect 2140 3180 2160 3220
rect 2200 3180 2220 3220
rect 2140 3150 2220 3180
rect 2250 3520 2330 3550
rect 2250 3480 2270 3520
rect 2310 3480 2330 3520
rect 2250 3420 2330 3480
rect 2250 3380 2270 3420
rect 2310 3380 2330 3420
rect 2250 3320 2330 3380
rect 2250 3280 2270 3320
rect 2310 3280 2330 3320
rect 2250 3220 2330 3280
rect 2250 3180 2270 3220
rect 2310 3180 2330 3220
rect 2250 3150 2330 3180
rect 2360 3520 2440 3550
rect 2360 3480 2380 3520
rect 2420 3480 2440 3520
rect 2360 3420 2440 3480
rect 2360 3380 2380 3420
rect 2420 3380 2440 3420
rect 2360 3320 2440 3380
rect 2360 3280 2380 3320
rect 2420 3280 2440 3320
rect 2360 3220 2440 3280
rect 2360 3180 2380 3220
rect 2420 3180 2440 3220
rect 2360 3150 2440 3180
rect 2660 3520 2740 3550
rect 2660 3480 2680 3520
rect 2720 3480 2740 3520
rect 2660 3420 2740 3480
rect 2660 3380 2680 3420
rect 2720 3380 2740 3420
rect 2660 3320 2740 3380
rect 2660 3280 2680 3320
rect 2720 3280 2740 3320
rect 2660 3220 2740 3280
rect 2660 3180 2680 3220
rect 2720 3180 2740 3220
rect 2660 3150 2740 3180
rect 2770 3520 2850 3550
rect 2770 3480 2790 3520
rect 2830 3480 2850 3520
rect 2770 3420 2850 3480
rect 2770 3380 2790 3420
rect 2830 3380 2850 3420
rect 2770 3320 2850 3380
rect 2770 3280 2790 3320
rect 2830 3280 2850 3320
rect 2770 3220 2850 3280
rect 2770 3180 2790 3220
rect 2830 3180 2850 3220
rect 2770 3150 2850 3180
rect 2880 3520 2960 3550
rect 3040 3520 3120 3550
rect 2880 3480 2900 3520
rect 2940 3480 2960 3520
rect 3040 3480 3060 3520
rect 3100 3480 3120 3520
rect 2880 3420 2960 3480
rect 3040 3420 3120 3480
rect 2880 3380 2900 3420
rect 2940 3380 2960 3420
rect 3040 3380 3060 3420
rect 3100 3380 3120 3420
rect 2880 3320 2960 3380
rect 3040 3320 3120 3380
rect 2880 3280 2900 3320
rect 2940 3280 2960 3320
rect 3040 3280 3060 3320
rect 3100 3280 3120 3320
rect 2880 3220 2960 3280
rect 3040 3220 3120 3280
rect 2880 3180 2900 3220
rect 2940 3180 2960 3220
rect 3040 3180 3060 3220
rect 3100 3180 3120 3220
rect 2880 3150 2960 3180
rect 3040 3150 3120 3180
rect 3150 3520 3230 3550
rect 3150 3480 3170 3520
rect 3210 3480 3230 3520
rect 3150 3420 3230 3480
rect 3150 3380 3170 3420
rect 3210 3380 3230 3420
rect 3150 3320 3230 3380
rect 3150 3280 3170 3320
rect 3210 3280 3230 3320
rect 3150 3220 3230 3280
rect 3150 3180 3170 3220
rect 3210 3180 3230 3220
rect 3150 3150 3230 3180
rect 3260 3520 3340 3550
rect 3260 3480 3280 3520
rect 3320 3480 3340 3520
rect 3260 3420 3340 3480
rect 3260 3380 3280 3420
rect 3320 3380 3340 3420
rect 3260 3320 3340 3380
rect 3260 3280 3280 3320
rect 3320 3280 3340 3320
rect 3260 3220 3340 3280
rect 3260 3180 3280 3220
rect 3320 3180 3340 3220
rect 3260 3150 3340 3180
rect 3560 3520 3640 3550
rect 3560 3480 3580 3520
rect 3620 3480 3640 3520
rect 3560 3420 3640 3480
rect 3560 3380 3580 3420
rect 3620 3380 3640 3420
rect 3560 3320 3640 3380
rect 3560 3280 3580 3320
rect 3620 3280 3640 3320
rect 3560 3220 3640 3280
rect 3560 3180 3580 3220
rect 3620 3180 3640 3220
rect 3560 3150 3640 3180
rect 3670 3520 3750 3550
rect 3670 3480 3690 3520
rect 3730 3480 3750 3520
rect 3670 3420 3750 3480
rect 3670 3380 3690 3420
rect 3730 3380 3750 3420
rect 3670 3320 3750 3380
rect 3670 3280 3690 3320
rect 3730 3280 3750 3320
rect 3670 3220 3750 3280
rect 3670 3180 3690 3220
rect 3730 3180 3750 3220
rect 3670 3150 3750 3180
rect 3780 3520 3860 3550
rect 3780 3480 3800 3520
rect 3840 3480 3860 3520
rect 3780 3420 3860 3480
rect 3780 3380 3800 3420
rect 3840 3380 3860 3420
rect 3780 3320 3860 3380
rect 3780 3280 3800 3320
rect 3840 3280 3860 3320
rect 3780 3220 3860 3280
rect 3780 3180 3800 3220
rect 3840 3180 3860 3220
rect 3780 3150 3860 3180
rect 4070 3520 4150 3550
rect 4070 3480 4090 3520
rect 4130 3480 4150 3520
rect 4070 3420 4150 3480
rect 4070 3380 4090 3420
rect 4130 3380 4150 3420
rect 4070 3320 4150 3380
rect 4070 3280 4090 3320
rect 4130 3280 4150 3320
rect 4070 3220 4150 3280
rect 4070 3180 4090 3220
rect 4130 3180 4150 3220
rect 4070 3150 4150 3180
rect 4180 3520 4260 3550
rect 4180 3480 4200 3520
rect 4240 3480 4260 3520
rect 4180 3420 4260 3480
rect 4180 3380 4200 3420
rect 4240 3380 4260 3420
rect 4180 3320 4260 3380
rect 4180 3280 4200 3320
rect 4240 3280 4260 3320
rect 4180 3220 4260 3280
rect 4180 3180 4200 3220
rect 4240 3180 4260 3220
rect 4180 3150 4260 3180
rect 4400 3520 4480 3550
rect 4400 3480 4420 3520
rect 4460 3480 4480 3520
rect 4400 3420 4480 3480
rect 4400 3380 4420 3420
rect 4460 3380 4480 3420
rect 4400 3320 4480 3380
rect 4400 3280 4420 3320
rect 4460 3280 4480 3320
rect 4400 3220 4480 3280
rect 4400 3180 4420 3220
rect 4460 3180 4480 3220
rect 4400 3150 4480 3180
rect 4510 3520 4590 3550
rect 4510 3480 4530 3520
rect 4570 3480 4590 3520
rect 4510 3420 4590 3480
rect 4510 3380 4530 3420
rect 4570 3380 4590 3420
rect 4510 3320 4590 3380
rect 4510 3280 4530 3320
rect 4570 3280 4590 3320
rect 4510 3220 4590 3280
rect 4510 3180 4530 3220
rect 4570 3180 4590 3220
rect 4510 3150 4590 3180
rect 4730 3520 4810 3550
rect 4730 3480 4750 3520
rect 4790 3480 4810 3520
rect 4730 3420 4810 3480
rect 4730 3380 4750 3420
rect 4790 3380 4810 3420
rect 4730 3320 4810 3380
rect 4730 3280 4750 3320
rect 4790 3280 4810 3320
rect 4730 3220 4810 3280
rect 4730 3180 4750 3220
rect 4790 3180 4810 3220
rect 4730 3150 4810 3180
rect 4840 3520 4920 3550
rect 4840 3480 4860 3520
rect 4900 3480 4920 3520
rect 4840 3420 4920 3480
rect 4840 3380 4860 3420
rect 4900 3380 4920 3420
rect 4840 3320 4920 3380
rect 4840 3280 4860 3320
rect 4900 3280 4920 3320
rect 4840 3220 4920 3280
rect 4840 3180 4860 3220
rect 4900 3180 4920 3220
rect 4840 3150 4920 3180
rect 5270 3520 5370 3550
rect 5270 3480 5300 3520
rect 5340 3480 5370 3520
rect 5270 3420 5370 3480
rect 5270 3380 5300 3420
rect 5340 3380 5370 3420
rect 5270 3320 5370 3380
rect 5270 3280 5300 3320
rect 5340 3280 5370 3320
rect 5270 3220 5370 3280
rect 5270 3180 5300 3220
rect 5340 3180 5370 3220
rect 5270 3150 5370 3180
rect 5400 3520 5500 3550
rect 5400 3480 5430 3520
rect 5470 3480 5500 3520
rect 5400 3420 5500 3480
rect 5400 3380 5430 3420
rect 5470 3380 5500 3420
rect 5400 3320 5500 3380
rect 5400 3280 5430 3320
rect 5470 3280 5500 3320
rect 5400 3220 5500 3280
rect 5400 3180 5430 3220
rect 5470 3180 5500 3220
rect 5400 3150 5500 3180
rect 5660 3520 5760 3550
rect 5660 3480 5690 3520
rect 5730 3480 5760 3520
rect 5660 3420 5760 3480
rect 5660 3380 5690 3420
rect 5730 3380 5760 3420
rect 5660 3320 5760 3380
rect 5660 3280 5690 3320
rect 5730 3280 5760 3320
rect 5660 3220 5760 3280
rect 5660 3180 5690 3220
rect 5730 3180 5760 3220
rect 5660 3150 5760 3180
rect 5790 3520 5890 3550
rect 5790 3480 5820 3520
rect 5860 3480 5890 3520
rect 5790 3420 5890 3480
rect 5790 3380 5820 3420
rect 5860 3380 5890 3420
rect 5790 3320 5890 3380
rect 5790 3280 5820 3320
rect 5860 3280 5890 3320
rect 5790 3220 5890 3280
rect 5790 3180 5820 3220
rect 5860 3180 5890 3220
rect 5790 3150 5890 3180
rect 6050 3520 6150 3550
rect 6050 3480 6080 3520
rect 6120 3480 6150 3520
rect 6050 3420 6150 3480
rect 6050 3380 6080 3420
rect 6120 3380 6150 3420
rect 6050 3320 6150 3380
rect 6050 3280 6080 3320
rect 6120 3280 6150 3320
rect 6050 3220 6150 3280
rect 6050 3180 6080 3220
rect 6120 3180 6150 3220
rect 6050 3150 6150 3180
rect 6180 3520 6280 3550
rect 6180 3480 6210 3520
rect 6250 3480 6280 3520
rect 6180 3420 6280 3480
rect 6180 3380 6210 3420
rect 6250 3380 6280 3420
rect 6180 3320 6280 3380
rect 6180 3280 6210 3320
rect 6250 3280 6280 3320
rect 6180 3220 6280 3280
rect 6180 3180 6210 3220
rect 6250 3180 6280 3220
rect 6180 3150 6280 3180
rect 6340 3520 6440 3550
rect 6340 3480 6370 3520
rect 6410 3480 6440 3520
rect 6340 3420 6440 3480
rect 6340 3380 6370 3420
rect 6410 3380 6440 3420
rect 6340 3320 6440 3380
rect 6340 3280 6370 3320
rect 6410 3280 6440 3320
rect 6340 3220 6440 3280
rect 6340 3180 6370 3220
rect 6410 3180 6440 3220
rect 6340 3150 6440 3180
rect 6470 3520 6570 3550
rect 6470 3480 6500 3520
rect 6540 3480 6570 3520
rect 6470 3420 6570 3480
rect 6470 3380 6500 3420
rect 6540 3380 6570 3420
rect 6470 3320 6570 3380
rect 6470 3280 6500 3320
rect 6540 3280 6570 3320
rect 6470 3220 6570 3280
rect 6470 3180 6500 3220
rect 6540 3180 6570 3220
rect 6470 3150 6570 3180
rect 1990 1090 2070 1120
rect 1990 1050 2010 1090
rect 2050 1050 2070 1090
rect 1990 1020 2070 1050
rect 2100 1090 2180 1120
rect 2100 1050 2120 1090
rect 2160 1050 2180 1090
rect 2100 1020 2180 1050
rect 2410 1090 2490 1120
rect 2410 1050 2430 1090
rect 2470 1050 2490 1090
rect 2410 1020 2490 1050
rect 2520 1090 2600 1120
rect 2520 1050 2540 1090
rect 2580 1050 2600 1090
rect 2520 1020 2600 1050
rect 2630 1090 2710 1120
rect 2630 1050 2650 1090
rect 2690 1050 2710 1090
rect 2630 1020 2710 1050
rect 3080 1090 3160 1120
rect 3080 1050 3100 1090
rect 3140 1050 3160 1090
rect 3080 1020 3160 1050
rect 3190 1090 3270 1120
rect 3190 1050 3210 1090
rect 3250 1050 3270 1090
rect 3190 1020 3270 1050
rect 3300 1090 3380 1120
rect 3300 1050 3320 1090
rect 3360 1050 3380 1090
rect 3300 1020 3380 1050
rect 3520 1090 3600 1120
rect 3520 1050 3540 1090
rect 3580 1050 3600 1090
rect 3520 1020 3600 1050
rect 3630 1090 3710 1120
rect 3630 1050 3650 1090
rect 3690 1050 3710 1090
rect 3630 1020 3710 1050
rect 3740 1090 3820 1120
rect 3740 1050 3760 1090
rect 3800 1050 3820 1090
rect 3740 1020 3820 1050
rect 3850 1090 3930 1120
rect 3850 1050 3870 1090
rect 3910 1050 3930 1090
rect 3850 1020 3930 1050
rect 4360 1090 4440 1120
rect 4360 1050 4380 1090
rect 4420 1050 4440 1090
rect 4360 1020 4440 1050
rect 4470 1090 4550 1120
rect 4470 1050 4490 1090
rect 4530 1050 4550 1090
rect 4470 1020 4550 1050
rect 4780 1090 4860 1120
rect 4780 1050 4800 1090
rect 4840 1050 4860 1090
rect 4780 1020 4860 1050
rect 4890 1090 4970 1120
rect 4890 1050 4910 1090
rect 4950 1050 4970 1090
rect 4890 1020 4970 1050
rect 5000 1090 5080 1120
rect 5000 1050 5020 1090
rect 5060 1050 5080 1090
rect 5000 1020 5080 1050
rect 5230 1090 5310 1120
rect 5230 1050 5250 1090
rect 5290 1050 5310 1090
rect 5230 1020 5310 1050
rect 5340 1090 5420 1120
rect 5340 1050 5360 1090
rect 5400 1050 5420 1090
rect 5340 1020 5420 1050
rect 5450 1090 5530 1120
rect 5450 1050 5470 1090
rect 5510 1050 5530 1090
rect 5450 1020 5530 1050
rect 5590 1090 5670 1120
rect 5590 1050 5610 1090
rect 5650 1050 5670 1090
rect 5590 1020 5670 1050
rect 5700 1090 5780 1120
rect 5700 1050 5720 1090
rect 5760 1050 5780 1090
rect 5700 1020 5780 1050
rect 5810 1090 5890 1120
rect 5810 1050 5830 1090
rect 5870 1050 5890 1090
rect 5810 1020 5890 1050
rect 6170 1090 6250 1120
rect 6170 1050 6190 1090
rect 6230 1050 6250 1090
rect 6170 1020 6250 1050
rect 6280 1090 6360 1120
rect 6280 1050 6300 1090
rect 6340 1050 6360 1090
rect 6280 1020 6360 1050
rect 6390 1090 6470 1120
rect 6390 1050 6410 1090
rect 6450 1050 6470 1090
rect 6390 1020 6470 1050
rect 6610 1090 6690 1120
rect 6610 1050 6630 1090
rect 6670 1050 6690 1090
rect 6610 1020 6690 1050
rect 6720 1090 6800 1120
rect 6720 1050 6740 1090
rect 6780 1050 6800 1090
rect 6720 1020 6800 1050
rect 6830 1090 6910 1120
rect 6830 1050 6850 1090
rect 6890 1050 6910 1090
rect 12400 1190 12480 1220
rect 12400 1150 12420 1190
rect 12460 1150 12480 1190
rect 6830 1020 6910 1050
rect 7230 1090 7310 1120
rect 7230 1050 7250 1090
rect 7290 1050 7310 1090
rect 7230 1020 7310 1050
rect 7340 1090 7420 1120
rect 7340 1050 7360 1090
rect 7400 1050 7420 1090
rect 7340 1020 7420 1050
rect 7570 1090 7650 1120
rect 7570 1050 7590 1090
rect 7630 1050 7650 1090
rect 7570 1020 7650 1050
rect 7680 1090 7760 1120
rect 7680 1050 7700 1090
rect 7740 1050 7760 1090
rect 7680 1020 7760 1050
rect 7790 1090 7870 1120
rect 7790 1050 7810 1090
rect 7850 1050 7870 1090
rect 7790 1020 7870 1050
rect 7930 1090 8010 1120
rect 7930 1050 7950 1090
rect 7990 1050 8010 1090
rect 7930 1020 8010 1050
rect 8040 1090 8120 1120
rect 8040 1050 8060 1090
rect 8100 1050 8120 1090
rect 8040 1020 8120 1050
rect 8150 1090 8230 1120
rect 8150 1050 8170 1090
rect 8210 1050 8230 1090
rect 8150 1020 8230 1050
rect 8530 1090 8610 1120
rect 8530 1050 8550 1090
rect 8590 1050 8610 1090
rect 8530 1020 8610 1050
rect 8640 1090 8720 1120
rect 8640 1050 8660 1090
rect 8700 1050 8720 1090
rect 8640 1020 8720 1050
rect 8870 1090 8950 1120
rect 8870 1050 8890 1090
rect 8930 1050 8950 1090
rect 8870 1020 8950 1050
rect 8980 1090 9060 1120
rect 8980 1050 9000 1090
rect 9040 1050 9060 1090
rect 8980 1020 9060 1050
rect 9090 1090 9170 1120
rect 9090 1050 9110 1090
rect 9150 1050 9170 1090
rect 9090 1020 9170 1050
rect 9230 1090 9310 1120
rect 9230 1050 9250 1090
rect 9290 1050 9310 1090
rect 9230 1020 9310 1050
rect 9340 1090 9420 1120
rect 9340 1050 9360 1090
rect 9400 1050 9420 1090
rect 9340 1020 9420 1050
rect 9450 1090 9530 1120
rect 9450 1050 9470 1090
rect 9510 1050 9530 1090
rect 9450 1020 9530 1050
rect 9830 1090 9910 1120
rect 9830 1050 9850 1090
rect 9890 1050 9910 1090
rect 9830 1020 9910 1050
rect 9940 1090 10020 1120
rect 9940 1050 9960 1090
rect 10000 1050 10020 1090
rect 9940 1020 10020 1050
rect 10170 1090 10250 1120
rect 10170 1050 10190 1090
rect 10230 1050 10250 1090
rect 10170 1020 10250 1050
rect 10280 1090 10360 1120
rect 10280 1050 10300 1090
rect 10340 1050 10360 1090
rect 10280 1020 10360 1050
rect 10390 1090 10470 1120
rect 10390 1050 10410 1090
rect 10450 1050 10470 1090
rect 10390 1020 10470 1050
rect 10530 1090 10610 1120
rect 10530 1050 10550 1090
rect 10590 1050 10610 1090
rect 10530 1020 10610 1050
rect 10640 1090 10720 1120
rect 10640 1050 10660 1090
rect 10700 1050 10720 1090
rect 10640 1020 10720 1050
rect 10750 1090 10830 1120
rect 10750 1050 10770 1090
rect 10810 1050 10830 1090
rect 10750 1020 10830 1050
rect 11130 1090 11210 1120
rect 11130 1050 11150 1090
rect 11190 1050 11210 1090
rect 11130 1020 11210 1050
rect 11240 1090 11320 1120
rect 11240 1050 11260 1090
rect 11300 1050 11320 1090
rect 11240 1020 11320 1050
rect 11470 1090 11550 1120
rect 11470 1050 11490 1090
rect 11530 1050 11550 1090
rect 11470 1020 11550 1050
rect 11580 1090 11660 1120
rect 11580 1050 11600 1090
rect 11640 1050 11660 1090
rect 11580 1020 11660 1050
rect 11690 1090 11770 1120
rect 11690 1050 11710 1090
rect 11750 1050 11770 1090
rect 11690 1020 11770 1050
rect 11830 1090 11910 1120
rect 11830 1050 11850 1090
rect 11890 1050 11910 1090
rect 11830 1020 11910 1050
rect 11940 1090 12020 1120
rect 11940 1050 11960 1090
rect 12000 1050 12020 1090
rect 11940 1020 12020 1050
rect 12050 1090 12130 1120
rect 12050 1050 12070 1090
rect 12110 1050 12130 1090
rect 12050 1020 12130 1050
rect 12400 1090 12480 1150
rect 12400 1050 12420 1090
rect 12460 1050 12480 1090
rect 12400 1020 12480 1050
rect 12510 1190 12590 1220
rect 12510 1150 12530 1190
rect 12570 1150 12590 1190
rect 12510 1090 12590 1150
rect 12510 1050 12530 1090
rect 12570 1050 12590 1090
rect 12510 1020 12590 1050
rect 13000 1190 13080 1220
rect 13000 1150 13020 1190
rect 13060 1150 13080 1190
rect 13000 1090 13080 1150
rect 13000 1050 13020 1090
rect 13060 1050 13080 1090
rect 13000 1020 13080 1050
rect 13110 1190 13190 1220
rect 13110 1150 13130 1190
rect 13170 1150 13190 1190
rect 13110 1090 13190 1150
rect 13110 1050 13130 1090
rect 13170 1050 13190 1090
rect 13110 1020 13190 1050
rect 13600 1190 13680 1220
rect 13600 1150 13620 1190
rect 13660 1150 13680 1190
rect 13600 1090 13680 1150
rect 13600 1050 13620 1090
rect 13660 1050 13680 1090
rect 13600 1020 13680 1050
rect 13710 1190 13790 1220
rect 13710 1150 13730 1190
rect 13770 1150 13790 1190
rect 13710 1090 13790 1150
rect 13710 1050 13730 1090
rect 13770 1050 13790 1090
rect 13710 1020 13790 1050
rect 12400 850 12480 880
rect 12400 810 12420 850
rect 12460 810 12480 850
rect 12400 750 12480 810
rect 12400 710 12420 750
rect 12460 710 12480 750
rect 12400 680 12480 710
rect 12510 850 12590 880
rect 12510 810 12530 850
rect 12570 810 12590 850
rect 12510 750 12590 810
rect 12510 710 12530 750
rect 12570 710 12590 750
rect 12510 680 12590 710
rect 13000 850 13080 880
rect 13000 810 13020 850
rect 13060 810 13080 850
rect 13000 750 13080 810
rect 13000 710 13020 750
rect 13060 710 13080 750
rect 13000 680 13080 710
rect 13110 850 13190 880
rect 13110 810 13130 850
rect 13170 810 13190 850
rect 13110 750 13190 810
rect 13110 710 13130 750
rect 13170 710 13190 750
rect 13110 680 13190 710
rect 13600 850 13680 880
rect 13600 810 13620 850
rect 13660 810 13680 850
rect 13600 750 13680 810
rect 13600 710 13620 750
rect 13660 710 13680 750
rect 13600 680 13680 710
rect 13710 850 13790 880
rect 13710 810 13730 850
rect 13770 810 13790 850
rect 13710 750 13790 810
rect 13710 710 13730 750
rect 13770 710 13790 750
rect 13710 680 13790 710
rect 12400 500 12480 530
rect 12400 460 12420 500
rect 12460 460 12480 500
rect 12400 400 12480 460
rect 12400 360 12420 400
rect 12460 360 12480 400
rect 12400 300 12480 360
rect 12400 260 12420 300
rect 12460 260 12480 300
rect 12400 200 12480 260
rect 12400 160 12420 200
rect 12460 160 12480 200
rect 12400 130 12480 160
rect 12780 500 12860 530
rect 12780 460 12800 500
rect 12840 460 12860 500
rect 12780 400 12860 460
rect 12780 360 12800 400
rect 12840 360 12860 400
rect 12780 300 12860 360
rect 12780 260 12800 300
rect 12840 260 12860 300
rect 12780 200 12860 260
rect 12780 160 12800 200
rect 12840 160 12860 200
rect 12780 130 12860 160
rect 13000 500 13080 530
rect 13000 460 13020 500
rect 13060 460 13080 500
rect 13000 400 13080 460
rect 13000 360 13020 400
rect 13060 360 13080 400
rect 13000 300 13080 360
rect 13000 260 13020 300
rect 13060 260 13080 300
rect 13000 200 13080 260
rect 13000 160 13020 200
rect 13060 160 13080 200
rect 13000 130 13080 160
rect 13380 500 13460 530
rect 13380 460 13400 500
rect 13440 460 13460 500
rect 13380 400 13460 460
rect 13380 360 13400 400
rect 13440 360 13460 400
rect 13380 300 13460 360
rect 13380 260 13400 300
rect 13440 260 13460 300
rect 13380 200 13460 260
rect 13380 160 13400 200
rect 13440 160 13460 200
rect 13380 130 13460 160
rect 13600 500 13680 530
rect 13600 460 13620 500
rect 13660 460 13680 500
rect 13600 400 13680 460
rect 13600 360 13620 400
rect 13660 360 13680 400
rect 13600 300 13680 360
rect 13600 260 13620 300
rect 13660 260 13680 300
rect 13600 200 13680 260
rect 13600 160 13620 200
rect 13660 160 13680 200
rect 13600 130 13680 160
rect 13980 500 14060 530
rect 14140 500 14220 530
rect 13980 460 14000 500
rect 14040 460 14060 500
rect 14140 460 14160 500
rect 14200 460 14220 500
rect 13980 400 14060 460
rect 14140 400 14220 460
rect 13980 360 14000 400
rect 14040 360 14060 400
rect 14140 360 14160 400
rect 14200 360 14220 400
rect 13980 300 14060 360
rect 14140 300 14220 360
rect 13980 260 14000 300
rect 14040 260 14060 300
rect 14140 260 14160 300
rect 14200 260 14220 300
rect 13980 200 14060 260
rect 14140 200 14220 260
rect 13980 160 14000 200
rect 14040 160 14060 200
rect 14140 160 14160 200
rect 14200 160 14220 200
rect 13980 130 14060 160
rect 14140 130 14220 160
rect 14520 500 14600 530
rect 14520 460 14540 500
rect 14580 460 14600 500
rect 14520 400 14600 460
rect 14520 360 14540 400
rect 14580 360 14600 400
rect 14520 300 14600 360
rect 14520 260 14540 300
rect 14580 260 14600 300
rect 14520 200 14600 260
rect 14520 160 14540 200
rect 14580 160 14600 200
rect 14520 130 14600 160
<< ndiffc >>
rect 1170 10220 1210 10260
rect 1170 10120 1210 10160
rect 3250 10220 3290 10260
rect 3250 10120 3290 10160
rect 5330 10220 5370 10260
rect 5330 10120 5370 10160
rect 750 9610 790 9650
rect 750 9510 790 9550
rect 750 9410 790 9450
rect 750 9310 790 9350
rect 750 9210 790 9250
rect 1830 9610 1870 9650
rect 1990 9610 2030 9650
rect 1830 9510 1870 9550
rect 1990 9510 2030 9550
rect 1830 9410 1870 9450
rect 1990 9410 2030 9450
rect 1830 9310 1870 9350
rect 1990 9310 2030 9350
rect 1830 9210 1870 9250
rect 1990 9210 2030 9250
rect 3070 9610 3110 9650
rect 3070 9510 3110 9550
rect 3070 9410 3110 9450
rect 3070 9310 3110 9350
rect 3070 9210 3110 9250
rect 3430 9610 3470 9650
rect 3430 9510 3470 9550
rect 3430 9410 3470 9450
rect 3430 9310 3470 9350
rect 3430 9210 3470 9250
rect 4510 9610 4550 9650
rect 4670 9610 4710 9650
rect 4510 9510 4550 9550
rect 4670 9510 4710 9550
rect 4510 9410 4550 9450
rect 4670 9410 4710 9450
rect 4510 9310 4550 9350
rect 4670 9310 4710 9350
rect 4510 9210 4550 9250
rect 4670 9210 4710 9250
rect 5750 9610 5790 9650
rect 5750 9510 5790 9550
rect 5750 9410 5790 9450
rect 5750 9310 5790 9350
rect 5750 9210 5790 9250
rect 1370 8600 1410 8640
rect 1490 8600 1530 8640
rect 1610 8600 1650 8640
rect 1730 8600 1770 8640
rect 1850 8600 1890 8640
rect 1970 8600 2010 8640
rect 2090 8600 2130 8640
rect 2210 8600 2250 8640
rect 2330 8600 2370 8640
rect 2450 8600 2490 8640
rect 2570 8600 2610 8640
rect 3930 8600 3970 8640
rect 4050 8600 4090 8640
rect 4170 8600 4210 8640
rect 4290 8600 4330 8640
rect 4410 8600 4450 8640
rect 4530 8600 4570 8640
rect 4650 8600 4690 8640
rect 4770 8600 4810 8640
rect 4890 8600 4930 8640
rect 5010 8600 5050 8640
rect 5130 8600 5170 8640
rect 8230 8530 8270 8580
rect 8230 8390 8270 8440
rect 8430 8530 8470 8580
rect 8430 8390 8470 8440
rect 8630 8530 8670 8580
rect 8630 8390 8670 8440
rect 8830 8530 8870 8580
rect 8830 8390 8870 8440
rect 9030 8530 9070 8580
rect 9030 8390 9070 8440
rect 9230 8530 9270 8580
rect 9230 8390 9270 8440
rect 9430 8530 9470 8580
rect 9430 8390 9470 8440
rect 9630 8530 9670 8580
rect 9630 8390 9670 8440
rect 9830 8530 9870 8580
rect 9830 8390 9870 8440
rect 10030 8530 10070 8580
rect 10030 8390 10070 8440
rect 10230 8530 10270 8580
rect 10230 8390 10270 8440
rect 8280 7850 8320 7890
rect 8410 7850 8450 7890
rect 8540 7850 8580 7890
rect 8670 7850 8710 7890
rect 8800 7850 8840 7890
rect 8930 7850 8970 7890
rect 9060 7850 9100 7890
rect 9420 7850 9460 7890
rect 9550 7850 9590 7890
rect 9680 7850 9720 7890
rect 9810 7850 9850 7890
rect 9940 7850 9980 7890
rect 10070 7850 10110 7890
rect 10200 7850 10240 7890
rect 10560 7850 10600 7890
rect 10690 7850 10730 7890
rect 10820 7850 10860 7890
rect 10950 7850 10990 7890
rect 11080 7850 11120 7890
rect 11210 7850 11250 7890
rect 11340 7850 11380 7890
rect 2160 4660 2200 4700
rect 2160 4560 2200 4600
rect 2270 4660 2310 4700
rect 2270 4560 2310 4600
rect 2380 4660 2420 4700
rect 2380 4560 2420 4600
rect 2680 4660 2720 4700
rect 2680 4560 2720 4600
rect 2790 4660 2830 4700
rect 2790 4560 2830 4600
rect 2900 4660 2940 4700
rect 3060 4660 3100 4700
rect 2900 4560 2940 4600
rect 3060 4560 3100 4600
rect 3170 4660 3210 4700
rect 3170 4560 3210 4600
rect 3280 4660 3320 4700
rect 3280 4560 3320 4600
rect 3580 4660 3620 4700
rect 3580 4560 3620 4600
rect 3690 4660 3730 4700
rect 3690 4560 3730 4600
rect 3800 4660 3840 4700
rect 3800 4560 3840 4600
rect 4100 4660 4140 4700
rect 4100 4560 4140 4600
rect 4210 4660 4250 4700
rect 4210 4560 4250 4600
rect 4320 4660 4360 4700
rect 4320 4560 4360 4600
rect 4540 4660 4580 4700
rect 4540 4560 4580 4600
rect 4650 4660 4690 4700
rect 4650 4560 4690 4600
rect 4870 4660 4910 4700
rect 4870 4560 4910 4600
rect 4980 4660 5020 4700
rect 4980 4560 5020 4600
rect 5300 4660 5340 4700
rect 5300 4560 5340 4600
rect 5430 4660 5470 4700
rect 5430 4560 5470 4600
rect 5690 4660 5730 4700
rect 5690 4560 5730 4600
rect 5820 4660 5860 4700
rect 5820 4560 5860 4600
rect 6080 4660 6120 4700
rect 6080 4560 6120 4600
rect 6210 4660 6250 4700
rect 6210 4560 6250 4600
rect 6370 4660 6410 4700
rect 6370 4560 6410 4600
rect 6500 4660 6540 4700
rect 6500 4560 6540 4600
rect 7970 3310 8010 3350
rect 7970 3210 8010 3250
rect 7970 3110 8010 3150
rect 7970 3010 8010 3050
rect 8190 3310 8230 3350
rect 8190 3210 8230 3250
rect 8190 3110 8230 3150
rect 8190 3010 8230 3050
rect 8410 3310 8450 3350
rect 8410 3210 8450 3250
rect 8410 3110 8450 3150
rect 8410 3010 8450 3050
rect 8630 3310 8670 3350
rect 8630 3210 8670 3250
rect 8630 3110 8670 3150
rect 8630 3010 8670 3050
rect 8850 3310 8890 3350
rect 9050 3310 9090 3350
rect 8850 3210 8890 3250
rect 9050 3210 9090 3250
rect 8850 3110 8890 3150
rect 9050 3110 9090 3150
rect 8850 3010 8890 3050
rect 9050 3010 9090 3050
rect 9270 3310 9310 3350
rect 9270 3210 9310 3250
rect 9270 3110 9310 3150
rect 9270 3010 9310 3050
rect 9490 3310 9530 3350
rect 9490 3210 9530 3250
rect 9490 3110 9530 3150
rect 9490 3010 9530 3050
rect 9710 3310 9750 3350
rect 9710 3210 9750 3250
rect 9710 3110 9750 3150
rect 9710 3010 9750 3050
rect 9930 3310 9970 3350
rect 10130 3310 10170 3350
rect 9930 3210 9970 3250
rect 10130 3210 10170 3250
rect 9930 3110 9970 3150
rect 10130 3110 10170 3150
rect 9930 3010 9970 3050
rect 10130 3010 10170 3050
rect 10350 3310 10390 3350
rect 10350 3210 10390 3250
rect 10350 3110 10390 3150
rect 10350 3010 10390 3050
rect 10570 3310 10610 3350
rect 10570 3210 10610 3250
rect 10570 3110 10610 3150
rect 10570 3010 10610 3050
rect 10790 3310 10830 3350
rect 10790 3210 10830 3250
rect 10790 3110 10830 3150
rect 10790 3010 10830 3050
rect 11010 3310 11050 3350
rect 11010 3210 11050 3250
rect 11010 3110 11050 3150
rect 11010 3010 11050 3050
rect 2160 2860 2200 2900
rect 2160 2760 2200 2800
rect 2270 2860 2310 2900
rect 2270 2760 2310 2800
rect 2380 2860 2420 2900
rect 2380 2760 2420 2800
rect 2680 2860 2720 2900
rect 2680 2760 2720 2800
rect 2790 2860 2830 2900
rect 2790 2760 2830 2800
rect 2900 2860 2940 2900
rect 3060 2860 3100 2900
rect 2900 2760 2940 2800
rect 3060 2760 3100 2800
rect 3170 2860 3210 2900
rect 3170 2760 3210 2800
rect 3280 2860 3320 2900
rect 3280 2760 3320 2800
rect 3580 2860 3620 2900
rect 3580 2760 3620 2800
rect 3690 2860 3730 2900
rect 3690 2760 3730 2800
rect 3800 2860 3840 2900
rect 3800 2760 3840 2800
rect 4090 2860 4130 2900
rect 4090 2760 4130 2800
rect 4200 2860 4240 2900
rect 4200 2760 4240 2800
rect 4420 2860 4460 2900
rect 4420 2760 4460 2800
rect 4530 2860 4570 2900
rect 4530 2760 4570 2800
rect 4750 2860 4790 2900
rect 4750 2760 4790 2800
rect 4860 2860 4900 2900
rect 4860 2760 4900 2800
rect 5300 2860 5340 2900
rect 5300 2760 5340 2800
rect 5430 2860 5470 2900
rect 5430 2760 5470 2800
rect 5690 2860 5730 2900
rect 5690 2760 5730 2800
rect 5820 2860 5860 2900
rect 5820 2760 5860 2800
rect 6080 2860 6120 2900
rect 6080 2760 6120 2800
rect 6210 2860 6250 2900
rect 6210 2760 6250 2800
rect 6370 2860 6410 2900
rect 6370 2760 6410 2800
rect 6500 2860 6540 2900
rect 6500 2760 6540 2800
rect 6760 2860 6800 2900
rect 6760 2760 6800 2800
rect 6890 2860 6930 2900
rect 6890 2760 6930 2800
rect 12420 1930 12460 1970
rect 12420 1830 12460 1870
rect 12530 1930 12570 1970
rect 12530 1830 12570 1870
rect 13020 1930 13060 1970
rect 13020 1830 13060 1870
rect 13130 1930 13170 1970
rect 13130 1830 13170 1870
rect 13620 1930 13660 1970
rect 13620 1830 13660 1870
rect 13730 1930 13770 1970
rect 13890 1930 13930 1970
rect 13730 1830 13770 1870
rect 13890 1830 13930 1870
rect 14000 1930 14040 1970
rect 14000 1830 14040 1870
rect 12420 1600 12460 1640
rect 12530 1600 12570 1640
rect 13020 1600 13060 1640
rect 13130 1600 13170 1640
rect 13620 1600 13660 1640
rect 13730 1600 13770 1640
rect 1850 1370 1890 1410
rect 1960 1370 2000 1410
rect 2070 1370 2110 1410
rect 2180 1370 2220 1410
rect 2290 1370 2330 1410
rect 2430 1370 2470 1410
rect 2540 1370 2580 1410
rect 2650 1370 2690 1410
rect 2880 1370 2920 1410
rect 2990 1370 3030 1410
rect 3100 1370 3140 1410
rect 3210 1370 3250 1410
rect 3320 1370 3360 1410
rect 3540 1370 3580 1410
rect 3650 1370 3690 1410
rect 3760 1370 3800 1410
rect 3870 1370 3910 1410
rect 3980 1370 4020 1410
rect 4220 1370 4260 1410
rect 4330 1370 4370 1410
rect 4440 1370 4480 1410
rect 4550 1370 4590 1410
rect 4660 1370 4700 1410
rect 4800 1370 4840 1410
rect 4910 1370 4950 1410
rect 5020 1370 5060 1410
rect 5360 1370 5400 1410
rect 5470 1370 5510 1410
rect 5720 1370 5760 1410
rect 5830 1370 5870 1410
rect 5970 1370 6010 1410
rect 6080 1370 6120 1410
rect 6190 1370 6230 1410
rect 6300 1370 6340 1410
rect 6410 1370 6450 1410
rect 6630 1370 6670 1410
rect 6740 1370 6780 1410
rect 6850 1370 6890 1410
rect 6960 1370 7000 1410
rect 7180 1370 7220 1410
rect 7290 1370 7330 1410
rect 7400 1370 7440 1410
rect 7510 1370 7550 1410
rect 7620 1370 7660 1410
rect 7840 1370 7880 1410
rect 7950 1370 7990 1410
rect 8060 1370 8100 1410
rect 8480 1460 8520 1500
rect 8590 1460 8630 1500
rect 8700 1460 8740 1500
rect 8810 1460 8850 1500
rect 8920 1460 8960 1500
rect 9140 1460 9180 1500
rect 9250 1460 9290 1500
rect 9360 1460 9400 1500
rect 9470 1460 9510 1500
rect 9780 1460 9820 1500
rect 9890 1460 9930 1500
rect 10000 1460 10040 1500
rect 10110 1460 10150 1500
rect 10220 1460 10260 1500
rect 10440 1460 10480 1500
rect 10550 1460 10590 1500
rect 10660 1460 10700 1500
rect 10770 1460 10810 1500
rect 11080 1460 11120 1500
rect 11190 1460 11230 1500
rect 11300 1460 11340 1500
rect 11410 1460 11450 1500
rect 11520 1460 11560 1500
rect 11740 1460 11780 1500
rect 11850 1460 11890 1500
rect 11960 1460 12000 1500
rect 12070 1460 12110 1500
rect 8170 1370 8210 1410
rect 12420 1360 12460 1400
rect 12530 1360 12570 1400
rect 13020 1360 13060 1400
rect 13130 1360 13170 1400
rect 13620 1360 13660 1400
rect 13730 1360 13770 1400
<< pdiffc >>
rect 1622 14402 1656 14436
rect 1712 14402 1746 14436
rect 1802 14402 1836 14436
rect 1892 14402 1926 14436
rect 1982 14402 2016 14436
rect 2072 14402 2106 14436
rect 2162 14402 2196 14436
rect 1622 14312 1656 14346
rect 1712 14312 1746 14346
rect 1802 14312 1836 14346
rect 1892 14312 1926 14346
rect 1982 14312 2016 14346
rect 2072 14312 2106 14346
rect 2162 14312 2196 14346
rect 1622 14222 1656 14256
rect 1712 14222 1746 14256
rect 1802 14222 1836 14256
rect 1892 14222 1926 14256
rect 1982 14222 2016 14256
rect 2072 14222 2106 14256
rect 2162 14222 2196 14256
rect 1622 14132 1656 14166
rect 1712 14132 1746 14166
rect 1802 14132 1836 14166
rect 1892 14132 1926 14166
rect 1982 14132 2016 14166
rect 2072 14132 2106 14166
rect 2162 14132 2196 14166
rect 1622 14042 1656 14076
rect 1712 14042 1746 14076
rect 1802 14042 1836 14076
rect 1892 14042 1926 14076
rect 1982 14042 2016 14076
rect 2072 14042 2106 14076
rect 2162 14042 2196 14076
rect 1622 13952 1656 13986
rect 1712 13952 1746 13986
rect 1802 13952 1836 13986
rect 1892 13952 1926 13986
rect 1982 13952 2016 13986
rect 2072 13952 2106 13986
rect 2162 13952 2196 13986
rect 1622 13862 1656 13896
rect 1712 13862 1746 13896
rect 1802 13862 1836 13896
rect 1892 13862 1926 13896
rect 1982 13862 2016 13896
rect 2072 13862 2106 13896
rect 2162 13862 2196 13896
rect 2982 14402 3016 14436
rect 3072 14402 3106 14436
rect 3162 14402 3196 14436
rect 3252 14402 3286 14436
rect 3342 14402 3376 14436
rect 3432 14402 3466 14436
rect 3522 14402 3556 14436
rect 2982 14312 3016 14346
rect 3072 14312 3106 14346
rect 3162 14312 3196 14346
rect 3252 14312 3286 14346
rect 3342 14312 3376 14346
rect 3432 14312 3466 14346
rect 3522 14312 3556 14346
rect 2982 14222 3016 14256
rect 3072 14222 3106 14256
rect 3162 14222 3196 14256
rect 3252 14222 3286 14256
rect 3342 14222 3376 14256
rect 3432 14222 3466 14256
rect 3522 14222 3556 14256
rect 2982 14132 3016 14166
rect 3072 14132 3106 14166
rect 3162 14132 3196 14166
rect 3252 14132 3286 14166
rect 3342 14132 3376 14166
rect 3432 14132 3466 14166
rect 3522 14132 3556 14166
rect 2982 14042 3016 14076
rect 3072 14042 3106 14076
rect 3162 14042 3196 14076
rect 3252 14042 3286 14076
rect 3342 14042 3376 14076
rect 3432 14042 3466 14076
rect 3522 14042 3556 14076
rect 2982 13952 3016 13986
rect 3072 13952 3106 13986
rect 3162 13952 3196 13986
rect 3252 13952 3286 13986
rect 3342 13952 3376 13986
rect 3432 13952 3466 13986
rect 3522 13952 3556 13986
rect 2982 13862 3016 13896
rect 3072 13862 3106 13896
rect 3162 13862 3196 13896
rect 3252 13862 3286 13896
rect 3342 13862 3376 13896
rect 3432 13862 3466 13896
rect 3522 13862 3556 13896
rect 4342 14402 4376 14436
rect 4432 14402 4466 14436
rect 4522 14402 4556 14436
rect 4612 14402 4646 14436
rect 4702 14402 4736 14436
rect 4792 14402 4826 14436
rect 4882 14402 4916 14436
rect 4342 14312 4376 14346
rect 4432 14312 4466 14346
rect 4522 14312 4556 14346
rect 4612 14312 4646 14346
rect 4702 14312 4736 14346
rect 4792 14312 4826 14346
rect 4882 14312 4916 14346
rect 4342 14222 4376 14256
rect 4432 14222 4466 14256
rect 4522 14222 4556 14256
rect 4612 14222 4646 14256
rect 4702 14222 4736 14256
rect 4792 14222 4826 14256
rect 4882 14222 4916 14256
rect 4342 14132 4376 14166
rect 4432 14132 4466 14166
rect 4522 14132 4556 14166
rect 4612 14132 4646 14166
rect 4702 14132 4736 14166
rect 4792 14132 4826 14166
rect 4882 14132 4916 14166
rect 4342 14042 4376 14076
rect 4432 14042 4466 14076
rect 4522 14042 4556 14076
rect 4612 14042 4646 14076
rect 4702 14042 4736 14076
rect 4792 14042 4826 14076
rect 4882 14042 4916 14076
rect 4342 13952 4376 13986
rect 4432 13952 4466 13986
rect 4522 13952 4556 13986
rect 4612 13952 4646 13986
rect 4702 13952 4736 13986
rect 4792 13952 4826 13986
rect 4882 13952 4916 13986
rect 4342 13862 4376 13896
rect 4432 13862 4466 13896
rect 4522 13862 4556 13896
rect 4612 13862 4646 13896
rect 4702 13862 4736 13896
rect 4792 13862 4826 13896
rect 4882 13862 4916 13896
rect 1622 13042 1656 13076
rect 1712 13042 1746 13076
rect 1802 13042 1836 13076
rect 1892 13042 1926 13076
rect 1982 13042 2016 13076
rect 2072 13042 2106 13076
rect 2162 13042 2196 13076
rect 1622 12952 1656 12986
rect 1712 12952 1746 12986
rect 1802 12952 1836 12986
rect 1892 12952 1926 12986
rect 1982 12952 2016 12986
rect 2072 12952 2106 12986
rect 2162 12952 2196 12986
rect 1622 12862 1656 12896
rect 1712 12862 1746 12896
rect 1802 12862 1836 12896
rect 1892 12862 1926 12896
rect 1982 12862 2016 12896
rect 2072 12862 2106 12896
rect 2162 12862 2196 12896
rect 1622 12772 1656 12806
rect 1712 12772 1746 12806
rect 1802 12772 1836 12806
rect 1892 12772 1926 12806
rect 1982 12772 2016 12806
rect 2072 12772 2106 12806
rect 2162 12772 2196 12806
rect 1622 12682 1656 12716
rect 1712 12682 1746 12716
rect 1802 12682 1836 12716
rect 1892 12682 1926 12716
rect 1982 12682 2016 12716
rect 2072 12682 2106 12716
rect 2162 12682 2196 12716
rect 1622 12592 1656 12626
rect 1712 12592 1746 12626
rect 1802 12592 1836 12626
rect 1892 12592 1926 12626
rect 1982 12592 2016 12626
rect 2072 12592 2106 12626
rect 2162 12592 2196 12626
rect 1622 12502 1656 12536
rect 1712 12502 1746 12536
rect 1802 12502 1836 12536
rect 1892 12502 1926 12536
rect 1982 12502 2016 12536
rect 2072 12502 2106 12536
rect 2162 12502 2196 12536
rect 2982 13042 3016 13076
rect 3072 13042 3106 13076
rect 3162 13042 3196 13076
rect 3252 13042 3286 13076
rect 3342 13042 3376 13076
rect 3432 13042 3466 13076
rect 3522 13042 3556 13076
rect 2982 12952 3016 12986
rect 3072 12952 3106 12986
rect 3162 12952 3196 12986
rect 3252 12952 3286 12986
rect 3342 12952 3376 12986
rect 3432 12952 3466 12986
rect 3522 12952 3556 12986
rect 2982 12862 3016 12896
rect 3072 12862 3106 12896
rect 3162 12862 3196 12896
rect 3252 12862 3286 12896
rect 3342 12862 3376 12896
rect 3432 12862 3466 12896
rect 3522 12862 3556 12896
rect 2982 12772 3016 12806
rect 3072 12772 3106 12806
rect 3162 12772 3196 12806
rect 3252 12772 3286 12806
rect 3342 12772 3376 12806
rect 3432 12772 3466 12806
rect 3522 12772 3556 12806
rect 2982 12682 3016 12716
rect 3072 12682 3106 12716
rect 3162 12682 3196 12716
rect 3252 12682 3286 12716
rect 3342 12682 3376 12716
rect 3432 12682 3466 12716
rect 3522 12682 3556 12716
rect 2982 12592 3016 12626
rect 3072 12592 3106 12626
rect 3162 12592 3196 12626
rect 3252 12592 3286 12626
rect 3342 12592 3376 12626
rect 3432 12592 3466 12626
rect 3522 12592 3556 12626
rect 2982 12502 3016 12536
rect 3072 12502 3106 12536
rect 3162 12502 3196 12536
rect 3252 12502 3286 12536
rect 3342 12502 3376 12536
rect 3432 12502 3466 12536
rect 3522 12502 3556 12536
rect 4342 13042 4376 13076
rect 4432 13042 4466 13076
rect 4522 13042 4556 13076
rect 4612 13042 4646 13076
rect 4702 13042 4736 13076
rect 4792 13042 4826 13076
rect 4882 13042 4916 13076
rect 4342 12952 4376 12986
rect 4432 12952 4466 12986
rect 4522 12952 4556 12986
rect 4612 12952 4646 12986
rect 4702 12952 4736 12986
rect 4792 12952 4826 12986
rect 4882 12952 4916 12986
rect 4342 12862 4376 12896
rect 4432 12862 4466 12896
rect 4522 12862 4556 12896
rect 4612 12862 4646 12896
rect 4702 12862 4736 12896
rect 4792 12862 4826 12896
rect 4882 12862 4916 12896
rect 4342 12772 4376 12806
rect 4432 12772 4466 12806
rect 4522 12772 4556 12806
rect 4612 12772 4646 12806
rect 4702 12772 4736 12806
rect 4792 12772 4826 12806
rect 4882 12772 4916 12806
rect 4342 12682 4376 12716
rect 4432 12682 4466 12716
rect 4522 12682 4556 12716
rect 4612 12682 4646 12716
rect 4702 12682 4736 12716
rect 4792 12682 4826 12716
rect 4882 12682 4916 12716
rect 4342 12592 4376 12626
rect 4432 12592 4466 12626
rect 4522 12592 4556 12626
rect 4612 12592 4646 12626
rect 4702 12592 4736 12626
rect 4792 12592 4826 12626
rect 4882 12592 4916 12626
rect 4342 12502 4376 12536
rect 4432 12502 4466 12536
rect 4522 12502 4556 12536
rect 4612 12502 4646 12536
rect 4702 12502 4736 12536
rect 4792 12502 4826 12536
rect 4882 12502 4916 12536
rect 1622 11682 1656 11716
rect 1712 11682 1746 11716
rect 1802 11682 1836 11716
rect 1892 11682 1926 11716
rect 1982 11682 2016 11716
rect 2072 11682 2106 11716
rect 2162 11682 2196 11716
rect 1622 11592 1656 11626
rect 1712 11592 1746 11626
rect 1802 11592 1836 11626
rect 1892 11592 1926 11626
rect 1982 11592 2016 11626
rect 2072 11592 2106 11626
rect 2162 11592 2196 11626
rect 1622 11502 1656 11536
rect 1712 11502 1746 11536
rect 1802 11502 1836 11536
rect 1892 11502 1926 11536
rect 1982 11502 2016 11536
rect 2072 11502 2106 11536
rect 2162 11502 2196 11536
rect 1622 11412 1656 11446
rect 1712 11412 1746 11446
rect 1802 11412 1836 11446
rect 1892 11412 1926 11446
rect 1982 11412 2016 11446
rect 2072 11412 2106 11446
rect 2162 11412 2196 11446
rect 1622 11322 1656 11356
rect 1712 11322 1746 11356
rect 1802 11322 1836 11356
rect 1892 11322 1926 11356
rect 1982 11322 2016 11356
rect 2072 11322 2106 11356
rect 2162 11322 2196 11356
rect 1622 11232 1656 11266
rect 1712 11232 1746 11266
rect 1802 11232 1836 11266
rect 1892 11232 1926 11266
rect 1982 11232 2016 11266
rect 2072 11232 2106 11266
rect 2162 11232 2196 11266
rect 1622 11142 1656 11176
rect 1712 11142 1746 11176
rect 1802 11142 1836 11176
rect 1892 11142 1926 11176
rect 1982 11142 2016 11176
rect 2072 11142 2106 11176
rect 2162 11142 2196 11176
rect 2982 11682 3016 11716
rect 3072 11682 3106 11716
rect 3162 11682 3196 11716
rect 3252 11682 3286 11716
rect 3342 11682 3376 11716
rect 3432 11682 3466 11716
rect 3522 11682 3556 11716
rect 2982 11592 3016 11626
rect 3072 11592 3106 11626
rect 3162 11592 3196 11626
rect 3252 11592 3286 11626
rect 3342 11592 3376 11626
rect 3432 11592 3466 11626
rect 3522 11592 3556 11626
rect 2982 11502 3016 11536
rect 3072 11502 3106 11536
rect 3162 11502 3196 11536
rect 3252 11502 3286 11536
rect 3342 11502 3376 11536
rect 3432 11502 3466 11536
rect 3522 11502 3556 11536
rect 2982 11412 3016 11446
rect 3072 11412 3106 11446
rect 3162 11412 3196 11446
rect 3252 11412 3286 11446
rect 3342 11412 3376 11446
rect 3432 11412 3466 11446
rect 3522 11412 3556 11446
rect 2982 11322 3016 11356
rect 3072 11322 3106 11356
rect 3162 11322 3196 11356
rect 3252 11322 3286 11356
rect 3342 11322 3376 11356
rect 3432 11322 3466 11356
rect 3522 11322 3556 11356
rect 2982 11232 3016 11266
rect 3072 11232 3106 11266
rect 3162 11232 3196 11266
rect 3252 11232 3286 11266
rect 3342 11232 3376 11266
rect 3432 11232 3466 11266
rect 3522 11232 3556 11266
rect 2982 11142 3016 11176
rect 3072 11142 3106 11176
rect 3162 11142 3196 11176
rect 3252 11142 3286 11176
rect 3342 11142 3376 11176
rect 3432 11142 3466 11176
rect 3522 11142 3556 11176
rect 4342 11682 4376 11716
rect 4432 11682 4466 11716
rect 4522 11682 4556 11716
rect 4612 11682 4646 11716
rect 4702 11682 4736 11716
rect 4792 11682 4826 11716
rect 4882 11682 4916 11716
rect 4342 11592 4376 11626
rect 4432 11592 4466 11626
rect 4522 11592 4556 11626
rect 4612 11592 4646 11626
rect 4702 11592 4736 11626
rect 4792 11592 4826 11626
rect 4882 11592 4916 11626
rect 4342 11502 4376 11536
rect 4432 11502 4466 11536
rect 4522 11502 4556 11536
rect 4612 11502 4646 11536
rect 4702 11502 4736 11536
rect 4792 11502 4826 11536
rect 4882 11502 4916 11536
rect 4342 11412 4376 11446
rect 4432 11412 4466 11446
rect 4522 11412 4556 11446
rect 4612 11412 4646 11446
rect 4702 11412 4736 11446
rect 4792 11412 4826 11446
rect 4882 11412 4916 11446
rect 4342 11322 4376 11356
rect 4432 11322 4466 11356
rect 4522 11322 4556 11356
rect 4612 11322 4646 11356
rect 4702 11322 4736 11356
rect 4792 11322 4826 11356
rect 4882 11322 4916 11356
rect 4342 11232 4376 11266
rect 4432 11232 4466 11266
rect 4522 11232 4556 11266
rect 4612 11232 4646 11266
rect 4702 11232 4736 11266
rect 4792 11232 4826 11266
rect 4882 11232 4916 11266
rect 4342 11142 4376 11176
rect 4432 11142 4466 11176
rect 4522 11142 4556 11176
rect 4612 11142 4646 11176
rect 4702 11142 4736 11176
rect 4792 11142 4826 11176
rect 4882 11142 4916 11176
rect 530 7760 570 7800
rect 530 7660 570 7700
rect 650 7760 690 7800
rect 650 7660 690 7700
rect 770 7760 810 7800
rect 770 7660 810 7700
rect 890 7760 930 7800
rect 890 7660 930 7700
rect 1010 7760 1050 7800
rect 1010 7660 1050 7700
rect 1130 7760 1170 7800
rect 1130 7660 1170 7700
rect 1250 7760 1290 7800
rect 1250 7660 1290 7700
rect 1370 7760 1410 7800
rect 1370 7660 1410 7700
rect 1490 7760 1530 7800
rect 1490 7660 1530 7700
rect 1610 7760 1650 7800
rect 1610 7660 1650 7700
rect 1730 7760 1770 7800
rect 1730 7660 1770 7700
rect 1850 7760 1890 7800
rect 1850 7660 1890 7700
rect 1970 7760 2010 7800
rect 1970 7660 2010 7700
rect 2090 7760 2130 7800
rect 2090 7660 2130 7700
rect 2210 7760 2250 7800
rect 2210 7660 2250 7700
rect 2330 7760 2370 7800
rect 2330 7660 2370 7700
rect 2450 7760 2490 7800
rect 2450 7660 2490 7700
rect 2570 7760 2610 7800
rect 2570 7660 2610 7700
rect 2690 7760 2730 7800
rect 2690 7660 2730 7700
rect 2810 7760 2850 7800
rect 2810 7660 2850 7700
rect 2930 7760 2970 7800
rect 2930 7660 2970 7700
rect 3570 7760 3610 7800
rect 3570 7660 3610 7700
rect 3690 7760 3730 7800
rect 3690 7660 3730 7700
rect 3810 7760 3850 7800
rect 3810 7660 3850 7700
rect 3930 7760 3970 7800
rect 3930 7660 3970 7700
rect 4050 7760 4090 7800
rect 4050 7660 4090 7700
rect 4170 7760 4210 7800
rect 4170 7660 4210 7700
rect 4290 7760 4330 7800
rect 4290 7660 4330 7700
rect 4410 7760 4450 7800
rect 4410 7660 4450 7700
rect 4530 7760 4570 7800
rect 4530 7660 4570 7700
rect 4650 7760 4690 7800
rect 4650 7660 4690 7700
rect 4770 7760 4810 7800
rect 4770 7660 4810 7700
rect 4890 7760 4930 7800
rect 4890 7660 4930 7700
rect 5010 7760 5050 7800
rect 5010 7660 5050 7700
rect 5130 7760 5170 7800
rect 5130 7660 5170 7700
rect 5250 7760 5290 7800
rect 5250 7660 5290 7700
rect 5370 7760 5410 7800
rect 5370 7660 5410 7700
rect 5490 7760 5530 7800
rect 5490 7660 5530 7700
rect 5610 7760 5650 7800
rect 5610 7660 5650 7700
rect 5730 7760 5770 7800
rect 5730 7660 5770 7700
rect 5850 7760 5890 7800
rect 5850 7660 5890 7700
rect 5970 7760 6010 7800
rect 5970 7660 6010 7700
rect 8280 7280 8320 7320
rect 8280 7180 8320 7220
rect 8410 7280 8450 7320
rect 8410 7180 8450 7220
rect 8540 7280 8580 7320
rect 8540 7180 8580 7220
rect 8670 7280 8710 7320
rect 8670 7180 8710 7220
rect 8800 7280 8840 7320
rect 8800 7180 8840 7220
rect 8930 7280 8970 7320
rect 8930 7180 8970 7220
rect 9060 7280 9100 7320
rect 9060 7180 9100 7220
rect 9420 7280 9460 7320
rect 9420 7180 9460 7220
rect 9550 7280 9590 7320
rect 9550 7180 9590 7220
rect 9680 7280 9720 7320
rect 9680 7180 9720 7220
rect 9810 7280 9850 7320
rect 9810 7180 9850 7220
rect 9940 7280 9980 7320
rect 9940 7180 9980 7220
rect 10070 7280 10110 7320
rect 10070 7180 10110 7220
rect 10200 7280 10240 7320
rect 10200 7180 10240 7220
rect 10560 7280 10600 7320
rect 10560 7180 10600 7220
rect 10690 7280 10730 7320
rect 10690 7180 10730 7220
rect 10820 7280 10860 7320
rect 10820 7180 10860 7220
rect 10950 7280 10990 7320
rect 10950 7180 10990 7220
rect 11080 7280 11120 7320
rect 11080 7180 11120 7220
rect 11210 7280 11250 7320
rect 11210 7180 11250 7220
rect 11340 7280 11380 7320
rect 11340 7180 11380 7220
rect 1630 6600 1670 6640
rect 1630 6500 1670 6540
rect 1630 6400 1670 6440
rect 1630 6300 1670 6340
rect 1630 6200 1670 6240
rect 1630 6100 1670 6140
rect 1810 6600 1850 6640
rect 1810 6500 1850 6540
rect 1810 6400 1850 6440
rect 1810 6300 1850 6340
rect 1810 6200 1850 6240
rect 1810 6100 1850 6140
rect 1990 6600 2030 6640
rect 1990 6500 2030 6540
rect 1990 6400 2030 6440
rect 1990 6300 2030 6340
rect 1990 6200 2030 6240
rect 1990 6100 2030 6140
rect 2170 6600 2210 6640
rect 2170 6500 2210 6540
rect 2170 6400 2210 6440
rect 2170 6300 2210 6340
rect 2170 6200 2210 6240
rect 2170 6100 2210 6140
rect 2350 6600 2390 6640
rect 2350 6500 2390 6540
rect 2350 6400 2390 6440
rect 2350 6300 2390 6340
rect 2350 6200 2390 6240
rect 2350 6100 2390 6140
rect 2530 6600 2570 6640
rect 2530 6500 2570 6540
rect 2530 6400 2570 6440
rect 2530 6300 2570 6340
rect 2530 6200 2570 6240
rect 2530 6100 2570 6140
rect 2710 6600 2750 6640
rect 2710 6500 2750 6540
rect 2710 6400 2750 6440
rect 2710 6300 2750 6340
rect 2710 6200 2750 6240
rect 2710 6100 2750 6140
rect 2890 6600 2930 6640
rect 2890 6500 2930 6540
rect 2890 6400 2930 6440
rect 2890 6300 2930 6340
rect 2890 6200 2930 6240
rect 2890 6100 2930 6140
rect 3070 6600 3110 6640
rect 3070 6500 3110 6540
rect 3070 6400 3110 6440
rect 3070 6300 3110 6340
rect 3070 6200 3110 6240
rect 3070 6100 3110 6140
rect 3250 6600 3290 6640
rect 3250 6500 3290 6540
rect 3250 6400 3290 6440
rect 3250 6300 3290 6340
rect 3250 6200 3290 6240
rect 3250 6100 3290 6140
rect 3430 6600 3470 6640
rect 3430 6500 3470 6540
rect 3430 6400 3470 6440
rect 3430 6300 3470 6340
rect 3430 6200 3470 6240
rect 3430 6100 3470 6140
rect 3610 6600 3650 6640
rect 3610 6500 3650 6540
rect 3610 6400 3650 6440
rect 3610 6300 3650 6340
rect 3610 6200 3650 6240
rect 3610 6100 3650 6140
rect 3790 6600 3830 6640
rect 3790 6500 3830 6540
rect 3790 6400 3830 6440
rect 3790 6300 3830 6340
rect 3790 6200 3830 6240
rect 3790 6100 3830 6140
rect 3970 6600 4010 6640
rect 3970 6500 4010 6540
rect 3970 6400 4010 6440
rect 3970 6300 4010 6340
rect 3970 6200 4010 6240
rect 3970 6100 4010 6140
rect 4150 6600 4190 6640
rect 4150 6500 4190 6540
rect 4150 6400 4190 6440
rect 4150 6300 4190 6340
rect 4150 6200 4190 6240
rect 4150 6100 4190 6140
rect 4330 6600 4370 6640
rect 4330 6500 4370 6540
rect 4330 6400 4370 6440
rect 4330 6300 4370 6340
rect 4330 6200 4370 6240
rect 4330 6100 4370 6140
rect 4510 6600 4550 6640
rect 4510 6500 4550 6540
rect 4510 6400 4550 6440
rect 4510 6300 4550 6340
rect 4510 6200 4550 6240
rect 4510 6100 4550 6140
rect 4690 6600 4730 6640
rect 4690 6500 4730 6540
rect 4690 6400 4730 6440
rect 4690 6300 4730 6340
rect 4690 6200 4730 6240
rect 4690 6100 4730 6140
rect 4870 6600 4910 6640
rect 8350 6630 8390 6670
rect 4870 6500 4910 6540
rect 8350 6530 8390 6570
rect 4870 6400 4910 6440
rect 4870 6300 4910 6340
rect 5500 6400 5540 6440
rect 5500 6300 5540 6340
rect 5610 6400 5650 6440
rect 5610 6300 5650 6340
rect 5720 6400 5760 6440
rect 5720 6300 5760 6340
rect 5830 6400 5870 6440
rect 5830 6300 5870 6340
rect 5940 6400 5980 6440
rect 5940 6300 5980 6340
rect 8350 6430 8390 6470
rect 8350 6330 8390 6370
rect 4870 6200 4910 6240
rect 8350 6230 8390 6270
rect 8550 6630 8590 6670
rect 8550 6530 8590 6570
rect 8550 6430 8590 6470
rect 8550 6330 8590 6370
rect 8550 6230 8590 6270
rect 8750 6630 8790 6670
rect 8750 6530 8790 6570
rect 8750 6430 8790 6470
rect 8750 6330 8790 6370
rect 8750 6230 8790 6270
rect 8950 6630 8990 6670
rect 8950 6530 8990 6570
rect 8950 6430 8990 6470
rect 8950 6330 8990 6370
rect 8950 6230 8990 6270
rect 9150 6630 9190 6670
rect 9150 6530 9190 6570
rect 9150 6430 9190 6470
rect 9150 6330 9190 6370
rect 9150 6230 9190 6270
rect 9350 6630 9390 6670
rect 9350 6530 9390 6570
rect 9350 6430 9390 6470
rect 9350 6330 9390 6370
rect 9350 6230 9390 6270
rect 9550 6630 9590 6670
rect 9550 6530 9590 6570
rect 9550 6430 9590 6470
rect 9550 6330 9590 6370
rect 9550 6230 9590 6270
rect 9750 6630 9790 6670
rect 9750 6530 9790 6570
rect 9750 6430 9790 6470
rect 9750 6330 9790 6370
rect 9750 6230 9790 6270
rect 9950 6630 9990 6670
rect 9950 6530 9990 6570
rect 9950 6430 9990 6470
rect 9950 6330 9990 6370
rect 9950 6230 9990 6270
rect 10150 6630 10190 6670
rect 10150 6530 10190 6570
rect 10150 6430 10190 6470
rect 10150 6330 10190 6370
rect 10150 6230 10190 6270
rect 10350 6630 10390 6670
rect 10350 6530 10390 6570
rect 10350 6430 10390 6470
rect 10350 6330 10390 6370
rect 10350 6230 10390 6270
rect 4870 6100 4910 6140
rect 1640 5600 1680 5640
rect 1640 5500 1680 5540
rect 1750 5600 1790 5640
rect 1750 5500 1790 5540
rect 1860 5600 1900 5640
rect 1860 5500 1900 5540
rect 1970 5600 2010 5640
rect 1970 5500 2010 5540
rect 2080 5600 2120 5640
rect 2080 5500 2120 5540
rect 2190 5600 2230 5640
rect 2190 5500 2230 5540
rect 2300 5600 2340 5640
rect 2300 5500 2340 5540
rect 2410 5600 2450 5640
rect 2410 5500 2450 5540
rect 2520 5600 2560 5640
rect 2520 5500 2560 5540
rect 2630 5600 2670 5640
rect 2630 5500 2670 5540
rect 2740 5600 2780 5640
rect 2740 5500 2780 5540
rect 2850 5600 2890 5640
rect 2850 5500 2890 5540
rect 2960 5600 3000 5640
rect 2960 5500 3000 5540
rect 3540 5600 3580 5640
rect 3540 5500 3580 5540
rect 3650 5600 3690 5640
rect 3650 5500 3690 5540
rect 3760 5600 3800 5640
rect 3760 5500 3800 5540
rect 3870 5600 3910 5640
rect 3870 5500 3910 5540
rect 3980 5600 4020 5640
rect 3980 5500 4020 5540
rect 4090 5600 4130 5640
rect 4090 5500 4130 5540
rect 4200 5600 4240 5640
rect 4200 5500 4240 5540
rect 4310 5600 4350 5640
rect 4310 5500 4350 5540
rect 4420 5600 4460 5640
rect 4420 5500 4460 5540
rect 4530 5600 4570 5640
rect 4530 5500 4570 5540
rect 4640 5600 4680 5640
rect 4640 5500 4680 5540
rect 4750 5600 4790 5640
rect 4750 5500 4790 5540
rect 4860 5600 4900 5640
rect 4860 5500 4900 5540
rect 2160 4240 2200 4280
rect 2160 4140 2200 4180
rect 2160 4040 2200 4080
rect 2160 3940 2200 3980
rect 2270 4240 2310 4280
rect 2270 4140 2310 4180
rect 2270 4040 2310 4080
rect 2270 3940 2310 3980
rect 2380 4240 2420 4280
rect 2380 4140 2420 4180
rect 2380 4040 2420 4080
rect 2380 3940 2420 3980
rect 2680 4240 2720 4280
rect 2680 4140 2720 4180
rect 2680 4040 2720 4080
rect 2680 3940 2720 3980
rect 2790 4240 2830 4280
rect 2790 4140 2830 4180
rect 2790 4040 2830 4080
rect 2790 3940 2830 3980
rect 2900 4240 2940 4280
rect 3060 4240 3100 4280
rect 2900 4140 2940 4180
rect 3060 4140 3100 4180
rect 2900 4040 2940 4080
rect 3060 4040 3100 4080
rect 2900 3940 2940 3980
rect 3060 3940 3100 3980
rect 3170 4240 3210 4280
rect 3170 4140 3210 4180
rect 3170 4040 3210 4080
rect 3170 3940 3210 3980
rect 3280 4240 3320 4280
rect 3280 4140 3320 4180
rect 3280 4040 3320 4080
rect 3280 3940 3320 3980
rect 3580 4240 3620 4280
rect 3580 4140 3620 4180
rect 3580 4040 3620 4080
rect 3580 3940 3620 3980
rect 3690 4240 3730 4280
rect 3690 4140 3730 4180
rect 3690 4040 3730 4080
rect 3690 3940 3730 3980
rect 3800 4240 3840 4280
rect 3800 4140 3840 4180
rect 3800 4040 3840 4080
rect 3800 3940 3840 3980
rect 4100 4240 4140 4280
rect 4100 4140 4140 4180
rect 4100 4040 4140 4080
rect 4100 3940 4140 3980
rect 4210 4240 4250 4280
rect 4210 4140 4250 4180
rect 4210 4040 4250 4080
rect 4210 3940 4250 3980
rect 4320 4240 4360 4280
rect 4320 4140 4360 4180
rect 4320 4040 4360 4080
rect 4320 3940 4360 3980
rect 4540 4240 4580 4280
rect 4540 4140 4580 4180
rect 4540 4040 4580 4080
rect 4540 3940 4580 3980
rect 4650 4240 4690 4280
rect 4650 4140 4690 4180
rect 4650 4040 4690 4080
rect 4650 3940 4690 3980
rect 4870 4240 4910 4280
rect 4870 4140 4910 4180
rect 4870 4040 4910 4080
rect 4870 3940 4910 3980
rect 4980 4240 5020 4280
rect 4980 4140 5020 4180
rect 4980 4040 5020 4080
rect 4980 3940 5020 3980
rect 5300 4240 5340 4280
rect 5300 4140 5340 4180
rect 5300 4040 5340 4080
rect 5300 3940 5340 3980
rect 5430 4240 5470 4280
rect 5430 4140 5470 4180
rect 5430 4040 5470 4080
rect 5430 3940 5470 3980
rect 5690 4240 5730 4280
rect 5690 4140 5730 4180
rect 5690 4040 5730 4080
rect 5690 3940 5730 3980
rect 5820 4240 5860 4280
rect 5820 4140 5860 4180
rect 5820 4040 5860 4080
rect 5820 3940 5860 3980
rect 6080 4240 6120 4280
rect 6080 4140 6120 4180
rect 6080 4040 6120 4080
rect 6080 3940 6120 3980
rect 6210 4240 6250 4280
rect 6210 4140 6250 4180
rect 6210 4040 6250 4080
rect 6210 3940 6250 3980
rect 6370 4240 6410 4280
rect 6370 4140 6410 4180
rect 6370 4040 6410 4080
rect 6370 3940 6410 3980
rect 6500 4240 6540 4280
rect 6500 4140 6540 4180
rect 6500 4040 6540 4080
rect 6500 3940 6540 3980
rect 6760 4240 6800 4280
rect 6760 4140 6800 4180
rect 6760 4040 6800 4080
rect 6760 3940 6800 3980
rect 6890 4240 6930 4280
rect 6890 4140 6930 4180
rect 6890 4040 6930 4080
rect 6890 3940 6930 3980
rect 8170 4290 8210 4330
rect 8170 4190 8210 4230
rect 8170 4090 8210 4130
rect 8170 3990 8210 4030
rect 8390 4290 8430 4330
rect 8390 4190 8430 4230
rect 8390 4090 8430 4130
rect 8390 3990 8430 4030
rect 8610 4290 8650 4330
rect 8610 4190 8650 4230
rect 8610 4090 8650 4130
rect 8610 3990 8650 4030
rect 8830 4290 8870 4330
rect 8830 4190 8870 4230
rect 8830 4090 8870 4130
rect 8830 3990 8870 4030
rect 9050 4290 9090 4330
rect 9050 4190 9090 4230
rect 9050 4090 9090 4130
rect 9050 3990 9090 4030
rect 9270 4290 9310 4330
rect 9270 4190 9310 4230
rect 9270 4090 9310 4130
rect 9270 3990 9310 4030
rect 9490 4290 9530 4330
rect 9690 4290 9730 4330
rect 9490 4190 9530 4230
rect 9690 4190 9730 4230
rect 9490 4090 9530 4130
rect 9690 4090 9730 4130
rect 9490 3990 9530 4030
rect 9690 3990 9730 4030
rect 9910 4290 9950 4330
rect 9910 4190 9950 4230
rect 9910 4090 9950 4130
rect 9910 3990 9950 4030
rect 10130 4290 10170 4330
rect 10130 4190 10170 4230
rect 10130 4090 10170 4130
rect 10130 3990 10170 4030
rect 10350 4290 10390 4330
rect 10350 4190 10390 4230
rect 10350 4090 10390 4130
rect 10350 3990 10390 4030
rect 10570 4290 10610 4330
rect 10570 4190 10610 4230
rect 10570 4090 10610 4130
rect 10570 3990 10610 4030
rect 10790 4290 10830 4330
rect 10790 4190 10830 4230
rect 10790 4090 10830 4130
rect 10790 3990 10830 4030
rect 11010 4290 11050 4330
rect 11010 4190 11050 4230
rect 11010 4090 11050 4130
rect 11010 3990 11050 4030
rect 2160 3480 2200 3520
rect 2160 3380 2200 3420
rect 2160 3280 2200 3320
rect 2160 3180 2200 3220
rect 2270 3480 2310 3520
rect 2270 3380 2310 3420
rect 2270 3280 2310 3320
rect 2270 3180 2310 3220
rect 2380 3480 2420 3520
rect 2380 3380 2420 3420
rect 2380 3280 2420 3320
rect 2380 3180 2420 3220
rect 2680 3480 2720 3520
rect 2680 3380 2720 3420
rect 2680 3280 2720 3320
rect 2680 3180 2720 3220
rect 2790 3480 2830 3520
rect 2790 3380 2830 3420
rect 2790 3280 2830 3320
rect 2790 3180 2830 3220
rect 2900 3480 2940 3520
rect 3060 3480 3100 3520
rect 2900 3380 2940 3420
rect 3060 3380 3100 3420
rect 2900 3280 2940 3320
rect 3060 3280 3100 3320
rect 2900 3180 2940 3220
rect 3060 3180 3100 3220
rect 3170 3480 3210 3520
rect 3170 3380 3210 3420
rect 3170 3280 3210 3320
rect 3170 3180 3210 3220
rect 3280 3480 3320 3520
rect 3280 3380 3320 3420
rect 3280 3280 3320 3320
rect 3280 3180 3320 3220
rect 3580 3480 3620 3520
rect 3580 3380 3620 3420
rect 3580 3280 3620 3320
rect 3580 3180 3620 3220
rect 3690 3480 3730 3520
rect 3690 3380 3730 3420
rect 3690 3280 3730 3320
rect 3690 3180 3730 3220
rect 3800 3480 3840 3520
rect 3800 3380 3840 3420
rect 3800 3280 3840 3320
rect 3800 3180 3840 3220
rect 4090 3480 4130 3520
rect 4090 3380 4130 3420
rect 4090 3280 4130 3320
rect 4090 3180 4130 3220
rect 4200 3480 4240 3520
rect 4200 3380 4240 3420
rect 4200 3280 4240 3320
rect 4200 3180 4240 3220
rect 4420 3480 4460 3520
rect 4420 3380 4460 3420
rect 4420 3280 4460 3320
rect 4420 3180 4460 3220
rect 4530 3480 4570 3520
rect 4530 3380 4570 3420
rect 4530 3280 4570 3320
rect 4530 3180 4570 3220
rect 4750 3480 4790 3520
rect 4750 3380 4790 3420
rect 4750 3280 4790 3320
rect 4750 3180 4790 3220
rect 4860 3480 4900 3520
rect 4860 3380 4900 3420
rect 4860 3280 4900 3320
rect 4860 3180 4900 3220
rect 5300 3480 5340 3520
rect 5300 3380 5340 3420
rect 5300 3280 5340 3320
rect 5300 3180 5340 3220
rect 5430 3480 5470 3520
rect 5430 3380 5470 3420
rect 5430 3280 5470 3320
rect 5430 3180 5470 3220
rect 5690 3480 5730 3520
rect 5690 3380 5730 3420
rect 5690 3280 5730 3320
rect 5690 3180 5730 3220
rect 5820 3480 5860 3520
rect 5820 3380 5860 3420
rect 5820 3280 5860 3320
rect 5820 3180 5860 3220
rect 6080 3480 6120 3520
rect 6080 3380 6120 3420
rect 6080 3280 6120 3320
rect 6080 3180 6120 3220
rect 6210 3480 6250 3520
rect 6210 3380 6250 3420
rect 6210 3280 6250 3320
rect 6210 3180 6250 3220
rect 6370 3480 6410 3520
rect 6370 3380 6410 3420
rect 6370 3280 6410 3320
rect 6370 3180 6410 3220
rect 6500 3480 6540 3520
rect 6500 3380 6540 3420
rect 6500 3280 6540 3320
rect 6500 3180 6540 3220
rect 2010 1050 2050 1090
rect 2120 1050 2160 1090
rect 2430 1050 2470 1090
rect 2540 1050 2580 1090
rect 2650 1050 2690 1090
rect 3100 1050 3140 1090
rect 3210 1050 3250 1090
rect 3320 1050 3360 1090
rect 3540 1050 3580 1090
rect 3650 1050 3690 1090
rect 3760 1050 3800 1090
rect 3870 1050 3910 1090
rect 4380 1050 4420 1090
rect 4490 1050 4530 1090
rect 4800 1050 4840 1090
rect 4910 1050 4950 1090
rect 5020 1050 5060 1090
rect 5250 1050 5290 1090
rect 5360 1050 5400 1090
rect 5470 1050 5510 1090
rect 5610 1050 5650 1090
rect 5720 1050 5760 1090
rect 5830 1050 5870 1090
rect 6190 1050 6230 1090
rect 6300 1050 6340 1090
rect 6410 1050 6450 1090
rect 6630 1050 6670 1090
rect 6740 1050 6780 1090
rect 6850 1050 6890 1090
rect 12420 1150 12460 1190
rect 7250 1050 7290 1090
rect 7360 1050 7400 1090
rect 7590 1050 7630 1090
rect 7700 1050 7740 1090
rect 7810 1050 7850 1090
rect 7950 1050 7990 1090
rect 8060 1050 8100 1090
rect 8170 1050 8210 1090
rect 8550 1050 8590 1090
rect 8660 1050 8700 1090
rect 8890 1050 8930 1090
rect 9000 1050 9040 1090
rect 9110 1050 9150 1090
rect 9250 1050 9290 1090
rect 9360 1050 9400 1090
rect 9470 1050 9510 1090
rect 9850 1050 9890 1090
rect 9960 1050 10000 1090
rect 10190 1050 10230 1090
rect 10300 1050 10340 1090
rect 10410 1050 10450 1090
rect 10550 1050 10590 1090
rect 10660 1050 10700 1090
rect 10770 1050 10810 1090
rect 11150 1050 11190 1090
rect 11260 1050 11300 1090
rect 11490 1050 11530 1090
rect 11600 1050 11640 1090
rect 11710 1050 11750 1090
rect 11850 1050 11890 1090
rect 11960 1050 12000 1090
rect 12070 1050 12110 1090
rect 12420 1050 12460 1090
rect 12530 1150 12570 1190
rect 12530 1050 12570 1090
rect 13020 1150 13060 1190
rect 13020 1050 13060 1090
rect 13130 1150 13170 1190
rect 13130 1050 13170 1090
rect 13620 1150 13660 1190
rect 13620 1050 13660 1090
rect 13730 1150 13770 1190
rect 13730 1050 13770 1090
rect 12420 810 12460 850
rect 12420 710 12460 750
rect 12530 810 12570 850
rect 12530 710 12570 750
rect 13020 810 13060 850
rect 13020 710 13060 750
rect 13130 810 13170 850
rect 13130 710 13170 750
rect 13620 810 13660 850
rect 13620 710 13660 750
rect 13730 810 13770 850
rect 13730 710 13770 750
rect 12420 460 12460 500
rect 12420 360 12460 400
rect 12420 260 12460 300
rect 12420 160 12460 200
rect 12800 460 12840 500
rect 12800 360 12840 400
rect 12800 260 12840 300
rect 12800 160 12840 200
rect 13020 460 13060 500
rect 13020 360 13060 400
rect 13020 260 13060 300
rect 13020 160 13060 200
rect 13400 460 13440 500
rect 13400 360 13440 400
rect 13400 260 13440 300
rect 13400 160 13440 200
rect 13620 460 13660 500
rect 13620 360 13660 400
rect 13620 260 13660 300
rect 13620 160 13660 200
rect 14000 460 14040 500
rect 14160 460 14200 500
rect 14000 360 14040 400
rect 14160 360 14200 400
rect 14000 260 14040 300
rect 14160 260 14200 300
rect 14000 160 14040 200
rect 14160 160 14200 200
rect 14540 460 14580 500
rect 14540 360 14580 400
rect 14540 260 14580 300
rect 14540 160 14580 200
<< psubdiff >>
rect 3220 15080 3320 15110
rect 3220 15040 3250 15080
rect 3290 15040 3320 15080
rect 3220 15000 3320 15040
rect 3220 14960 3250 15000
rect 3290 14960 3320 15000
rect 3220 14920 3320 14960
rect 3220 14880 3250 14920
rect 3290 14880 3320 14920
rect 3220 14850 3320 14880
rect 1266 14762 2554 14794
rect 1266 14728 1400 14762
rect 1434 14728 1490 14762
rect 1524 14728 1580 14762
rect 1614 14728 1670 14762
rect 1704 14728 1760 14762
rect 1794 14728 1850 14762
rect 1884 14728 1940 14762
rect 1974 14728 2030 14762
rect 2064 14728 2120 14762
rect 2154 14728 2210 14762
rect 2244 14728 2300 14762
rect 2334 14728 2390 14762
rect 2424 14728 2554 14762
rect 1266 14693 2554 14728
rect 1266 14678 1367 14693
rect 1266 14644 1299 14678
rect 1333 14644 1367 14678
rect 1266 14588 1367 14644
rect 2453 14678 2554 14693
rect 2453 14644 2486 14678
rect 2520 14644 2554 14678
rect 1266 14554 1299 14588
rect 1333 14554 1367 14588
rect 1266 14498 1367 14554
rect 1266 14464 1299 14498
rect 1333 14464 1367 14498
rect 1266 14408 1367 14464
rect 1266 14374 1299 14408
rect 1333 14374 1367 14408
rect 1266 14318 1367 14374
rect 1266 14284 1299 14318
rect 1333 14284 1367 14318
rect 1266 14228 1367 14284
rect 1266 14194 1299 14228
rect 1333 14194 1367 14228
rect 1266 14138 1367 14194
rect 1266 14104 1299 14138
rect 1333 14104 1367 14138
rect 1266 14048 1367 14104
rect 1266 14014 1299 14048
rect 1333 14014 1367 14048
rect 1266 13958 1367 14014
rect 1266 13924 1299 13958
rect 1333 13924 1367 13958
rect 1266 13868 1367 13924
rect 1266 13834 1299 13868
rect 1333 13834 1367 13868
rect 1266 13778 1367 13834
rect 1266 13744 1299 13778
rect 1333 13744 1367 13778
rect 1266 13688 1367 13744
rect 1266 13654 1299 13688
rect 1333 13654 1367 13688
rect 2453 14588 2554 14644
rect 2453 14554 2486 14588
rect 2520 14554 2554 14588
rect 2453 14498 2554 14554
rect 2453 14464 2486 14498
rect 2520 14464 2554 14498
rect 2453 14408 2554 14464
rect 2453 14374 2486 14408
rect 2520 14374 2554 14408
rect 2453 14318 2554 14374
rect 2453 14284 2486 14318
rect 2520 14284 2554 14318
rect 2453 14228 2554 14284
rect 2453 14194 2486 14228
rect 2520 14194 2554 14228
rect 2453 14138 2554 14194
rect 2453 14104 2486 14138
rect 2520 14104 2554 14138
rect 2453 14048 2554 14104
rect 2453 14014 2486 14048
rect 2520 14014 2554 14048
rect 2453 13958 2554 14014
rect 2453 13924 2486 13958
rect 2520 13924 2554 13958
rect 2453 13868 2554 13924
rect 2453 13834 2486 13868
rect 2520 13834 2554 13868
rect 2453 13778 2554 13834
rect 2453 13744 2486 13778
rect 2520 13744 2554 13778
rect 2453 13688 2554 13744
rect 1266 13607 1367 13654
rect 2453 13654 2486 13688
rect 2520 13654 2554 13688
rect 2453 13607 2554 13654
rect 1266 13598 2554 13607
rect 1266 13564 1299 13598
rect 1333 13575 2486 13598
rect 1333 13564 1400 13575
rect 1266 13541 1400 13564
rect 1434 13541 1490 13575
rect 1524 13541 1580 13575
rect 1614 13541 1670 13575
rect 1704 13541 1760 13575
rect 1794 13541 1850 13575
rect 1884 13541 1940 13575
rect 1974 13541 2030 13575
rect 2064 13541 2120 13575
rect 2154 13541 2210 13575
rect 2244 13541 2300 13575
rect 2334 13541 2390 13575
rect 2424 13564 2486 13575
rect 2520 13564 2554 13598
rect 2424 13541 2554 13564
rect 1266 13506 2554 13541
rect 2626 14762 3914 14794
rect 2626 14728 2760 14762
rect 2794 14728 2850 14762
rect 2884 14728 2940 14762
rect 2974 14728 3030 14762
rect 3064 14728 3120 14762
rect 3154 14728 3210 14762
rect 3244 14728 3300 14762
rect 3334 14728 3390 14762
rect 3424 14728 3480 14762
rect 3514 14728 3570 14762
rect 3604 14728 3660 14762
rect 3694 14728 3750 14762
rect 3784 14728 3914 14762
rect 2626 14693 3914 14728
rect 2626 14678 2727 14693
rect 2626 14644 2659 14678
rect 2693 14644 2727 14678
rect 2626 14588 2727 14644
rect 3813 14678 3914 14693
rect 3813 14644 3846 14678
rect 3880 14644 3914 14678
rect 2626 14554 2659 14588
rect 2693 14554 2727 14588
rect 2626 14498 2727 14554
rect 2626 14464 2659 14498
rect 2693 14464 2727 14498
rect 2626 14408 2727 14464
rect 2626 14374 2659 14408
rect 2693 14374 2727 14408
rect 2626 14318 2727 14374
rect 2626 14284 2659 14318
rect 2693 14284 2727 14318
rect 2626 14228 2727 14284
rect 2626 14194 2659 14228
rect 2693 14194 2727 14228
rect 2626 14138 2727 14194
rect 2626 14104 2659 14138
rect 2693 14104 2727 14138
rect 2626 14048 2727 14104
rect 2626 14014 2659 14048
rect 2693 14014 2727 14048
rect 2626 13958 2727 14014
rect 2626 13924 2659 13958
rect 2693 13924 2727 13958
rect 2626 13868 2727 13924
rect 2626 13834 2659 13868
rect 2693 13834 2727 13868
rect 2626 13778 2727 13834
rect 2626 13744 2659 13778
rect 2693 13744 2727 13778
rect 2626 13688 2727 13744
rect 2626 13654 2659 13688
rect 2693 13654 2727 13688
rect 3813 14588 3914 14644
rect 3813 14554 3846 14588
rect 3880 14554 3914 14588
rect 3813 14498 3914 14554
rect 3813 14464 3846 14498
rect 3880 14464 3914 14498
rect 3813 14408 3914 14464
rect 3813 14374 3846 14408
rect 3880 14374 3914 14408
rect 3813 14318 3914 14374
rect 3813 14284 3846 14318
rect 3880 14284 3914 14318
rect 3813 14228 3914 14284
rect 3813 14194 3846 14228
rect 3880 14194 3914 14228
rect 3813 14138 3914 14194
rect 3813 14104 3846 14138
rect 3880 14104 3914 14138
rect 3813 14048 3914 14104
rect 3813 14014 3846 14048
rect 3880 14014 3914 14048
rect 3813 13958 3914 14014
rect 3813 13924 3846 13958
rect 3880 13924 3914 13958
rect 3813 13868 3914 13924
rect 3813 13834 3846 13868
rect 3880 13834 3914 13868
rect 3813 13778 3914 13834
rect 3813 13744 3846 13778
rect 3880 13744 3914 13778
rect 3813 13688 3914 13744
rect 2626 13607 2727 13654
rect 3813 13654 3846 13688
rect 3880 13654 3914 13688
rect 3813 13607 3914 13654
rect 2626 13598 3914 13607
rect 2626 13564 2659 13598
rect 2693 13575 3846 13598
rect 2693 13564 2760 13575
rect 2626 13541 2760 13564
rect 2794 13541 2850 13575
rect 2884 13541 2940 13575
rect 2974 13541 3030 13575
rect 3064 13541 3120 13575
rect 3154 13541 3210 13575
rect 3244 13541 3300 13575
rect 3334 13541 3390 13575
rect 3424 13541 3480 13575
rect 3514 13541 3570 13575
rect 3604 13541 3660 13575
rect 3694 13541 3750 13575
rect 3784 13564 3846 13575
rect 3880 13564 3914 13598
rect 3784 13541 3914 13564
rect 2626 13506 3914 13541
rect 3986 14762 5274 14794
rect 3986 14728 4120 14762
rect 4154 14728 4210 14762
rect 4244 14728 4300 14762
rect 4334 14728 4390 14762
rect 4424 14728 4480 14762
rect 4514 14728 4570 14762
rect 4604 14728 4660 14762
rect 4694 14728 4750 14762
rect 4784 14728 4840 14762
rect 4874 14728 4930 14762
rect 4964 14728 5020 14762
rect 5054 14728 5110 14762
rect 5144 14728 5274 14762
rect 3986 14693 5274 14728
rect 3986 14678 4087 14693
rect 3986 14644 4019 14678
rect 4053 14644 4087 14678
rect 3986 14588 4087 14644
rect 5173 14678 5274 14693
rect 5173 14644 5206 14678
rect 5240 14644 5274 14678
rect 3986 14554 4019 14588
rect 4053 14554 4087 14588
rect 3986 14498 4087 14554
rect 3986 14464 4019 14498
rect 4053 14464 4087 14498
rect 3986 14408 4087 14464
rect 3986 14374 4019 14408
rect 4053 14374 4087 14408
rect 3986 14318 4087 14374
rect 3986 14284 4019 14318
rect 4053 14284 4087 14318
rect 3986 14228 4087 14284
rect 3986 14194 4019 14228
rect 4053 14194 4087 14228
rect 3986 14138 4087 14194
rect 3986 14104 4019 14138
rect 4053 14104 4087 14138
rect 3986 14048 4087 14104
rect 3986 14014 4019 14048
rect 4053 14014 4087 14048
rect 3986 13958 4087 14014
rect 3986 13924 4019 13958
rect 4053 13924 4087 13958
rect 3986 13868 4087 13924
rect 3986 13834 4019 13868
rect 4053 13834 4087 13868
rect 3986 13778 4087 13834
rect 3986 13744 4019 13778
rect 4053 13744 4087 13778
rect 3986 13688 4087 13744
rect 3986 13654 4019 13688
rect 4053 13654 4087 13688
rect 5173 14588 5274 14644
rect 5173 14554 5206 14588
rect 5240 14554 5274 14588
rect 5173 14498 5274 14554
rect 5173 14464 5206 14498
rect 5240 14464 5274 14498
rect 5173 14408 5274 14464
rect 5173 14374 5206 14408
rect 5240 14374 5274 14408
rect 5173 14318 5274 14374
rect 5173 14284 5206 14318
rect 5240 14284 5274 14318
rect 5173 14228 5274 14284
rect 5173 14194 5206 14228
rect 5240 14194 5274 14228
rect 5173 14138 5274 14194
rect 5173 14104 5206 14138
rect 5240 14104 5274 14138
rect 5173 14048 5274 14104
rect 5173 14014 5206 14048
rect 5240 14014 5274 14048
rect 5173 13958 5274 14014
rect 5173 13924 5206 13958
rect 5240 13924 5274 13958
rect 5173 13868 5274 13924
rect 5173 13834 5206 13868
rect 5240 13834 5274 13868
rect 5173 13778 5274 13834
rect 5173 13744 5206 13778
rect 5240 13744 5274 13778
rect 5173 13688 5274 13744
rect 3986 13607 4087 13654
rect 5173 13654 5206 13688
rect 5240 13654 5274 13688
rect 5173 13607 5274 13654
rect 3986 13598 5274 13607
rect 3986 13564 4019 13598
rect 4053 13575 5206 13598
rect 4053 13564 4120 13575
rect 3986 13541 4120 13564
rect 4154 13541 4210 13575
rect 4244 13541 4300 13575
rect 4334 13541 4390 13575
rect 4424 13541 4480 13575
rect 4514 13541 4570 13575
rect 4604 13541 4660 13575
rect 4694 13541 4750 13575
rect 4784 13541 4840 13575
rect 4874 13541 4930 13575
rect 4964 13541 5020 13575
rect 5054 13541 5110 13575
rect 5144 13564 5206 13575
rect 5240 13564 5274 13598
rect 5144 13541 5274 13564
rect 3986 13506 5274 13541
rect 1266 13402 2554 13434
rect 1266 13368 1400 13402
rect 1434 13368 1490 13402
rect 1524 13368 1580 13402
rect 1614 13368 1670 13402
rect 1704 13368 1760 13402
rect 1794 13368 1850 13402
rect 1884 13368 1940 13402
rect 1974 13368 2030 13402
rect 2064 13368 2120 13402
rect 2154 13368 2210 13402
rect 2244 13368 2300 13402
rect 2334 13368 2390 13402
rect 2424 13368 2554 13402
rect 1266 13333 2554 13368
rect 1266 13318 1367 13333
rect 1266 13284 1299 13318
rect 1333 13284 1367 13318
rect 1266 13228 1367 13284
rect 2453 13318 2554 13333
rect 2453 13284 2486 13318
rect 2520 13284 2554 13318
rect 1266 13194 1299 13228
rect 1333 13194 1367 13228
rect 1266 13138 1367 13194
rect 1266 13104 1299 13138
rect 1333 13104 1367 13138
rect 1266 13048 1367 13104
rect 1266 13014 1299 13048
rect 1333 13014 1367 13048
rect 1266 12958 1367 13014
rect 1266 12924 1299 12958
rect 1333 12924 1367 12958
rect 1266 12868 1367 12924
rect 1266 12834 1299 12868
rect 1333 12834 1367 12868
rect 1266 12778 1367 12834
rect 1266 12744 1299 12778
rect 1333 12744 1367 12778
rect 1266 12688 1367 12744
rect 1266 12654 1299 12688
rect 1333 12654 1367 12688
rect 1266 12598 1367 12654
rect 1266 12564 1299 12598
rect 1333 12564 1367 12598
rect 1266 12508 1367 12564
rect 1266 12474 1299 12508
rect 1333 12474 1367 12508
rect 1266 12418 1367 12474
rect 1266 12384 1299 12418
rect 1333 12384 1367 12418
rect 1266 12328 1367 12384
rect 1266 12294 1299 12328
rect 1333 12294 1367 12328
rect 2453 13228 2554 13284
rect 2453 13194 2486 13228
rect 2520 13194 2554 13228
rect 2453 13138 2554 13194
rect 2453 13104 2486 13138
rect 2520 13104 2554 13138
rect 2453 13048 2554 13104
rect 2453 13014 2486 13048
rect 2520 13014 2554 13048
rect 2453 12958 2554 13014
rect 2453 12924 2486 12958
rect 2520 12924 2554 12958
rect 2453 12868 2554 12924
rect 2453 12834 2486 12868
rect 2520 12834 2554 12868
rect 2453 12778 2554 12834
rect 2453 12744 2486 12778
rect 2520 12744 2554 12778
rect 2453 12688 2554 12744
rect 2453 12654 2486 12688
rect 2520 12654 2554 12688
rect 2453 12598 2554 12654
rect 2453 12564 2486 12598
rect 2520 12564 2554 12598
rect 2453 12508 2554 12564
rect 2453 12474 2486 12508
rect 2520 12474 2554 12508
rect 2453 12418 2554 12474
rect 2453 12384 2486 12418
rect 2520 12384 2554 12418
rect 2453 12328 2554 12384
rect 1266 12247 1367 12294
rect 2453 12294 2486 12328
rect 2520 12294 2554 12328
rect 2453 12247 2554 12294
rect 1266 12238 2554 12247
rect 1266 12204 1299 12238
rect 1333 12215 2486 12238
rect 1333 12204 1400 12215
rect 1266 12181 1400 12204
rect 1434 12181 1490 12215
rect 1524 12181 1580 12215
rect 1614 12181 1670 12215
rect 1704 12181 1760 12215
rect 1794 12181 1850 12215
rect 1884 12181 1940 12215
rect 1974 12181 2030 12215
rect 2064 12181 2120 12215
rect 2154 12181 2210 12215
rect 2244 12181 2300 12215
rect 2334 12181 2390 12215
rect 2424 12204 2486 12215
rect 2520 12204 2554 12238
rect 2424 12181 2554 12204
rect 1266 12146 2554 12181
rect 2626 13402 3914 13434
rect 2626 13368 2760 13402
rect 2794 13368 2850 13402
rect 2884 13368 2940 13402
rect 2974 13368 3030 13402
rect 3064 13368 3120 13402
rect 3154 13368 3210 13402
rect 3244 13368 3300 13402
rect 3334 13368 3390 13402
rect 3424 13368 3480 13402
rect 3514 13368 3570 13402
rect 3604 13368 3660 13402
rect 3694 13368 3750 13402
rect 3784 13368 3914 13402
rect 2626 13333 3914 13368
rect 2626 13318 2727 13333
rect 2626 13284 2659 13318
rect 2693 13284 2727 13318
rect 2626 13228 2727 13284
rect 3813 13318 3914 13333
rect 3813 13284 3846 13318
rect 3880 13284 3914 13318
rect 2626 13194 2659 13228
rect 2693 13194 2727 13228
rect 2626 13138 2727 13194
rect 2626 13104 2659 13138
rect 2693 13104 2727 13138
rect 2626 13048 2727 13104
rect 2626 13014 2659 13048
rect 2693 13014 2727 13048
rect 2626 12958 2727 13014
rect 2626 12924 2659 12958
rect 2693 12924 2727 12958
rect 2626 12868 2727 12924
rect 2626 12834 2659 12868
rect 2693 12834 2727 12868
rect 2626 12778 2727 12834
rect 2626 12744 2659 12778
rect 2693 12744 2727 12778
rect 2626 12688 2727 12744
rect 2626 12654 2659 12688
rect 2693 12654 2727 12688
rect 2626 12598 2727 12654
rect 2626 12564 2659 12598
rect 2693 12564 2727 12598
rect 2626 12508 2727 12564
rect 2626 12474 2659 12508
rect 2693 12474 2727 12508
rect 2626 12418 2727 12474
rect 2626 12384 2659 12418
rect 2693 12384 2727 12418
rect 2626 12328 2727 12384
rect 2626 12294 2659 12328
rect 2693 12294 2727 12328
rect 3813 13228 3914 13284
rect 3813 13194 3846 13228
rect 3880 13194 3914 13228
rect 3813 13138 3914 13194
rect 3813 13104 3846 13138
rect 3880 13104 3914 13138
rect 3813 13048 3914 13104
rect 3813 13014 3846 13048
rect 3880 13014 3914 13048
rect 3813 12958 3914 13014
rect 3813 12924 3846 12958
rect 3880 12924 3914 12958
rect 3813 12868 3914 12924
rect 3813 12834 3846 12868
rect 3880 12834 3914 12868
rect 3813 12778 3914 12834
rect 3813 12744 3846 12778
rect 3880 12744 3914 12778
rect 3813 12688 3914 12744
rect 3813 12654 3846 12688
rect 3880 12654 3914 12688
rect 3813 12598 3914 12654
rect 3813 12564 3846 12598
rect 3880 12564 3914 12598
rect 3813 12508 3914 12564
rect 3813 12474 3846 12508
rect 3880 12474 3914 12508
rect 3813 12418 3914 12474
rect 3813 12384 3846 12418
rect 3880 12384 3914 12418
rect 3813 12328 3914 12384
rect 2626 12247 2727 12294
rect 3813 12294 3846 12328
rect 3880 12294 3914 12328
rect 3813 12247 3914 12294
rect 2626 12238 3914 12247
rect 2626 12204 2659 12238
rect 2693 12215 3846 12238
rect 2693 12204 2760 12215
rect 2626 12181 2760 12204
rect 2794 12181 2850 12215
rect 2884 12181 2940 12215
rect 2974 12181 3030 12215
rect 3064 12181 3120 12215
rect 3154 12181 3210 12215
rect 3244 12181 3300 12215
rect 3334 12181 3390 12215
rect 3424 12181 3480 12215
rect 3514 12181 3570 12215
rect 3604 12181 3660 12215
rect 3694 12181 3750 12215
rect 3784 12204 3846 12215
rect 3880 12204 3914 12238
rect 3784 12181 3914 12204
rect 2626 12146 3914 12181
rect 3986 13402 5274 13434
rect 3986 13368 4120 13402
rect 4154 13368 4210 13402
rect 4244 13368 4300 13402
rect 4334 13368 4390 13402
rect 4424 13368 4480 13402
rect 4514 13368 4570 13402
rect 4604 13368 4660 13402
rect 4694 13368 4750 13402
rect 4784 13368 4840 13402
rect 4874 13368 4930 13402
rect 4964 13368 5020 13402
rect 5054 13368 5110 13402
rect 5144 13368 5274 13402
rect 3986 13333 5274 13368
rect 3986 13318 4087 13333
rect 3986 13284 4019 13318
rect 4053 13284 4087 13318
rect 3986 13228 4087 13284
rect 5173 13318 5274 13333
rect 5173 13284 5206 13318
rect 5240 13284 5274 13318
rect 3986 13194 4019 13228
rect 4053 13194 4087 13228
rect 3986 13138 4087 13194
rect 3986 13104 4019 13138
rect 4053 13104 4087 13138
rect 3986 13048 4087 13104
rect 3986 13014 4019 13048
rect 4053 13014 4087 13048
rect 3986 12958 4087 13014
rect 3986 12924 4019 12958
rect 4053 12924 4087 12958
rect 3986 12868 4087 12924
rect 3986 12834 4019 12868
rect 4053 12834 4087 12868
rect 3986 12778 4087 12834
rect 3986 12744 4019 12778
rect 4053 12744 4087 12778
rect 3986 12688 4087 12744
rect 3986 12654 4019 12688
rect 4053 12654 4087 12688
rect 3986 12598 4087 12654
rect 3986 12564 4019 12598
rect 4053 12564 4087 12598
rect 3986 12508 4087 12564
rect 3986 12474 4019 12508
rect 4053 12474 4087 12508
rect 3986 12418 4087 12474
rect 3986 12384 4019 12418
rect 4053 12384 4087 12418
rect 3986 12328 4087 12384
rect 3986 12294 4019 12328
rect 4053 12294 4087 12328
rect 5173 13228 5274 13284
rect 5173 13194 5206 13228
rect 5240 13194 5274 13228
rect 5173 13138 5274 13194
rect 5173 13104 5206 13138
rect 5240 13104 5274 13138
rect 5173 13048 5274 13104
rect 5173 13014 5206 13048
rect 5240 13014 5274 13048
rect 5173 12958 5274 13014
rect 5173 12924 5206 12958
rect 5240 12924 5274 12958
rect 5173 12868 5274 12924
rect 5173 12834 5206 12868
rect 5240 12834 5274 12868
rect 5173 12778 5274 12834
rect 5173 12744 5206 12778
rect 5240 12744 5274 12778
rect 5173 12688 5274 12744
rect 5173 12654 5206 12688
rect 5240 12654 5274 12688
rect 5173 12598 5274 12654
rect 5173 12564 5206 12598
rect 5240 12564 5274 12598
rect 5173 12508 5274 12564
rect 5173 12474 5206 12508
rect 5240 12474 5274 12508
rect 5173 12418 5274 12474
rect 5173 12384 5206 12418
rect 5240 12384 5274 12418
rect 5173 12328 5274 12384
rect 3986 12247 4087 12294
rect 5173 12294 5206 12328
rect 5240 12294 5274 12328
rect 5173 12247 5274 12294
rect 3986 12238 5274 12247
rect 3986 12204 4019 12238
rect 4053 12215 5206 12238
rect 4053 12204 4120 12215
rect 3986 12181 4120 12204
rect 4154 12181 4210 12215
rect 4244 12181 4300 12215
rect 4334 12181 4390 12215
rect 4424 12181 4480 12215
rect 4514 12181 4570 12215
rect 4604 12181 4660 12215
rect 4694 12181 4750 12215
rect 4784 12181 4840 12215
rect 4874 12181 4930 12215
rect 4964 12181 5020 12215
rect 5054 12181 5110 12215
rect 5144 12204 5206 12215
rect 5240 12204 5274 12238
rect 5144 12181 5274 12204
rect 3986 12146 5274 12181
rect 1266 12042 2554 12074
rect 1266 12008 1400 12042
rect 1434 12008 1490 12042
rect 1524 12008 1580 12042
rect 1614 12008 1670 12042
rect 1704 12008 1760 12042
rect 1794 12008 1850 12042
rect 1884 12008 1940 12042
rect 1974 12008 2030 12042
rect 2064 12008 2120 12042
rect 2154 12008 2210 12042
rect 2244 12008 2300 12042
rect 2334 12008 2390 12042
rect 2424 12008 2554 12042
rect 1266 11973 2554 12008
rect 1266 11958 1367 11973
rect 1266 11924 1299 11958
rect 1333 11924 1367 11958
rect 1266 11868 1367 11924
rect 2453 11958 2554 11973
rect 2453 11924 2486 11958
rect 2520 11924 2554 11958
rect 1266 11834 1299 11868
rect 1333 11834 1367 11868
rect 1266 11778 1367 11834
rect 1266 11744 1299 11778
rect 1333 11744 1367 11778
rect 1266 11688 1367 11744
rect 1266 11654 1299 11688
rect 1333 11654 1367 11688
rect 1266 11598 1367 11654
rect 1266 11564 1299 11598
rect 1333 11564 1367 11598
rect 1266 11508 1367 11564
rect 1266 11474 1299 11508
rect 1333 11474 1367 11508
rect 1266 11418 1367 11474
rect 1266 11384 1299 11418
rect 1333 11384 1367 11418
rect 1266 11328 1367 11384
rect 1266 11294 1299 11328
rect 1333 11294 1367 11328
rect 1266 11238 1367 11294
rect 1266 11204 1299 11238
rect 1333 11204 1367 11238
rect 1266 11148 1367 11204
rect 1266 11114 1299 11148
rect 1333 11114 1367 11148
rect 1266 11058 1367 11114
rect 1266 11024 1299 11058
rect 1333 11024 1367 11058
rect 1266 10968 1367 11024
rect 1266 10934 1299 10968
rect 1333 10934 1367 10968
rect 2453 11868 2554 11924
rect 2453 11834 2486 11868
rect 2520 11834 2554 11868
rect 2453 11778 2554 11834
rect 2453 11744 2486 11778
rect 2520 11744 2554 11778
rect 2453 11688 2554 11744
rect 2453 11654 2486 11688
rect 2520 11654 2554 11688
rect 2453 11598 2554 11654
rect 2453 11564 2486 11598
rect 2520 11564 2554 11598
rect 2453 11508 2554 11564
rect 2453 11474 2486 11508
rect 2520 11474 2554 11508
rect 2453 11418 2554 11474
rect 2453 11384 2486 11418
rect 2520 11384 2554 11418
rect 2453 11328 2554 11384
rect 2453 11294 2486 11328
rect 2520 11294 2554 11328
rect 2453 11238 2554 11294
rect 2453 11204 2486 11238
rect 2520 11204 2554 11238
rect 2453 11148 2554 11204
rect 2453 11114 2486 11148
rect 2520 11114 2554 11148
rect 2453 11058 2554 11114
rect 2453 11024 2486 11058
rect 2520 11024 2554 11058
rect 2453 10968 2554 11024
rect 1266 10887 1367 10934
rect 2453 10934 2486 10968
rect 2520 10934 2554 10968
rect 2453 10887 2554 10934
rect 1266 10878 2554 10887
rect 1266 10844 1299 10878
rect 1333 10855 2486 10878
rect 1333 10844 1400 10855
rect 1266 10821 1400 10844
rect 1434 10821 1490 10855
rect 1524 10821 1580 10855
rect 1614 10821 1670 10855
rect 1704 10821 1760 10855
rect 1794 10821 1850 10855
rect 1884 10821 1940 10855
rect 1974 10821 2030 10855
rect 2064 10821 2120 10855
rect 2154 10821 2210 10855
rect 2244 10821 2300 10855
rect 2334 10821 2390 10855
rect 2424 10844 2486 10855
rect 2520 10844 2554 10878
rect 2424 10821 2554 10844
rect 1266 10786 2554 10821
rect 2626 12042 3914 12074
rect 2626 12008 2760 12042
rect 2794 12008 2850 12042
rect 2884 12008 2940 12042
rect 2974 12008 3030 12042
rect 3064 12008 3120 12042
rect 3154 12008 3210 12042
rect 3244 12008 3300 12042
rect 3334 12008 3390 12042
rect 3424 12008 3480 12042
rect 3514 12008 3570 12042
rect 3604 12008 3660 12042
rect 3694 12008 3750 12042
rect 3784 12008 3914 12042
rect 2626 11973 3914 12008
rect 2626 11958 2727 11973
rect 2626 11924 2659 11958
rect 2693 11924 2727 11958
rect 2626 11868 2727 11924
rect 3813 11958 3914 11973
rect 3813 11924 3846 11958
rect 3880 11924 3914 11958
rect 2626 11834 2659 11868
rect 2693 11834 2727 11868
rect 2626 11778 2727 11834
rect 2626 11744 2659 11778
rect 2693 11744 2727 11778
rect 2626 11688 2727 11744
rect 2626 11654 2659 11688
rect 2693 11654 2727 11688
rect 2626 11598 2727 11654
rect 2626 11564 2659 11598
rect 2693 11564 2727 11598
rect 2626 11508 2727 11564
rect 2626 11474 2659 11508
rect 2693 11474 2727 11508
rect 2626 11418 2727 11474
rect 2626 11384 2659 11418
rect 2693 11384 2727 11418
rect 2626 11328 2727 11384
rect 2626 11294 2659 11328
rect 2693 11294 2727 11328
rect 2626 11238 2727 11294
rect 2626 11204 2659 11238
rect 2693 11204 2727 11238
rect 2626 11148 2727 11204
rect 2626 11114 2659 11148
rect 2693 11114 2727 11148
rect 2626 11058 2727 11114
rect 2626 11024 2659 11058
rect 2693 11024 2727 11058
rect 2626 10968 2727 11024
rect 2626 10934 2659 10968
rect 2693 10934 2727 10968
rect 3813 11868 3914 11924
rect 3813 11834 3846 11868
rect 3880 11834 3914 11868
rect 3813 11778 3914 11834
rect 3813 11744 3846 11778
rect 3880 11744 3914 11778
rect 3813 11688 3914 11744
rect 3813 11654 3846 11688
rect 3880 11654 3914 11688
rect 3813 11598 3914 11654
rect 3813 11564 3846 11598
rect 3880 11564 3914 11598
rect 3813 11508 3914 11564
rect 3813 11474 3846 11508
rect 3880 11474 3914 11508
rect 3813 11418 3914 11474
rect 3813 11384 3846 11418
rect 3880 11384 3914 11418
rect 3813 11328 3914 11384
rect 3813 11294 3846 11328
rect 3880 11294 3914 11328
rect 3813 11238 3914 11294
rect 3813 11204 3846 11238
rect 3880 11204 3914 11238
rect 3813 11148 3914 11204
rect 3813 11114 3846 11148
rect 3880 11114 3914 11148
rect 3813 11058 3914 11114
rect 3813 11024 3846 11058
rect 3880 11024 3914 11058
rect 3813 10968 3914 11024
rect 2626 10887 2727 10934
rect 3813 10934 3846 10968
rect 3880 10934 3914 10968
rect 3813 10887 3914 10934
rect 2626 10878 3914 10887
rect 2626 10844 2659 10878
rect 2693 10855 3846 10878
rect 2693 10844 2760 10855
rect 2626 10821 2760 10844
rect 2794 10821 2850 10855
rect 2884 10821 2940 10855
rect 2974 10821 3030 10855
rect 3064 10821 3120 10855
rect 3154 10821 3210 10855
rect 3244 10821 3300 10855
rect 3334 10821 3390 10855
rect 3424 10821 3480 10855
rect 3514 10821 3570 10855
rect 3604 10821 3660 10855
rect 3694 10821 3750 10855
rect 3784 10844 3846 10855
rect 3880 10844 3914 10878
rect 3784 10821 3914 10844
rect 2626 10786 3914 10821
rect 3986 12042 5274 12074
rect 3986 12008 4120 12042
rect 4154 12008 4210 12042
rect 4244 12008 4300 12042
rect 4334 12008 4390 12042
rect 4424 12008 4480 12042
rect 4514 12008 4570 12042
rect 4604 12008 4660 12042
rect 4694 12008 4750 12042
rect 4784 12008 4840 12042
rect 4874 12008 4930 12042
rect 4964 12008 5020 12042
rect 5054 12008 5110 12042
rect 5144 12008 5274 12042
rect 3986 11973 5274 12008
rect 3986 11958 4087 11973
rect 3986 11924 4019 11958
rect 4053 11924 4087 11958
rect 3986 11868 4087 11924
rect 5173 11958 5274 11973
rect 5173 11924 5206 11958
rect 5240 11924 5274 11958
rect 3986 11834 4019 11868
rect 4053 11834 4087 11868
rect 3986 11778 4087 11834
rect 3986 11744 4019 11778
rect 4053 11744 4087 11778
rect 3986 11688 4087 11744
rect 3986 11654 4019 11688
rect 4053 11654 4087 11688
rect 3986 11598 4087 11654
rect 3986 11564 4019 11598
rect 4053 11564 4087 11598
rect 3986 11508 4087 11564
rect 3986 11474 4019 11508
rect 4053 11474 4087 11508
rect 3986 11418 4087 11474
rect 3986 11384 4019 11418
rect 4053 11384 4087 11418
rect 3986 11328 4087 11384
rect 3986 11294 4019 11328
rect 4053 11294 4087 11328
rect 3986 11238 4087 11294
rect 3986 11204 4019 11238
rect 4053 11204 4087 11238
rect 3986 11148 4087 11204
rect 3986 11114 4019 11148
rect 4053 11114 4087 11148
rect 3986 11058 4087 11114
rect 3986 11024 4019 11058
rect 4053 11024 4087 11058
rect 3986 10968 4087 11024
rect 3986 10934 4019 10968
rect 4053 10934 4087 10968
rect 5173 11868 5274 11924
rect 5173 11834 5206 11868
rect 5240 11834 5274 11868
rect 5173 11778 5274 11834
rect 5173 11744 5206 11778
rect 5240 11744 5274 11778
rect 5173 11688 5274 11744
rect 5173 11654 5206 11688
rect 5240 11654 5274 11688
rect 5173 11598 5274 11654
rect 5173 11564 5206 11598
rect 5240 11564 5274 11598
rect 5173 11508 5274 11564
rect 5173 11474 5206 11508
rect 5240 11474 5274 11508
rect 5173 11418 5274 11474
rect 5173 11384 5206 11418
rect 5240 11384 5274 11418
rect 5173 11328 5274 11384
rect 5173 11294 5206 11328
rect 5240 11294 5274 11328
rect 5173 11238 5274 11294
rect 5173 11204 5206 11238
rect 5240 11204 5274 11238
rect 5173 11148 5274 11204
rect 5173 11114 5206 11148
rect 5240 11114 5274 11148
rect 5173 11058 5274 11114
rect 5173 11024 5206 11058
rect 5240 11024 5274 11058
rect 5173 10968 5274 11024
rect 3986 10887 4087 10934
rect 5173 10934 5206 10968
rect 5240 10934 5274 10968
rect 5173 10887 5274 10934
rect 3986 10878 5274 10887
rect 3986 10844 4019 10878
rect 4053 10855 5206 10878
rect 4053 10844 4120 10855
rect 3986 10821 4120 10844
rect 4154 10821 4210 10855
rect 4244 10821 4300 10855
rect 4334 10821 4390 10855
rect 4424 10821 4480 10855
rect 4514 10821 4570 10855
rect 4604 10821 4660 10855
rect 4694 10821 4750 10855
rect 4784 10821 4840 10855
rect 4874 10821 4930 10855
rect 4964 10821 5020 10855
rect 5054 10821 5110 10855
rect 5144 10844 5206 10855
rect 5240 10844 5274 10878
rect 5144 10821 5274 10844
rect 3986 10786 5274 10821
rect 5390 10260 5470 10290
rect 5390 10220 5410 10260
rect 5450 10220 5470 10260
rect 5390 10160 5470 10220
rect 5390 10120 5410 10160
rect 5450 10120 5470 10160
rect 5390 10090 5470 10120
rect 1890 9650 1970 9680
rect 1890 9610 1910 9650
rect 1950 9610 1970 9650
rect 1890 9550 1970 9610
rect 1890 9510 1910 9550
rect 1950 9510 1970 9550
rect 1890 9450 1970 9510
rect 1890 9410 1910 9450
rect 1950 9410 1970 9450
rect 1890 9350 1970 9410
rect 1890 9310 1910 9350
rect 1950 9310 1970 9350
rect 1890 9250 1970 9310
rect 1890 9210 1910 9250
rect 1950 9210 1970 9250
rect 1890 9180 1970 9210
rect 4570 9650 4650 9670
rect 4570 9610 4590 9650
rect 4630 9610 4650 9650
rect 4570 9550 4650 9610
rect 4570 9510 4590 9550
rect 4630 9510 4650 9550
rect 4570 9450 4650 9510
rect 4570 9410 4590 9450
rect 4630 9410 4650 9450
rect 4570 9350 4650 9410
rect 4570 9310 4590 9350
rect 4630 9310 4650 9350
rect 4570 9250 4650 9310
rect 4570 9210 4590 9250
rect 4630 9210 4650 9250
rect 4570 9180 4650 9210
rect 2790 8730 2870 8760
rect 2790 8690 2810 8730
rect 2850 8690 2870 8730
rect 2790 8650 2870 8690
rect 2790 8610 2810 8650
rect 2850 8610 2870 8650
rect 2790 8570 2870 8610
rect 2790 8530 2810 8570
rect 2850 8530 2870 8570
rect 2790 8500 2870 8530
rect 3670 8730 3750 8760
rect 3670 8690 3690 8730
rect 3730 8690 3750 8730
rect 3670 8650 3750 8690
rect 3670 8610 3690 8650
rect 3730 8610 3750 8650
rect 3670 8570 3750 8610
rect 8100 8580 8200 8610
rect 3670 8530 3690 8570
rect 3730 8530 3750 8570
rect 3670 8500 3750 8530
rect 8100 8530 8130 8580
rect 8170 8530 8200 8580
rect 8100 8440 8200 8530
rect 8100 8390 8130 8440
rect 8170 8390 8200 8440
rect 8100 8360 8200 8390
rect 10300 8580 10400 8610
rect 10300 8530 10330 8580
rect 10370 8530 10400 8580
rect 10300 8440 10400 8530
rect 10300 8390 10330 8440
rect 10370 8390 10400 8440
rect 10300 8360 10400 8390
rect 8150 7890 8250 7920
rect 8150 7850 8180 7890
rect 8220 7850 8250 7890
rect 8150 7820 8250 7850
rect 9130 7890 9230 7920
rect 9130 7850 9160 7890
rect 9200 7850 9230 7890
rect 9130 7820 9230 7850
rect 10430 7890 10530 7920
rect 10430 7850 10460 7890
rect 10500 7850 10530 7890
rect 10430 7820 10530 7850
rect 11410 7890 11510 7920
rect 11410 7850 11440 7890
rect 11480 7850 11510 7890
rect 11410 7820 11510 7850
rect 2060 4700 2140 4730
rect 2060 4660 2080 4700
rect 2120 4660 2140 4700
rect 2060 4600 2140 4660
rect 2060 4560 2080 4600
rect 2120 4560 2140 4600
rect 2060 4530 2140 4560
rect 2960 4700 3040 4730
rect 2960 4660 2980 4700
rect 3020 4660 3040 4700
rect 2960 4600 3040 4660
rect 2960 4560 2980 4600
rect 3020 4560 3040 4600
rect 2960 4530 3040 4560
rect 3860 4700 3940 4730
rect 3860 4660 3880 4700
rect 3920 4660 3940 4700
rect 3860 4600 3940 4660
rect 3860 4560 3880 4600
rect 3920 4560 3940 4600
rect 3860 4530 3940 4560
rect 4000 4700 4080 4730
rect 4000 4660 4020 4700
rect 4060 4660 4080 4700
rect 4000 4600 4080 4660
rect 4000 4560 4020 4600
rect 4060 4560 4080 4600
rect 4000 4530 4080 4560
rect 4440 4700 4520 4730
rect 4440 4660 4460 4700
rect 4500 4660 4520 4700
rect 4440 4600 4520 4660
rect 4440 4560 4460 4600
rect 4500 4560 4520 4600
rect 4440 4530 4520 4560
rect 4770 4700 4850 4730
rect 4770 4660 4790 4700
rect 4830 4660 4850 4700
rect 4770 4600 4850 4660
rect 4770 4560 4790 4600
rect 4830 4560 4850 4600
rect 4770 4530 4850 4560
rect 5190 4700 5270 4730
rect 5190 4660 5210 4700
rect 5250 4660 5270 4700
rect 5190 4600 5270 4660
rect 5190 4560 5210 4600
rect 5250 4560 5270 4600
rect 5190 4530 5270 4560
rect 5580 4700 5660 4730
rect 5580 4660 5600 4700
rect 5640 4660 5660 4700
rect 5580 4600 5660 4660
rect 5580 4560 5600 4600
rect 5640 4560 5660 4600
rect 5580 4530 5660 4560
rect 5970 4700 6050 4730
rect 5970 4660 5990 4700
rect 6030 4660 6050 4700
rect 5970 4600 6050 4660
rect 5970 4560 5990 4600
rect 6030 4560 6050 4600
rect 5970 4530 6050 4560
rect 7840 3350 7940 3380
rect 7840 3310 7870 3350
rect 7910 3310 7940 3350
rect 7840 3250 7940 3310
rect 7840 3210 7870 3250
rect 7910 3210 7940 3250
rect 7840 3150 7940 3210
rect 7840 3110 7870 3150
rect 7910 3110 7940 3150
rect 7840 3050 7940 3110
rect 7840 3010 7870 3050
rect 7910 3010 7940 3050
rect 7840 2980 7940 3010
rect 8920 3350 9020 3380
rect 8920 3310 8950 3350
rect 8990 3310 9020 3350
rect 8920 3250 9020 3310
rect 8920 3210 8950 3250
rect 8990 3210 9020 3250
rect 8920 3150 9020 3210
rect 8920 3110 8950 3150
rect 8990 3110 9020 3150
rect 8920 3050 9020 3110
rect 8920 3010 8950 3050
rect 8990 3010 9020 3050
rect 8920 2980 9020 3010
rect 10000 3350 10100 3380
rect 10000 3310 10030 3350
rect 10070 3310 10100 3350
rect 10000 3250 10100 3310
rect 10000 3210 10030 3250
rect 10070 3210 10100 3250
rect 10000 3150 10100 3210
rect 10000 3110 10030 3150
rect 10070 3110 10100 3150
rect 10000 3050 10100 3110
rect 10000 3010 10030 3050
rect 10070 3010 10100 3050
rect 10000 2980 10100 3010
rect 11080 3350 11180 3380
rect 11080 3310 11110 3350
rect 11150 3310 11180 3350
rect 11080 3250 11180 3310
rect 11080 3210 11110 3250
rect 11150 3210 11180 3250
rect 11080 3150 11180 3210
rect 11080 3110 11110 3150
rect 11150 3110 11180 3150
rect 11080 3050 11180 3110
rect 11080 3010 11110 3050
rect 11150 3010 11180 3050
rect 11080 2980 11180 3010
rect 2060 2900 2140 2930
rect 2060 2860 2080 2900
rect 2120 2860 2140 2900
rect 2060 2800 2140 2860
rect 2060 2760 2080 2800
rect 2120 2760 2140 2800
rect 2060 2730 2140 2760
rect 2960 2900 3040 2930
rect 2960 2860 2980 2900
rect 3020 2860 3040 2900
rect 2960 2800 3040 2860
rect 2960 2760 2980 2800
rect 3020 2760 3040 2800
rect 2960 2730 3040 2760
rect 3860 2900 3940 2930
rect 3860 2860 3880 2900
rect 3920 2860 3940 2900
rect 3860 2800 3940 2860
rect 3860 2760 3880 2800
rect 3920 2760 3940 2800
rect 3860 2730 3940 2760
rect 4260 2900 4340 2930
rect 4260 2860 4280 2900
rect 4320 2860 4340 2900
rect 4260 2800 4340 2860
rect 4260 2760 4280 2800
rect 4320 2760 4340 2800
rect 4260 2730 4340 2760
rect 4590 2900 4670 2930
rect 4590 2860 4610 2900
rect 4650 2860 4670 2900
rect 4590 2800 4670 2860
rect 4590 2760 4610 2800
rect 4650 2760 4670 2800
rect 4590 2730 4670 2760
rect 4920 2900 5000 2930
rect 4920 2860 4940 2900
rect 4980 2860 5000 2900
rect 4920 2800 5000 2860
rect 4920 2760 4940 2800
rect 4980 2760 5000 2800
rect 4920 2730 5000 2760
rect 5170 2900 5270 2930
rect 5170 2860 5200 2900
rect 5240 2860 5270 2900
rect 5170 2800 5270 2860
rect 5170 2760 5200 2800
rect 5240 2760 5270 2800
rect 5170 2730 5270 2760
rect 5950 2900 6050 2930
rect 5950 2860 5980 2900
rect 6020 2860 6050 2900
rect 5950 2800 6050 2860
rect 5950 2760 5980 2800
rect 6020 2760 6050 2800
rect 5950 2730 6050 2760
rect 6630 2900 6730 2930
rect 6630 2860 6660 2900
rect 6700 2860 6730 2900
rect 6630 2800 6730 2860
rect 6630 2760 6660 2800
rect 6700 2760 6730 2800
rect 6630 2730 6730 2760
rect 17350 2650 17450 2680
rect 17350 2610 17380 2650
rect 17420 2610 17450 2650
rect 17350 2580 17450 2610
rect 12590 1970 12670 2000
rect 12590 1930 12610 1970
rect 12650 1930 12670 1970
rect 12590 1870 12670 1930
rect 12590 1830 12610 1870
rect 12650 1830 12670 1870
rect 12590 1800 12670 1830
rect 13190 1970 13270 2000
rect 13190 1930 13210 1970
rect 13250 1930 13270 1970
rect 13190 1870 13270 1930
rect 13190 1830 13210 1870
rect 13250 1830 13270 1870
rect 13190 1800 13270 1830
rect 13790 1970 13870 2000
rect 13790 1930 13810 1970
rect 13850 1930 13870 1970
rect 13790 1870 13870 1930
rect 13790 1830 13810 1870
rect 13850 1830 13870 1870
rect 13790 1800 13870 1830
rect 12590 1640 12670 1670
rect 12590 1600 12610 1640
rect 12650 1600 12670 1640
rect 12590 1570 12670 1600
rect 13190 1640 13270 1670
rect 13190 1600 13210 1640
rect 13250 1600 13270 1640
rect 13190 1570 13270 1600
rect 13790 1640 13870 1670
rect 13790 1600 13810 1640
rect 13850 1600 13870 1640
rect 13790 1570 13870 1600
rect 8320 1500 8400 1530
rect 8320 1460 8340 1500
rect 8380 1460 8400 1500
rect 5080 1410 5160 1440
rect 5080 1370 5100 1410
rect 5140 1370 5160 1410
rect 5080 1340 5160 1370
rect 6530 1410 6610 1440
rect 6530 1370 6550 1410
rect 6590 1370 6610 1410
rect 6530 1340 6610 1370
rect 8320 1430 8400 1460
rect 9620 1500 9700 1530
rect 9620 1460 9640 1500
rect 9680 1460 9700 1500
rect 9620 1430 9700 1460
rect 10920 1500 11000 1530
rect 10920 1460 10940 1500
rect 10980 1460 11000 1500
rect 10920 1430 11000 1460
<< nsubdiff >>
rect 1429 14612 2391 14631
rect 1429 14578 1540 14612
rect 1574 14578 1630 14612
rect 1664 14578 1720 14612
rect 1754 14578 1810 14612
rect 1844 14578 1900 14612
rect 1934 14578 1990 14612
rect 2024 14578 2080 14612
rect 2114 14578 2170 14612
rect 2204 14578 2260 14612
rect 2294 14578 2391 14612
rect 1429 14559 2391 14578
rect 1429 14518 1501 14559
rect 1429 14484 1448 14518
rect 1482 14484 1501 14518
rect 2319 14499 2391 14559
rect 1429 14428 1501 14484
rect 1429 14394 1448 14428
rect 1482 14394 1501 14428
rect 1429 14338 1501 14394
rect 1429 14304 1448 14338
rect 1482 14304 1501 14338
rect 1429 14248 1501 14304
rect 1429 14214 1448 14248
rect 1482 14214 1501 14248
rect 1429 14158 1501 14214
rect 1429 14124 1448 14158
rect 1482 14124 1501 14158
rect 1429 14068 1501 14124
rect 1429 14034 1448 14068
rect 1482 14034 1501 14068
rect 1429 13978 1501 14034
rect 1429 13944 1448 13978
rect 1482 13944 1501 13978
rect 1429 13888 1501 13944
rect 1429 13854 1448 13888
rect 1482 13854 1501 13888
rect 1429 13798 1501 13854
rect 2319 14465 2338 14499
rect 2372 14465 2391 14499
rect 2319 14409 2391 14465
rect 2319 14375 2338 14409
rect 2372 14375 2391 14409
rect 2319 14319 2391 14375
rect 2319 14285 2338 14319
rect 2372 14285 2391 14319
rect 2319 14229 2391 14285
rect 2319 14195 2338 14229
rect 2372 14195 2391 14229
rect 2319 14139 2391 14195
rect 2319 14105 2338 14139
rect 2372 14105 2391 14139
rect 2319 14049 2391 14105
rect 2319 14015 2338 14049
rect 2372 14015 2391 14049
rect 2319 13959 2391 14015
rect 2319 13925 2338 13959
rect 2372 13925 2391 13959
rect 2319 13869 2391 13925
rect 2319 13835 2338 13869
rect 2372 13835 2391 13869
rect 1429 13764 1448 13798
rect 1482 13764 1501 13798
rect 1429 13741 1501 13764
rect 2319 13779 2391 13835
rect 2319 13745 2338 13779
rect 2372 13745 2391 13779
rect 2319 13741 2391 13745
rect 1429 13722 2391 13741
rect 1429 13688 1506 13722
rect 1540 13688 1596 13722
rect 1630 13688 1686 13722
rect 1720 13688 1776 13722
rect 1810 13688 1866 13722
rect 1900 13688 1956 13722
rect 1990 13688 2046 13722
rect 2080 13688 2136 13722
rect 2170 13688 2226 13722
rect 2260 13688 2391 13722
rect 1429 13669 2391 13688
rect 2789 14612 3751 14631
rect 2789 14578 2900 14612
rect 2934 14578 2990 14612
rect 3024 14578 3080 14612
rect 3114 14578 3170 14612
rect 3204 14578 3260 14612
rect 3294 14578 3350 14612
rect 3384 14578 3440 14612
rect 3474 14578 3530 14612
rect 3564 14578 3620 14612
rect 3654 14578 3751 14612
rect 2789 14559 3751 14578
rect 2789 14518 2861 14559
rect 2789 14484 2808 14518
rect 2842 14484 2861 14518
rect 3679 14499 3751 14559
rect 2789 14428 2861 14484
rect 2789 14394 2808 14428
rect 2842 14394 2861 14428
rect 2789 14338 2861 14394
rect 2789 14304 2808 14338
rect 2842 14304 2861 14338
rect 2789 14248 2861 14304
rect 2789 14214 2808 14248
rect 2842 14214 2861 14248
rect 2789 14158 2861 14214
rect 2789 14124 2808 14158
rect 2842 14124 2861 14158
rect 2789 14068 2861 14124
rect 2789 14034 2808 14068
rect 2842 14034 2861 14068
rect 2789 13978 2861 14034
rect 2789 13944 2808 13978
rect 2842 13944 2861 13978
rect 2789 13888 2861 13944
rect 2789 13854 2808 13888
rect 2842 13854 2861 13888
rect 2789 13798 2861 13854
rect 3679 14465 3698 14499
rect 3732 14465 3751 14499
rect 3679 14409 3751 14465
rect 3679 14375 3698 14409
rect 3732 14375 3751 14409
rect 3679 14319 3751 14375
rect 3679 14285 3698 14319
rect 3732 14285 3751 14319
rect 3679 14229 3751 14285
rect 3679 14195 3698 14229
rect 3732 14195 3751 14229
rect 3679 14139 3751 14195
rect 3679 14105 3698 14139
rect 3732 14105 3751 14139
rect 3679 14049 3751 14105
rect 3679 14015 3698 14049
rect 3732 14015 3751 14049
rect 3679 13959 3751 14015
rect 3679 13925 3698 13959
rect 3732 13925 3751 13959
rect 3679 13869 3751 13925
rect 3679 13835 3698 13869
rect 3732 13835 3751 13869
rect 2789 13764 2808 13798
rect 2842 13764 2861 13798
rect 2789 13741 2861 13764
rect 3679 13779 3751 13835
rect 3679 13745 3698 13779
rect 3732 13745 3751 13779
rect 3679 13741 3751 13745
rect 2789 13722 3751 13741
rect 2789 13688 2866 13722
rect 2900 13688 2956 13722
rect 2990 13688 3046 13722
rect 3080 13688 3136 13722
rect 3170 13688 3226 13722
rect 3260 13688 3316 13722
rect 3350 13688 3406 13722
rect 3440 13688 3496 13722
rect 3530 13688 3586 13722
rect 3620 13688 3751 13722
rect 2789 13669 3751 13688
rect 4149 14612 5111 14631
rect 4149 14578 4260 14612
rect 4294 14578 4350 14612
rect 4384 14578 4440 14612
rect 4474 14578 4530 14612
rect 4564 14578 4620 14612
rect 4654 14578 4710 14612
rect 4744 14578 4800 14612
rect 4834 14578 4890 14612
rect 4924 14578 4980 14612
rect 5014 14578 5111 14612
rect 4149 14559 5111 14578
rect 4149 14518 4221 14559
rect 4149 14484 4168 14518
rect 4202 14484 4221 14518
rect 5039 14499 5111 14559
rect 4149 14428 4221 14484
rect 4149 14394 4168 14428
rect 4202 14394 4221 14428
rect 4149 14338 4221 14394
rect 4149 14304 4168 14338
rect 4202 14304 4221 14338
rect 4149 14248 4221 14304
rect 4149 14214 4168 14248
rect 4202 14214 4221 14248
rect 4149 14158 4221 14214
rect 4149 14124 4168 14158
rect 4202 14124 4221 14158
rect 4149 14068 4221 14124
rect 4149 14034 4168 14068
rect 4202 14034 4221 14068
rect 4149 13978 4221 14034
rect 4149 13944 4168 13978
rect 4202 13944 4221 13978
rect 4149 13888 4221 13944
rect 4149 13854 4168 13888
rect 4202 13854 4221 13888
rect 4149 13798 4221 13854
rect 5039 14465 5058 14499
rect 5092 14465 5111 14499
rect 5039 14409 5111 14465
rect 5039 14375 5058 14409
rect 5092 14375 5111 14409
rect 5039 14319 5111 14375
rect 5039 14285 5058 14319
rect 5092 14285 5111 14319
rect 5039 14229 5111 14285
rect 5039 14195 5058 14229
rect 5092 14195 5111 14229
rect 5039 14139 5111 14195
rect 5039 14105 5058 14139
rect 5092 14105 5111 14139
rect 5039 14049 5111 14105
rect 5039 14015 5058 14049
rect 5092 14015 5111 14049
rect 5039 13959 5111 14015
rect 5039 13925 5058 13959
rect 5092 13925 5111 13959
rect 5039 13869 5111 13925
rect 5039 13835 5058 13869
rect 5092 13835 5111 13869
rect 4149 13764 4168 13798
rect 4202 13764 4221 13798
rect 4149 13741 4221 13764
rect 5039 13779 5111 13835
rect 5039 13745 5058 13779
rect 5092 13745 5111 13779
rect 5039 13741 5111 13745
rect 4149 13722 5111 13741
rect 4149 13688 4226 13722
rect 4260 13688 4316 13722
rect 4350 13688 4406 13722
rect 4440 13688 4496 13722
rect 4530 13688 4586 13722
rect 4620 13688 4676 13722
rect 4710 13688 4766 13722
rect 4800 13688 4856 13722
rect 4890 13688 4946 13722
rect 4980 13688 5111 13722
rect 4149 13669 5111 13688
rect 1429 13252 2391 13271
rect 1429 13218 1540 13252
rect 1574 13218 1630 13252
rect 1664 13218 1720 13252
rect 1754 13218 1810 13252
rect 1844 13218 1900 13252
rect 1934 13218 1990 13252
rect 2024 13218 2080 13252
rect 2114 13218 2170 13252
rect 2204 13218 2260 13252
rect 2294 13218 2391 13252
rect 1429 13199 2391 13218
rect 1429 13158 1501 13199
rect 1429 13124 1448 13158
rect 1482 13124 1501 13158
rect 2319 13139 2391 13199
rect 1429 13068 1501 13124
rect 1429 13034 1448 13068
rect 1482 13034 1501 13068
rect 1429 12978 1501 13034
rect 1429 12944 1448 12978
rect 1482 12944 1501 12978
rect 1429 12888 1501 12944
rect 1429 12854 1448 12888
rect 1482 12854 1501 12888
rect 1429 12798 1501 12854
rect 1429 12764 1448 12798
rect 1482 12764 1501 12798
rect 1429 12708 1501 12764
rect 1429 12674 1448 12708
rect 1482 12674 1501 12708
rect 1429 12618 1501 12674
rect 1429 12584 1448 12618
rect 1482 12584 1501 12618
rect 1429 12528 1501 12584
rect 1429 12494 1448 12528
rect 1482 12494 1501 12528
rect 1429 12438 1501 12494
rect 2319 13105 2338 13139
rect 2372 13105 2391 13139
rect 2319 13049 2391 13105
rect 2319 13015 2338 13049
rect 2372 13015 2391 13049
rect 2319 12959 2391 13015
rect 2319 12925 2338 12959
rect 2372 12925 2391 12959
rect 2319 12869 2391 12925
rect 2319 12835 2338 12869
rect 2372 12835 2391 12869
rect 2319 12779 2391 12835
rect 2319 12745 2338 12779
rect 2372 12745 2391 12779
rect 2319 12689 2391 12745
rect 2319 12655 2338 12689
rect 2372 12655 2391 12689
rect 2319 12599 2391 12655
rect 2319 12565 2338 12599
rect 2372 12565 2391 12599
rect 2319 12509 2391 12565
rect 2319 12475 2338 12509
rect 2372 12475 2391 12509
rect 1429 12404 1448 12438
rect 1482 12404 1501 12438
rect 1429 12381 1501 12404
rect 2319 12419 2391 12475
rect 2319 12385 2338 12419
rect 2372 12385 2391 12419
rect 2319 12381 2391 12385
rect 1429 12362 2391 12381
rect 1429 12328 1506 12362
rect 1540 12328 1596 12362
rect 1630 12328 1686 12362
rect 1720 12328 1776 12362
rect 1810 12328 1866 12362
rect 1900 12328 1956 12362
rect 1990 12328 2046 12362
rect 2080 12328 2136 12362
rect 2170 12328 2226 12362
rect 2260 12328 2391 12362
rect 1429 12309 2391 12328
rect 2789 13252 3751 13271
rect 2789 13218 2900 13252
rect 2934 13218 2990 13252
rect 3024 13218 3080 13252
rect 3114 13218 3170 13252
rect 3204 13218 3260 13252
rect 3294 13218 3350 13252
rect 3384 13218 3440 13252
rect 3474 13218 3530 13252
rect 3564 13218 3620 13252
rect 3654 13218 3751 13252
rect 2789 13199 3751 13218
rect 2789 13158 2861 13199
rect 2789 13124 2808 13158
rect 2842 13124 2861 13158
rect 3679 13139 3751 13199
rect 2789 13068 2861 13124
rect 2789 13034 2808 13068
rect 2842 13034 2861 13068
rect 2789 12978 2861 13034
rect 2789 12944 2808 12978
rect 2842 12944 2861 12978
rect 2789 12888 2861 12944
rect 2789 12854 2808 12888
rect 2842 12854 2861 12888
rect 2789 12798 2861 12854
rect 2789 12764 2808 12798
rect 2842 12764 2861 12798
rect 2789 12708 2861 12764
rect 2789 12674 2808 12708
rect 2842 12674 2861 12708
rect 2789 12618 2861 12674
rect 2789 12584 2808 12618
rect 2842 12584 2861 12618
rect 2789 12528 2861 12584
rect 2789 12494 2808 12528
rect 2842 12494 2861 12528
rect 2789 12438 2861 12494
rect 3679 13105 3698 13139
rect 3732 13105 3751 13139
rect 3679 13049 3751 13105
rect 3679 13015 3698 13049
rect 3732 13015 3751 13049
rect 3679 12959 3751 13015
rect 3679 12925 3698 12959
rect 3732 12925 3751 12959
rect 3679 12869 3751 12925
rect 3679 12835 3698 12869
rect 3732 12835 3751 12869
rect 3679 12779 3751 12835
rect 3679 12745 3698 12779
rect 3732 12745 3751 12779
rect 3679 12689 3751 12745
rect 3679 12655 3698 12689
rect 3732 12655 3751 12689
rect 3679 12599 3751 12655
rect 3679 12565 3698 12599
rect 3732 12565 3751 12599
rect 3679 12509 3751 12565
rect 3679 12475 3698 12509
rect 3732 12475 3751 12509
rect 2789 12404 2808 12438
rect 2842 12404 2861 12438
rect 2789 12381 2861 12404
rect 3679 12419 3751 12475
rect 3679 12385 3698 12419
rect 3732 12385 3751 12419
rect 3679 12381 3751 12385
rect 2789 12362 3751 12381
rect 2789 12328 2866 12362
rect 2900 12328 2956 12362
rect 2990 12328 3046 12362
rect 3080 12328 3136 12362
rect 3170 12328 3226 12362
rect 3260 12328 3316 12362
rect 3350 12328 3406 12362
rect 3440 12328 3496 12362
rect 3530 12328 3586 12362
rect 3620 12328 3751 12362
rect 2789 12309 3751 12328
rect 4149 13252 5111 13271
rect 4149 13218 4260 13252
rect 4294 13218 4350 13252
rect 4384 13218 4440 13252
rect 4474 13218 4530 13252
rect 4564 13218 4620 13252
rect 4654 13218 4710 13252
rect 4744 13218 4800 13252
rect 4834 13218 4890 13252
rect 4924 13218 4980 13252
rect 5014 13218 5111 13252
rect 4149 13199 5111 13218
rect 4149 13158 4221 13199
rect 4149 13124 4168 13158
rect 4202 13124 4221 13158
rect 5039 13139 5111 13199
rect 4149 13068 4221 13124
rect 4149 13034 4168 13068
rect 4202 13034 4221 13068
rect 4149 12978 4221 13034
rect 4149 12944 4168 12978
rect 4202 12944 4221 12978
rect 4149 12888 4221 12944
rect 4149 12854 4168 12888
rect 4202 12854 4221 12888
rect 4149 12798 4221 12854
rect 4149 12764 4168 12798
rect 4202 12764 4221 12798
rect 4149 12708 4221 12764
rect 4149 12674 4168 12708
rect 4202 12674 4221 12708
rect 4149 12618 4221 12674
rect 4149 12584 4168 12618
rect 4202 12584 4221 12618
rect 4149 12528 4221 12584
rect 4149 12494 4168 12528
rect 4202 12494 4221 12528
rect 4149 12438 4221 12494
rect 5039 13105 5058 13139
rect 5092 13105 5111 13139
rect 5039 13049 5111 13105
rect 5039 13015 5058 13049
rect 5092 13015 5111 13049
rect 5039 12959 5111 13015
rect 5039 12925 5058 12959
rect 5092 12925 5111 12959
rect 5039 12869 5111 12925
rect 5039 12835 5058 12869
rect 5092 12835 5111 12869
rect 5039 12779 5111 12835
rect 5039 12745 5058 12779
rect 5092 12745 5111 12779
rect 5039 12689 5111 12745
rect 5039 12655 5058 12689
rect 5092 12655 5111 12689
rect 5039 12599 5111 12655
rect 5039 12565 5058 12599
rect 5092 12565 5111 12599
rect 5039 12509 5111 12565
rect 5039 12475 5058 12509
rect 5092 12475 5111 12509
rect 4149 12404 4168 12438
rect 4202 12404 4221 12438
rect 4149 12381 4221 12404
rect 5039 12419 5111 12475
rect 5039 12385 5058 12419
rect 5092 12385 5111 12419
rect 5039 12381 5111 12385
rect 4149 12362 5111 12381
rect 4149 12328 4226 12362
rect 4260 12328 4316 12362
rect 4350 12328 4406 12362
rect 4440 12328 4496 12362
rect 4530 12328 4586 12362
rect 4620 12328 4676 12362
rect 4710 12328 4766 12362
rect 4800 12328 4856 12362
rect 4890 12328 4946 12362
rect 4980 12328 5111 12362
rect 4149 12309 5111 12328
rect 1429 11892 2391 11911
rect 1429 11858 1540 11892
rect 1574 11858 1630 11892
rect 1664 11858 1720 11892
rect 1754 11858 1810 11892
rect 1844 11858 1900 11892
rect 1934 11858 1990 11892
rect 2024 11858 2080 11892
rect 2114 11858 2170 11892
rect 2204 11858 2260 11892
rect 2294 11858 2391 11892
rect 1429 11839 2391 11858
rect 1429 11798 1501 11839
rect 1429 11764 1448 11798
rect 1482 11764 1501 11798
rect 2319 11779 2391 11839
rect 1429 11708 1501 11764
rect 1429 11674 1448 11708
rect 1482 11674 1501 11708
rect 1429 11618 1501 11674
rect 1429 11584 1448 11618
rect 1482 11584 1501 11618
rect 1429 11528 1501 11584
rect 1429 11494 1448 11528
rect 1482 11494 1501 11528
rect 1429 11438 1501 11494
rect 1429 11404 1448 11438
rect 1482 11404 1501 11438
rect 1429 11348 1501 11404
rect 1429 11314 1448 11348
rect 1482 11314 1501 11348
rect 1429 11258 1501 11314
rect 1429 11224 1448 11258
rect 1482 11224 1501 11258
rect 1429 11168 1501 11224
rect 1429 11134 1448 11168
rect 1482 11134 1501 11168
rect 1429 11078 1501 11134
rect 2319 11745 2338 11779
rect 2372 11745 2391 11779
rect 2319 11689 2391 11745
rect 2319 11655 2338 11689
rect 2372 11655 2391 11689
rect 2319 11599 2391 11655
rect 2319 11565 2338 11599
rect 2372 11565 2391 11599
rect 2319 11509 2391 11565
rect 2319 11475 2338 11509
rect 2372 11475 2391 11509
rect 2319 11419 2391 11475
rect 2319 11385 2338 11419
rect 2372 11385 2391 11419
rect 2319 11329 2391 11385
rect 2319 11295 2338 11329
rect 2372 11295 2391 11329
rect 2319 11239 2391 11295
rect 2319 11205 2338 11239
rect 2372 11205 2391 11239
rect 2319 11149 2391 11205
rect 2319 11115 2338 11149
rect 2372 11115 2391 11149
rect 1429 11044 1448 11078
rect 1482 11044 1501 11078
rect 1429 11021 1501 11044
rect 2319 11059 2391 11115
rect 2319 11025 2338 11059
rect 2372 11025 2391 11059
rect 2319 11021 2391 11025
rect 1429 11002 2391 11021
rect 1429 10968 1506 11002
rect 1540 10968 1596 11002
rect 1630 10968 1686 11002
rect 1720 10968 1776 11002
rect 1810 10968 1866 11002
rect 1900 10968 1956 11002
rect 1990 10968 2046 11002
rect 2080 10968 2136 11002
rect 2170 10968 2226 11002
rect 2260 10968 2391 11002
rect 1429 10949 2391 10968
rect 2789 11892 3751 11911
rect 2789 11858 2900 11892
rect 2934 11858 2990 11892
rect 3024 11858 3080 11892
rect 3114 11858 3170 11892
rect 3204 11858 3260 11892
rect 3294 11858 3350 11892
rect 3384 11858 3440 11892
rect 3474 11858 3530 11892
rect 3564 11858 3620 11892
rect 3654 11858 3751 11892
rect 2789 11839 3751 11858
rect 2789 11798 2861 11839
rect 2789 11764 2808 11798
rect 2842 11764 2861 11798
rect 3679 11779 3751 11839
rect 2789 11708 2861 11764
rect 2789 11674 2808 11708
rect 2842 11674 2861 11708
rect 2789 11618 2861 11674
rect 2789 11584 2808 11618
rect 2842 11584 2861 11618
rect 2789 11528 2861 11584
rect 2789 11494 2808 11528
rect 2842 11494 2861 11528
rect 2789 11438 2861 11494
rect 2789 11404 2808 11438
rect 2842 11404 2861 11438
rect 2789 11348 2861 11404
rect 2789 11314 2808 11348
rect 2842 11314 2861 11348
rect 2789 11258 2861 11314
rect 2789 11224 2808 11258
rect 2842 11224 2861 11258
rect 2789 11168 2861 11224
rect 2789 11134 2808 11168
rect 2842 11134 2861 11168
rect 2789 11078 2861 11134
rect 3679 11745 3698 11779
rect 3732 11745 3751 11779
rect 3679 11689 3751 11745
rect 3679 11655 3698 11689
rect 3732 11655 3751 11689
rect 3679 11599 3751 11655
rect 3679 11565 3698 11599
rect 3732 11565 3751 11599
rect 3679 11509 3751 11565
rect 3679 11475 3698 11509
rect 3732 11475 3751 11509
rect 3679 11419 3751 11475
rect 3679 11385 3698 11419
rect 3732 11385 3751 11419
rect 3679 11329 3751 11385
rect 3679 11295 3698 11329
rect 3732 11295 3751 11329
rect 3679 11239 3751 11295
rect 3679 11205 3698 11239
rect 3732 11205 3751 11239
rect 3679 11149 3751 11205
rect 3679 11115 3698 11149
rect 3732 11115 3751 11149
rect 2789 11044 2808 11078
rect 2842 11044 2861 11078
rect 2789 11021 2861 11044
rect 3679 11059 3751 11115
rect 3679 11025 3698 11059
rect 3732 11025 3751 11059
rect 3679 11021 3751 11025
rect 2789 11002 3751 11021
rect 2789 10968 2866 11002
rect 2900 10968 2956 11002
rect 2990 10968 3046 11002
rect 3080 10968 3136 11002
rect 3170 10968 3226 11002
rect 3260 10968 3316 11002
rect 3350 10968 3406 11002
rect 3440 10968 3496 11002
rect 3530 10968 3586 11002
rect 3620 10968 3751 11002
rect 2789 10949 3751 10968
rect 4149 11892 5111 11911
rect 4149 11858 4260 11892
rect 4294 11858 4350 11892
rect 4384 11858 4440 11892
rect 4474 11858 4530 11892
rect 4564 11858 4620 11892
rect 4654 11858 4710 11892
rect 4744 11858 4800 11892
rect 4834 11858 4890 11892
rect 4924 11858 4980 11892
rect 5014 11858 5111 11892
rect 4149 11839 5111 11858
rect 4149 11798 4221 11839
rect 4149 11764 4168 11798
rect 4202 11764 4221 11798
rect 5039 11779 5111 11839
rect 4149 11708 4221 11764
rect 4149 11674 4168 11708
rect 4202 11674 4221 11708
rect 4149 11618 4221 11674
rect 4149 11584 4168 11618
rect 4202 11584 4221 11618
rect 4149 11528 4221 11584
rect 4149 11494 4168 11528
rect 4202 11494 4221 11528
rect 4149 11438 4221 11494
rect 4149 11404 4168 11438
rect 4202 11404 4221 11438
rect 4149 11348 4221 11404
rect 4149 11314 4168 11348
rect 4202 11314 4221 11348
rect 4149 11258 4221 11314
rect 4149 11224 4168 11258
rect 4202 11224 4221 11258
rect 4149 11168 4221 11224
rect 4149 11134 4168 11168
rect 4202 11134 4221 11168
rect 4149 11078 4221 11134
rect 5039 11745 5058 11779
rect 5092 11745 5111 11779
rect 5039 11689 5111 11745
rect 5039 11655 5058 11689
rect 5092 11655 5111 11689
rect 5039 11599 5111 11655
rect 5039 11565 5058 11599
rect 5092 11565 5111 11599
rect 5039 11509 5111 11565
rect 5039 11475 5058 11509
rect 5092 11475 5111 11509
rect 5039 11419 5111 11475
rect 5039 11385 5058 11419
rect 5092 11385 5111 11419
rect 5039 11329 5111 11385
rect 5039 11295 5058 11329
rect 5092 11295 5111 11329
rect 5039 11239 5111 11295
rect 5039 11205 5058 11239
rect 5092 11205 5111 11239
rect 5039 11149 5111 11205
rect 5039 11115 5058 11149
rect 5092 11115 5111 11149
rect 4149 11044 4168 11078
rect 4202 11044 4221 11078
rect 4149 11021 4221 11044
rect 5039 11059 5111 11115
rect 5039 11025 5058 11059
rect 5092 11025 5111 11059
rect 5039 11021 5111 11025
rect 4149 11002 5111 11021
rect 4149 10968 4226 11002
rect 4260 10968 4316 11002
rect 4350 10968 4406 11002
rect 4440 10968 4496 11002
rect 4530 10968 4586 11002
rect 4620 10968 4676 11002
rect 4710 10968 4766 11002
rect 4800 10968 4856 11002
rect 4890 10968 4946 11002
rect 4980 10968 5111 11002
rect 4149 10949 5111 10968
rect 430 7800 510 7830
rect 430 7760 450 7800
rect 490 7760 510 7800
rect 430 7700 510 7760
rect 430 7660 450 7700
rect 490 7660 510 7700
rect 430 7630 510 7660
rect 2990 7800 3070 7830
rect 2990 7760 3010 7800
rect 3050 7760 3070 7800
rect 2990 7700 3070 7760
rect 2990 7660 3010 7700
rect 3050 7660 3070 7700
rect 2990 7630 3070 7660
rect 3470 7800 3550 7830
rect 3470 7760 3490 7800
rect 3530 7760 3550 7800
rect 3470 7700 3550 7760
rect 3470 7660 3490 7700
rect 3530 7660 3550 7700
rect 3470 7630 3550 7660
rect 6030 7800 6110 7830
rect 6030 7760 6050 7800
rect 6090 7760 6110 7800
rect 6030 7700 6110 7760
rect 6030 7660 6050 7700
rect 6090 7660 6110 7700
rect 6030 7630 6110 7660
rect 9290 7320 9390 7350
rect 9290 7280 9320 7320
rect 9360 7280 9390 7320
rect 9290 7220 9390 7280
rect 9290 7180 9320 7220
rect 9360 7180 9390 7220
rect 9290 7150 9390 7180
rect 10270 7320 10370 7350
rect 10270 7280 10300 7320
rect 10340 7280 10370 7320
rect 10270 7220 10370 7280
rect 10270 7180 10300 7220
rect 10340 7180 10370 7220
rect 10270 7150 10370 7180
rect 10430 7320 10530 7350
rect 10430 7280 10460 7320
rect 10500 7280 10530 7320
rect 10430 7220 10530 7280
rect 10430 7180 10460 7220
rect 10500 7180 10530 7220
rect 10430 7150 10530 7180
rect 11410 7320 11510 7350
rect 11410 7280 11440 7320
rect 11480 7280 11510 7320
rect 11410 7220 11510 7280
rect 11410 7180 11440 7220
rect 11480 7180 11510 7220
rect 11410 7150 11510 7180
rect 8220 6670 8320 6700
rect 1530 6640 1610 6670
rect 1530 6600 1550 6640
rect 1590 6600 1610 6640
rect 1530 6540 1610 6600
rect 1530 6500 1550 6540
rect 1590 6500 1610 6540
rect 1530 6440 1610 6500
rect 1530 6400 1550 6440
rect 1590 6400 1610 6440
rect 1530 6340 1610 6400
rect 1530 6300 1550 6340
rect 1590 6300 1610 6340
rect 1530 6240 1610 6300
rect 1530 6200 1550 6240
rect 1590 6200 1610 6240
rect 1530 6140 1610 6200
rect 1530 6100 1550 6140
rect 1590 6100 1610 6140
rect 1530 6070 1610 6100
rect 4930 6640 5010 6670
rect 4930 6600 4950 6640
rect 4990 6600 5010 6640
rect 4930 6540 5010 6600
rect 8220 6630 8250 6670
rect 8290 6630 8320 6670
rect 4930 6500 4950 6540
rect 4990 6500 5010 6540
rect 8220 6570 8320 6630
rect 8220 6530 8250 6570
rect 8290 6530 8320 6570
rect 4930 6440 5010 6500
rect 8220 6470 8320 6530
rect 4930 6400 4950 6440
rect 4990 6400 5010 6440
rect 4930 6340 5010 6400
rect 4930 6300 4950 6340
rect 4990 6300 5010 6340
rect 4930 6240 5010 6300
rect 5390 6440 5470 6470
rect 5390 6400 5410 6440
rect 5450 6400 5470 6440
rect 5390 6340 5470 6400
rect 5390 6300 5410 6340
rect 5450 6300 5470 6340
rect 5390 6270 5470 6300
rect 6000 6440 6080 6470
rect 6000 6400 6020 6440
rect 6060 6400 6080 6440
rect 6000 6340 6080 6400
rect 6000 6300 6020 6340
rect 6060 6300 6080 6340
rect 6000 6270 6080 6300
rect 8220 6430 8250 6470
rect 8290 6430 8320 6470
rect 8220 6370 8320 6430
rect 8220 6330 8250 6370
rect 8290 6330 8320 6370
rect 8220 6270 8320 6330
rect 4930 6200 4950 6240
rect 4990 6200 5010 6240
rect 4930 6140 5010 6200
rect 8220 6230 8250 6270
rect 8290 6230 8320 6270
rect 8220 6200 8320 6230
rect 10420 6670 10520 6700
rect 10420 6630 10450 6670
rect 10490 6630 10520 6670
rect 10420 6570 10520 6630
rect 10420 6530 10450 6570
rect 10490 6530 10520 6570
rect 10420 6470 10520 6530
rect 10420 6430 10450 6470
rect 10490 6430 10520 6470
rect 10420 6370 10520 6430
rect 10420 6330 10450 6370
rect 10490 6330 10520 6370
rect 10420 6270 10520 6330
rect 10420 6230 10450 6270
rect 10490 6230 10520 6270
rect 10420 6200 10520 6230
rect 4930 6100 4950 6140
rect 4990 6100 5010 6140
rect 4930 6070 5010 6100
rect 1540 5640 1620 5670
rect 1540 5600 1560 5640
rect 1600 5600 1620 5640
rect 1540 5540 1620 5600
rect 1540 5500 1560 5540
rect 1600 5500 1620 5540
rect 1540 5470 1620 5500
rect 3020 5640 3100 5670
rect 3020 5600 3040 5640
rect 3080 5600 3100 5640
rect 3020 5540 3100 5600
rect 3020 5500 3040 5540
rect 3080 5500 3100 5540
rect 3020 5470 3100 5500
rect 3440 5640 3520 5670
rect 3440 5600 3460 5640
rect 3500 5600 3520 5640
rect 3440 5540 3520 5600
rect 3440 5500 3460 5540
rect 3500 5500 3520 5540
rect 3440 5470 3520 5500
rect 4920 5640 5000 5670
rect 4920 5600 4940 5640
rect 4980 5600 5000 5640
rect 4920 5540 5000 5600
rect 4920 5500 4940 5540
rect 4980 5500 5000 5540
rect 4920 5470 5000 5500
rect 2060 4280 2140 4310
rect 2060 4240 2080 4280
rect 2120 4240 2140 4280
rect 2060 4180 2140 4240
rect 2060 4140 2080 4180
rect 2120 4140 2140 4180
rect 2060 4080 2140 4140
rect 2060 4040 2080 4080
rect 2120 4040 2140 4080
rect 2060 3980 2140 4040
rect 2060 3940 2080 3980
rect 2120 3940 2140 3980
rect 2060 3910 2140 3940
rect 2960 4280 3040 4310
rect 2960 4240 2980 4280
rect 3020 4240 3040 4280
rect 2960 4180 3040 4240
rect 2960 4140 2980 4180
rect 3020 4140 3040 4180
rect 2960 4080 3040 4140
rect 2960 4040 2980 4080
rect 3020 4040 3040 4080
rect 2960 3980 3040 4040
rect 2960 3940 2980 3980
rect 3020 3940 3040 3980
rect 2960 3910 3040 3940
rect 8040 4330 8140 4360
rect 3860 4280 3940 4310
rect 3860 4240 3880 4280
rect 3920 4240 3940 4280
rect 3860 4180 3940 4240
rect 3860 4140 3880 4180
rect 3920 4140 3940 4180
rect 3860 4080 3940 4140
rect 3860 4040 3880 4080
rect 3920 4040 3940 4080
rect 3860 3980 3940 4040
rect 3860 3940 3880 3980
rect 3920 3940 3940 3980
rect 3860 3910 3940 3940
rect 4000 4280 4080 4310
rect 4000 4240 4020 4280
rect 4060 4240 4080 4280
rect 4000 4180 4080 4240
rect 4000 4140 4020 4180
rect 4060 4140 4080 4180
rect 4000 4080 4080 4140
rect 4000 4040 4020 4080
rect 4060 4040 4080 4080
rect 4000 3980 4080 4040
rect 4000 3940 4020 3980
rect 4060 3940 4080 3980
rect 4000 3920 4080 3940
rect 4000 3910 4060 3920
rect 4440 4280 4520 4310
rect 4440 4240 4460 4280
rect 4500 4240 4520 4280
rect 4440 4180 4520 4240
rect 4440 4140 4460 4180
rect 4500 4140 4520 4180
rect 4440 4080 4520 4140
rect 4440 4040 4460 4080
rect 4500 4040 4520 4080
rect 4440 3980 4520 4040
rect 4440 3940 4460 3980
rect 4500 3940 4520 3980
rect 4440 3910 4520 3940
rect 4770 4280 4850 4310
rect 4770 4240 4790 4280
rect 4830 4240 4850 4280
rect 4770 4180 4850 4240
rect 4770 4140 4790 4180
rect 4830 4140 4850 4180
rect 4770 4080 4850 4140
rect 4770 4040 4790 4080
rect 4830 4040 4850 4080
rect 4770 3980 4850 4040
rect 4770 3940 4790 3980
rect 4830 3940 4850 3980
rect 4770 3910 4850 3940
rect 5170 4280 5270 4310
rect 5170 4240 5200 4280
rect 5240 4240 5270 4280
rect 5170 4180 5270 4240
rect 5170 4140 5200 4180
rect 5240 4140 5270 4180
rect 5170 4080 5270 4140
rect 5170 4040 5200 4080
rect 5240 4040 5270 4080
rect 5170 3980 5270 4040
rect 5170 3940 5200 3980
rect 5240 3940 5270 3980
rect 5170 3910 5270 3940
rect 5560 4280 5660 4310
rect 5560 4240 5590 4280
rect 5630 4240 5660 4280
rect 5560 4180 5660 4240
rect 5560 4140 5590 4180
rect 5630 4140 5660 4180
rect 5560 4080 5660 4140
rect 5560 4040 5590 4080
rect 5630 4040 5660 4080
rect 5560 3980 5660 4040
rect 5560 3940 5590 3980
rect 5630 3940 5660 3980
rect 5560 3910 5660 3940
rect 5950 4280 6050 4310
rect 5950 4240 5980 4280
rect 6020 4240 6050 4280
rect 5950 4180 6050 4240
rect 5950 4140 5980 4180
rect 6020 4140 6050 4180
rect 5950 4080 6050 4140
rect 5950 4040 5980 4080
rect 6020 4040 6050 4080
rect 5950 3980 6050 4040
rect 5950 3940 5980 3980
rect 6020 3940 6050 3980
rect 5950 3910 6050 3940
rect 6630 4280 6730 4310
rect 6630 4240 6660 4280
rect 6700 4240 6730 4280
rect 6630 4180 6730 4240
rect 6630 4140 6660 4180
rect 6700 4140 6730 4180
rect 6630 4080 6730 4140
rect 6630 4040 6660 4080
rect 6700 4040 6730 4080
rect 6630 3980 6730 4040
rect 6630 3940 6660 3980
rect 6700 3940 6730 3980
rect 6630 3910 6730 3940
rect 8040 4290 8070 4330
rect 8110 4290 8140 4330
rect 8040 4230 8140 4290
rect 8040 4190 8070 4230
rect 8110 4190 8140 4230
rect 8040 4130 8140 4190
rect 8040 4090 8070 4130
rect 8110 4090 8140 4130
rect 8040 4030 8140 4090
rect 8040 3990 8070 4030
rect 8110 3990 8140 4030
rect 8040 3960 8140 3990
rect 9560 4330 9660 4360
rect 9560 4290 9590 4330
rect 9630 4290 9660 4330
rect 9560 4230 9660 4290
rect 9560 4190 9590 4230
rect 9630 4190 9660 4230
rect 9560 4130 9660 4190
rect 9560 4090 9590 4130
rect 9630 4090 9660 4130
rect 9560 4030 9660 4090
rect 9560 3990 9590 4030
rect 9630 3990 9660 4030
rect 9560 3960 9660 3990
rect 11080 4330 11180 4360
rect 11080 4290 11110 4330
rect 11150 4290 11180 4330
rect 11080 4230 11180 4290
rect 11080 4190 11110 4230
rect 11150 4190 11180 4230
rect 11080 4130 11180 4190
rect 11080 4090 11110 4130
rect 11150 4090 11180 4130
rect 11080 4030 11180 4090
rect 11080 3990 11110 4030
rect 11150 3990 11180 4030
rect 11080 3960 11180 3990
rect 2060 3520 2140 3550
rect 2060 3480 2080 3520
rect 2120 3480 2140 3520
rect 2060 3420 2140 3480
rect 2060 3380 2080 3420
rect 2120 3380 2140 3420
rect 2060 3320 2140 3380
rect 2060 3280 2080 3320
rect 2120 3280 2140 3320
rect 2060 3220 2140 3280
rect 2060 3180 2080 3220
rect 2120 3180 2140 3220
rect 2060 3150 2140 3180
rect 2960 3520 3040 3550
rect 2960 3480 2980 3520
rect 3020 3480 3040 3520
rect 2960 3420 3040 3480
rect 2960 3380 2980 3420
rect 3020 3380 3040 3420
rect 2960 3320 3040 3380
rect 2960 3280 2980 3320
rect 3020 3280 3040 3320
rect 2960 3220 3040 3280
rect 2960 3180 2980 3220
rect 3020 3180 3040 3220
rect 2960 3150 3040 3180
rect 3860 3520 3940 3550
rect 3860 3480 3880 3520
rect 3920 3480 3940 3520
rect 3860 3420 3940 3480
rect 3860 3380 3880 3420
rect 3920 3380 3940 3420
rect 3860 3320 3940 3380
rect 3860 3280 3880 3320
rect 3920 3280 3940 3320
rect 3860 3220 3940 3280
rect 3860 3180 3880 3220
rect 3920 3180 3940 3220
rect 3860 3150 3940 3180
rect 4260 3520 4340 3550
rect 4260 3480 4280 3520
rect 4320 3480 4340 3520
rect 4260 3420 4340 3480
rect 4260 3380 4280 3420
rect 4320 3380 4340 3420
rect 4260 3320 4340 3380
rect 4260 3280 4280 3320
rect 4320 3280 4340 3320
rect 4260 3220 4340 3280
rect 4260 3180 4280 3220
rect 4320 3180 4340 3220
rect 4260 3150 4340 3180
rect 4590 3520 4670 3550
rect 4590 3480 4610 3520
rect 4650 3480 4670 3520
rect 4590 3420 4670 3480
rect 4590 3380 4610 3420
rect 4650 3380 4670 3420
rect 4590 3320 4670 3380
rect 4590 3280 4610 3320
rect 4650 3280 4670 3320
rect 4590 3220 4670 3280
rect 4590 3180 4610 3220
rect 4650 3180 4670 3220
rect 4590 3150 4670 3180
rect 4920 3520 5000 3550
rect 4920 3480 4940 3520
rect 4980 3480 5000 3520
rect 4920 3420 5000 3480
rect 4920 3380 4940 3420
rect 4980 3380 5000 3420
rect 4920 3320 5000 3380
rect 4920 3280 4940 3320
rect 4980 3280 5000 3320
rect 4920 3220 5000 3280
rect 4920 3180 4940 3220
rect 4980 3180 5000 3220
rect 4920 3150 5000 3180
rect 5170 3520 5270 3550
rect 5170 3480 5200 3520
rect 5240 3480 5270 3520
rect 5170 3420 5270 3480
rect 5170 3380 5200 3420
rect 5240 3380 5270 3420
rect 5170 3320 5270 3380
rect 5170 3280 5200 3320
rect 5240 3280 5270 3320
rect 5170 3220 5270 3280
rect 5170 3180 5200 3220
rect 5240 3180 5270 3220
rect 5170 3150 5270 3180
rect 5950 3520 6050 3550
rect 5950 3480 5980 3520
rect 6020 3480 6050 3520
rect 5950 3420 6050 3480
rect 5950 3380 5980 3420
rect 6020 3380 6050 3420
rect 5950 3320 6050 3380
rect 5950 3280 5980 3320
rect 6020 3280 6050 3320
rect 5950 3220 6050 3280
rect 5950 3180 5980 3220
rect 6020 3180 6050 3220
rect 5950 3150 6050 3180
rect 2180 1090 2260 1120
rect 2180 1050 2200 1090
rect 2240 1050 2260 1090
rect 2180 1020 2260 1050
rect 4550 1090 4630 1120
rect 4550 1050 4570 1090
rect 4610 1050 4630 1090
rect 4550 1020 4630 1050
rect 7420 1090 7500 1120
rect 7420 1050 7440 1090
rect 7480 1050 7500 1090
rect 7420 1020 7500 1050
rect 8720 1090 8800 1120
rect 8720 1050 8740 1090
rect 8780 1050 8800 1090
rect 8720 1020 8800 1050
rect 10020 1090 10100 1120
rect 10020 1050 10040 1090
rect 10080 1050 10100 1090
rect 10020 1020 10100 1050
rect 11320 1090 11400 1120
rect 11320 1050 11340 1090
rect 11380 1050 11400 1090
rect 11320 1020 11400 1050
rect 12590 850 12670 880
rect 12590 810 12610 850
rect 12650 810 12670 850
rect 12590 750 12670 810
rect 12590 710 12610 750
rect 12650 710 12670 750
rect 12590 680 12670 710
rect 13190 850 13270 880
rect 13190 810 13210 850
rect 13250 810 13270 850
rect 13190 750 13270 810
rect 13190 710 13210 750
rect 13250 710 13270 750
rect 13190 680 13270 710
rect 13790 850 13870 880
rect 13790 810 13810 850
rect 13850 810 13870 850
rect 13790 750 13870 810
rect 13790 710 13810 750
rect 13850 710 13870 750
rect 13790 680 13870 710
rect 12860 500 12940 530
rect 12860 460 12880 500
rect 12920 460 12940 500
rect 12860 400 12940 460
rect 12860 360 12880 400
rect 12920 360 12940 400
rect 12860 300 12940 360
rect 12860 260 12880 300
rect 12920 260 12940 300
rect 12860 200 12940 260
rect 12860 160 12880 200
rect 12920 160 12940 200
rect 12860 130 12940 160
rect 13460 500 13540 530
rect 13460 460 13480 500
rect 13520 460 13540 500
rect 13460 400 13540 460
rect 13460 360 13480 400
rect 13520 360 13540 400
rect 13460 300 13540 360
rect 13460 260 13480 300
rect 13520 260 13540 300
rect 13460 200 13540 260
rect 13460 160 13480 200
rect 13520 160 13540 200
rect 13460 130 13540 160
rect 14060 500 14140 530
rect 14060 460 14080 500
rect 14120 460 14140 500
rect 14060 400 14140 460
rect 14060 360 14080 400
rect 14120 360 14140 400
rect 14060 300 14140 360
rect 14060 260 14080 300
rect 14120 260 14140 300
rect 14060 200 14140 260
rect 14060 160 14080 200
rect 14120 160 14140 200
rect 14060 130 14140 160
<< psubdiffcont >>
rect 3250 15040 3290 15080
rect 3250 14960 3290 15000
rect 3250 14880 3290 14920
rect 1400 14728 1434 14762
rect 1490 14728 1524 14762
rect 1580 14728 1614 14762
rect 1670 14728 1704 14762
rect 1760 14728 1794 14762
rect 1850 14728 1884 14762
rect 1940 14728 1974 14762
rect 2030 14728 2064 14762
rect 2120 14728 2154 14762
rect 2210 14728 2244 14762
rect 2300 14728 2334 14762
rect 2390 14728 2424 14762
rect 1299 14644 1333 14678
rect 2486 14644 2520 14678
rect 1299 14554 1333 14588
rect 1299 14464 1333 14498
rect 1299 14374 1333 14408
rect 1299 14284 1333 14318
rect 1299 14194 1333 14228
rect 1299 14104 1333 14138
rect 1299 14014 1333 14048
rect 1299 13924 1333 13958
rect 1299 13834 1333 13868
rect 1299 13744 1333 13778
rect 1299 13654 1333 13688
rect 2486 14554 2520 14588
rect 2486 14464 2520 14498
rect 2486 14374 2520 14408
rect 2486 14284 2520 14318
rect 2486 14194 2520 14228
rect 2486 14104 2520 14138
rect 2486 14014 2520 14048
rect 2486 13924 2520 13958
rect 2486 13834 2520 13868
rect 2486 13744 2520 13778
rect 2486 13654 2520 13688
rect 1299 13564 1333 13598
rect 1400 13541 1434 13575
rect 1490 13541 1524 13575
rect 1580 13541 1614 13575
rect 1670 13541 1704 13575
rect 1760 13541 1794 13575
rect 1850 13541 1884 13575
rect 1940 13541 1974 13575
rect 2030 13541 2064 13575
rect 2120 13541 2154 13575
rect 2210 13541 2244 13575
rect 2300 13541 2334 13575
rect 2390 13541 2424 13575
rect 2486 13564 2520 13598
rect 2760 14728 2794 14762
rect 2850 14728 2884 14762
rect 2940 14728 2974 14762
rect 3030 14728 3064 14762
rect 3120 14728 3154 14762
rect 3210 14728 3244 14762
rect 3300 14728 3334 14762
rect 3390 14728 3424 14762
rect 3480 14728 3514 14762
rect 3570 14728 3604 14762
rect 3660 14728 3694 14762
rect 3750 14728 3784 14762
rect 2659 14644 2693 14678
rect 3846 14644 3880 14678
rect 2659 14554 2693 14588
rect 2659 14464 2693 14498
rect 2659 14374 2693 14408
rect 2659 14284 2693 14318
rect 2659 14194 2693 14228
rect 2659 14104 2693 14138
rect 2659 14014 2693 14048
rect 2659 13924 2693 13958
rect 2659 13834 2693 13868
rect 2659 13744 2693 13778
rect 2659 13654 2693 13688
rect 3846 14554 3880 14588
rect 3846 14464 3880 14498
rect 3846 14374 3880 14408
rect 3846 14284 3880 14318
rect 3846 14194 3880 14228
rect 3846 14104 3880 14138
rect 3846 14014 3880 14048
rect 3846 13924 3880 13958
rect 3846 13834 3880 13868
rect 3846 13744 3880 13778
rect 3846 13654 3880 13688
rect 2659 13564 2693 13598
rect 2760 13541 2794 13575
rect 2850 13541 2884 13575
rect 2940 13541 2974 13575
rect 3030 13541 3064 13575
rect 3120 13541 3154 13575
rect 3210 13541 3244 13575
rect 3300 13541 3334 13575
rect 3390 13541 3424 13575
rect 3480 13541 3514 13575
rect 3570 13541 3604 13575
rect 3660 13541 3694 13575
rect 3750 13541 3784 13575
rect 3846 13564 3880 13598
rect 4120 14728 4154 14762
rect 4210 14728 4244 14762
rect 4300 14728 4334 14762
rect 4390 14728 4424 14762
rect 4480 14728 4514 14762
rect 4570 14728 4604 14762
rect 4660 14728 4694 14762
rect 4750 14728 4784 14762
rect 4840 14728 4874 14762
rect 4930 14728 4964 14762
rect 5020 14728 5054 14762
rect 5110 14728 5144 14762
rect 4019 14644 4053 14678
rect 5206 14644 5240 14678
rect 4019 14554 4053 14588
rect 4019 14464 4053 14498
rect 4019 14374 4053 14408
rect 4019 14284 4053 14318
rect 4019 14194 4053 14228
rect 4019 14104 4053 14138
rect 4019 14014 4053 14048
rect 4019 13924 4053 13958
rect 4019 13834 4053 13868
rect 4019 13744 4053 13778
rect 4019 13654 4053 13688
rect 5206 14554 5240 14588
rect 5206 14464 5240 14498
rect 5206 14374 5240 14408
rect 5206 14284 5240 14318
rect 5206 14194 5240 14228
rect 5206 14104 5240 14138
rect 5206 14014 5240 14048
rect 5206 13924 5240 13958
rect 5206 13834 5240 13868
rect 5206 13744 5240 13778
rect 5206 13654 5240 13688
rect 4019 13564 4053 13598
rect 4120 13541 4154 13575
rect 4210 13541 4244 13575
rect 4300 13541 4334 13575
rect 4390 13541 4424 13575
rect 4480 13541 4514 13575
rect 4570 13541 4604 13575
rect 4660 13541 4694 13575
rect 4750 13541 4784 13575
rect 4840 13541 4874 13575
rect 4930 13541 4964 13575
rect 5020 13541 5054 13575
rect 5110 13541 5144 13575
rect 5206 13564 5240 13598
rect 1400 13368 1434 13402
rect 1490 13368 1524 13402
rect 1580 13368 1614 13402
rect 1670 13368 1704 13402
rect 1760 13368 1794 13402
rect 1850 13368 1884 13402
rect 1940 13368 1974 13402
rect 2030 13368 2064 13402
rect 2120 13368 2154 13402
rect 2210 13368 2244 13402
rect 2300 13368 2334 13402
rect 2390 13368 2424 13402
rect 1299 13284 1333 13318
rect 2486 13284 2520 13318
rect 1299 13194 1333 13228
rect 1299 13104 1333 13138
rect 1299 13014 1333 13048
rect 1299 12924 1333 12958
rect 1299 12834 1333 12868
rect 1299 12744 1333 12778
rect 1299 12654 1333 12688
rect 1299 12564 1333 12598
rect 1299 12474 1333 12508
rect 1299 12384 1333 12418
rect 1299 12294 1333 12328
rect 2486 13194 2520 13228
rect 2486 13104 2520 13138
rect 2486 13014 2520 13048
rect 2486 12924 2520 12958
rect 2486 12834 2520 12868
rect 2486 12744 2520 12778
rect 2486 12654 2520 12688
rect 2486 12564 2520 12598
rect 2486 12474 2520 12508
rect 2486 12384 2520 12418
rect 2486 12294 2520 12328
rect 1299 12204 1333 12238
rect 1400 12181 1434 12215
rect 1490 12181 1524 12215
rect 1580 12181 1614 12215
rect 1670 12181 1704 12215
rect 1760 12181 1794 12215
rect 1850 12181 1884 12215
rect 1940 12181 1974 12215
rect 2030 12181 2064 12215
rect 2120 12181 2154 12215
rect 2210 12181 2244 12215
rect 2300 12181 2334 12215
rect 2390 12181 2424 12215
rect 2486 12204 2520 12238
rect 2760 13368 2794 13402
rect 2850 13368 2884 13402
rect 2940 13368 2974 13402
rect 3030 13368 3064 13402
rect 3120 13368 3154 13402
rect 3210 13368 3244 13402
rect 3300 13368 3334 13402
rect 3390 13368 3424 13402
rect 3480 13368 3514 13402
rect 3570 13368 3604 13402
rect 3660 13368 3694 13402
rect 3750 13368 3784 13402
rect 2659 13284 2693 13318
rect 3846 13284 3880 13318
rect 2659 13194 2693 13228
rect 2659 13104 2693 13138
rect 2659 13014 2693 13048
rect 2659 12924 2693 12958
rect 2659 12834 2693 12868
rect 2659 12744 2693 12778
rect 2659 12654 2693 12688
rect 2659 12564 2693 12598
rect 2659 12474 2693 12508
rect 2659 12384 2693 12418
rect 2659 12294 2693 12328
rect 3846 13194 3880 13228
rect 3846 13104 3880 13138
rect 3846 13014 3880 13048
rect 3846 12924 3880 12958
rect 3846 12834 3880 12868
rect 3846 12744 3880 12778
rect 3846 12654 3880 12688
rect 3846 12564 3880 12598
rect 3846 12474 3880 12508
rect 3846 12384 3880 12418
rect 3846 12294 3880 12328
rect 2659 12204 2693 12238
rect 2760 12181 2794 12215
rect 2850 12181 2884 12215
rect 2940 12181 2974 12215
rect 3030 12181 3064 12215
rect 3120 12181 3154 12215
rect 3210 12181 3244 12215
rect 3300 12181 3334 12215
rect 3390 12181 3424 12215
rect 3480 12181 3514 12215
rect 3570 12181 3604 12215
rect 3660 12181 3694 12215
rect 3750 12181 3784 12215
rect 3846 12204 3880 12238
rect 4120 13368 4154 13402
rect 4210 13368 4244 13402
rect 4300 13368 4334 13402
rect 4390 13368 4424 13402
rect 4480 13368 4514 13402
rect 4570 13368 4604 13402
rect 4660 13368 4694 13402
rect 4750 13368 4784 13402
rect 4840 13368 4874 13402
rect 4930 13368 4964 13402
rect 5020 13368 5054 13402
rect 5110 13368 5144 13402
rect 4019 13284 4053 13318
rect 5206 13284 5240 13318
rect 4019 13194 4053 13228
rect 4019 13104 4053 13138
rect 4019 13014 4053 13048
rect 4019 12924 4053 12958
rect 4019 12834 4053 12868
rect 4019 12744 4053 12778
rect 4019 12654 4053 12688
rect 4019 12564 4053 12598
rect 4019 12474 4053 12508
rect 4019 12384 4053 12418
rect 4019 12294 4053 12328
rect 5206 13194 5240 13228
rect 5206 13104 5240 13138
rect 5206 13014 5240 13048
rect 5206 12924 5240 12958
rect 5206 12834 5240 12868
rect 5206 12744 5240 12778
rect 5206 12654 5240 12688
rect 5206 12564 5240 12598
rect 5206 12474 5240 12508
rect 5206 12384 5240 12418
rect 5206 12294 5240 12328
rect 4019 12204 4053 12238
rect 4120 12181 4154 12215
rect 4210 12181 4244 12215
rect 4300 12181 4334 12215
rect 4390 12181 4424 12215
rect 4480 12181 4514 12215
rect 4570 12181 4604 12215
rect 4660 12181 4694 12215
rect 4750 12181 4784 12215
rect 4840 12181 4874 12215
rect 4930 12181 4964 12215
rect 5020 12181 5054 12215
rect 5110 12181 5144 12215
rect 5206 12204 5240 12238
rect 1400 12008 1434 12042
rect 1490 12008 1524 12042
rect 1580 12008 1614 12042
rect 1670 12008 1704 12042
rect 1760 12008 1794 12042
rect 1850 12008 1884 12042
rect 1940 12008 1974 12042
rect 2030 12008 2064 12042
rect 2120 12008 2154 12042
rect 2210 12008 2244 12042
rect 2300 12008 2334 12042
rect 2390 12008 2424 12042
rect 1299 11924 1333 11958
rect 2486 11924 2520 11958
rect 1299 11834 1333 11868
rect 1299 11744 1333 11778
rect 1299 11654 1333 11688
rect 1299 11564 1333 11598
rect 1299 11474 1333 11508
rect 1299 11384 1333 11418
rect 1299 11294 1333 11328
rect 1299 11204 1333 11238
rect 1299 11114 1333 11148
rect 1299 11024 1333 11058
rect 1299 10934 1333 10968
rect 2486 11834 2520 11868
rect 2486 11744 2520 11778
rect 2486 11654 2520 11688
rect 2486 11564 2520 11598
rect 2486 11474 2520 11508
rect 2486 11384 2520 11418
rect 2486 11294 2520 11328
rect 2486 11204 2520 11238
rect 2486 11114 2520 11148
rect 2486 11024 2520 11058
rect 2486 10934 2520 10968
rect 1299 10844 1333 10878
rect 1400 10821 1434 10855
rect 1490 10821 1524 10855
rect 1580 10821 1614 10855
rect 1670 10821 1704 10855
rect 1760 10821 1794 10855
rect 1850 10821 1884 10855
rect 1940 10821 1974 10855
rect 2030 10821 2064 10855
rect 2120 10821 2154 10855
rect 2210 10821 2244 10855
rect 2300 10821 2334 10855
rect 2390 10821 2424 10855
rect 2486 10844 2520 10878
rect 2760 12008 2794 12042
rect 2850 12008 2884 12042
rect 2940 12008 2974 12042
rect 3030 12008 3064 12042
rect 3120 12008 3154 12042
rect 3210 12008 3244 12042
rect 3300 12008 3334 12042
rect 3390 12008 3424 12042
rect 3480 12008 3514 12042
rect 3570 12008 3604 12042
rect 3660 12008 3694 12042
rect 3750 12008 3784 12042
rect 2659 11924 2693 11958
rect 3846 11924 3880 11958
rect 2659 11834 2693 11868
rect 2659 11744 2693 11778
rect 2659 11654 2693 11688
rect 2659 11564 2693 11598
rect 2659 11474 2693 11508
rect 2659 11384 2693 11418
rect 2659 11294 2693 11328
rect 2659 11204 2693 11238
rect 2659 11114 2693 11148
rect 2659 11024 2693 11058
rect 2659 10934 2693 10968
rect 3846 11834 3880 11868
rect 3846 11744 3880 11778
rect 3846 11654 3880 11688
rect 3846 11564 3880 11598
rect 3846 11474 3880 11508
rect 3846 11384 3880 11418
rect 3846 11294 3880 11328
rect 3846 11204 3880 11238
rect 3846 11114 3880 11148
rect 3846 11024 3880 11058
rect 3846 10934 3880 10968
rect 2659 10844 2693 10878
rect 2760 10821 2794 10855
rect 2850 10821 2884 10855
rect 2940 10821 2974 10855
rect 3030 10821 3064 10855
rect 3120 10821 3154 10855
rect 3210 10821 3244 10855
rect 3300 10821 3334 10855
rect 3390 10821 3424 10855
rect 3480 10821 3514 10855
rect 3570 10821 3604 10855
rect 3660 10821 3694 10855
rect 3750 10821 3784 10855
rect 3846 10844 3880 10878
rect 4120 12008 4154 12042
rect 4210 12008 4244 12042
rect 4300 12008 4334 12042
rect 4390 12008 4424 12042
rect 4480 12008 4514 12042
rect 4570 12008 4604 12042
rect 4660 12008 4694 12042
rect 4750 12008 4784 12042
rect 4840 12008 4874 12042
rect 4930 12008 4964 12042
rect 5020 12008 5054 12042
rect 5110 12008 5144 12042
rect 4019 11924 4053 11958
rect 5206 11924 5240 11958
rect 4019 11834 4053 11868
rect 4019 11744 4053 11778
rect 4019 11654 4053 11688
rect 4019 11564 4053 11598
rect 4019 11474 4053 11508
rect 4019 11384 4053 11418
rect 4019 11294 4053 11328
rect 4019 11204 4053 11238
rect 4019 11114 4053 11148
rect 4019 11024 4053 11058
rect 4019 10934 4053 10968
rect 5206 11834 5240 11868
rect 5206 11744 5240 11778
rect 5206 11654 5240 11688
rect 5206 11564 5240 11598
rect 5206 11474 5240 11508
rect 5206 11384 5240 11418
rect 5206 11294 5240 11328
rect 5206 11204 5240 11238
rect 5206 11114 5240 11148
rect 5206 11024 5240 11058
rect 5206 10934 5240 10968
rect 4019 10844 4053 10878
rect 4120 10821 4154 10855
rect 4210 10821 4244 10855
rect 4300 10821 4334 10855
rect 4390 10821 4424 10855
rect 4480 10821 4514 10855
rect 4570 10821 4604 10855
rect 4660 10821 4694 10855
rect 4750 10821 4784 10855
rect 4840 10821 4874 10855
rect 4930 10821 4964 10855
rect 5020 10821 5054 10855
rect 5110 10821 5144 10855
rect 5206 10844 5240 10878
rect 5410 10220 5450 10260
rect 5410 10120 5450 10160
rect 1910 9610 1950 9650
rect 1910 9510 1950 9550
rect 1910 9410 1950 9450
rect 1910 9310 1950 9350
rect 1910 9210 1950 9250
rect 4590 9610 4630 9650
rect 4590 9510 4630 9550
rect 4590 9410 4630 9450
rect 4590 9310 4630 9350
rect 4590 9210 4630 9250
rect 2810 8690 2850 8730
rect 2810 8610 2850 8650
rect 2810 8530 2850 8570
rect 3690 8690 3730 8730
rect 3690 8610 3730 8650
rect 3690 8530 3730 8570
rect 8130 8530 8170 8580
rect 8130 8390 8170 8440
rect 10330 8530 10370 8580
rect 10330 8390 10370 8440
rect 8180 7850 8220 7890
rect 9160 7850 9200 7890
rect 10460 7850 10500 7890
rect 11440 7850 11480 7890
rect 2080 4660 2120 4700
rect 2080 4560 2120 4600
rect 2980 4660 3020 4700
rect 2980 4560 3020 4600
rect 3880 4660 3920 4700
rect 3880 4560 3920 4600
rect 4020 4660 4060 4700
rect 4020 4560 4060 4600
rect 4460 4660 4500 4700
rect 4460 4560 4500 4600
rect 4790 4660 4830 4700
rect 4790 4560 4830 4600
rect 5210 4660 5250 4700
rect 5210 4560 5250 4600
rect 5600 4660 5640 4700
rect 5600 4560 5640 4600
rect 5990 4660 6030 4700
rect 5990 4560 6030 4600
rect 7870 3310 7910 3350
rect 7870 3210 7910 3250
rect 7870 3110 7910 3150
rect 7870 3010 7910 3050
rect 8950 3310 8990 3350
rect 8950 3210 8990 3250
rect 8950 3110 8990 3150
rect 8950 3010 8990 3050
rect 10030 3310 10070 3350
rect 10030 3210 10070 3250
rect 10030 3110 10070 3150
rect 10030 3010 10070 3050
rect 11110 3310 11150 3350
rect 11110 3210 11150 3250
rect 11110 3110 11150 3150
rect 11110 3010 11150 3050
rect 2080 2860 2120 2900
rect 2080 2760 2120 2800
rect 2980 2860 3020 2900
rect 2980 2760 3020 2800
rect 3880 2860 3920 2900
rect 3880 2760 3920 2800
rect 4280 2860 4320 2900
rect 4280 2760 4320 2800
rect 4610 2860 4650 2900
rect 4610 2760 4650 2800
rect 4940 2860 4980 2900
rect 4940 2760 4980 2800
rect 5200 2860 5240 2900
rect 5200 2760 5240 2800
rect 5980 2860 6020 2900
rect 5980 2760 6020 2800
rect 6660 2860 6700 2900
rect 6660 2760 6700 2800
rect 17380 2610 17420 2650
rect 12610 1930 12650 1970
rect 12610 1830 12650 1870
rect 13210 1930 13250 1970
rect 13210 1830 13250 1870
rect 13810 1930 13850 1970
rect 13810 1830 13850 1870
rect 12610 1600 12650 1640
rect 13210 1600 13250 1640
rect 13810 1600 13850 1640
rect 8340 1460 8380 1500
rect 5100 1370 5140 1410
rect 6550 1370 6590 1410
rect 9640 1460 9680 1500
rect 10940 1460 10980 1500
<< nsubdiffcont >>
rect 1540 14578 1574 14612
rect 1630 14578 1664 14612
rect 1720 14578 1754 14612
rect 1810 14578 1844 14612
rect 1900 14578 1934 14612
rect 1990 14578 2024 14612
rect 2080 14578 2114 14612
rect 2170 14578 2204 14612
rect 2260 14578 2294 14612
rect 1448 14484 1482 14518
rect 1448 14394 1482 14428
rect 1448 14304 1482 14338
rect 1448 14214 1482 14248
rect 1448 14124 1482 14158
rect 1448 14034 1482 14068
rect 1448 13944 1482 13978
rect 1448 13854 1482 13888
rect 2338 14465 2372 14499
rect 2338 14375 2372 14409
rect 2338 14285 2372 14319
rect 2338 14195 2372 14229
rect 2338 14105 2372 14139
rect 2338 14015 2372 14049
rect 2338 13925 2372 13959
rect 2338 13835 2372 13869
rect 1448 13764 1482 13798
rect 2338 13745 2372 13779
rect 1506 13688 1540 13722
rect 1596 13688 1630 13722
rect 1686 13688 1720 13722
rect 1776 13688 1810 13722
rect 1866 13688 1900 13722
rect 1956 13688 1990 13722
rect 2046 13688 2080 13722
rect 2136 13688 2170 13722
rect 2226 13688 2260 13722
rect 2900 14578 2934 14612
rect 2990 14578 3024 14612
rect 3080 14578 3114 14612
rect 3170 14578 3204 14612
rect 3260 14578 3294 14612
rect 3350 14578 3384 14612
rect 3440 14578 3474 14612
rect 3530 14578 3564 14612
rect 3620 14578 3654 14612
rect 2808 14484 2842 14518
rect 2808 14394 2842 14428
rect 2808 14304 2842 14338
rect 2808 14214 2842 14248
rect 2808 14124 2842 14158
rect 2808 14034 2842 14068
rect 2808 13944 2842 13978
rect 2808 13854 2842 13888
rect 3698 14465 3732 14499
rect 3698 14375 3732 14409
rect 3698 14285 3732 14319
rect 3698 14195 3732 14229
rect 3698 14105 3732 14139
rect 3698 14015 3732 14049
rect 3698 13925 3732 13959
rect 3698 13835 3732 13869
rect 2808 13764 2842 13798
rect 3698 13745 3732 13779
rect 2866 13688 2900 13722
rect 2956 13688 2990 13722
rect 3046 13688 3080 13722
rect 3136 13688 3170 13722
rect 3226 13688 3260 13722
rect 3316 13688 3350 13722
rect 3406 13688 3440 13722
rect 3496 13688 3530 13722
rect 3586 13688 3620 13722
rect 4260 14578 4294 14612
rect 4350 14578 4384 14612
rect 4440 14578 4474 14612
rect 4530 14578 4564 14612
rect 4620 14578 4654 14612
rect 4710 14578 4744 14612
rect 4800 14578 4834 14612
rect 4890 14578 4924 14612
rect 4980 14578 5014 14612
rect 4168 14484 4202 14518
rect 4168 14394 4202 14428
rect 4168 14304 4202 14338
rect 4168 14214 4202 14248
rect 4168 14124 4202 14158
rect 4168 14034 4202 14068
rect 4168 13944 4202 13978
rect 4168 13854 4202 13888
rect 5058 14465 5092 14499
rect 5058 14375 5092 14409
rect 5058 14285 5092 14319
rect 5058 14195 5092 14229
rect 5058 14105 5092 14139
rect 5058 14015 5092 14049
rect 5058 13925 5092 13959
rect 5058 13835 5092 13869
rect 4168 13764 4202 13798
rect 5058 13745 5092 13779
rect 4226 13688 4260 13722
rect 4316 13688 4350 13722
rect 4406 13688 4440 13722
rect 4496 13688 4530 13722
rect 4586 13688 4620 13722
rect 4676 13688 4710 13722
rect 4766 13688 4800 13722
rect 4856 13688 4890 13722
rect 4946 13688 4980 13722
rect 1540 13218 1574 13252
rect 1630 13218 1664 13252
rect 1720 13218 1754 13252
rect 1810 13218 1844 13252
rect 1900 13218 1934 13252
rect 1990 13218 2024 13252
rect 2080 13218 2114 13252
rect 2170 13218 2204 13252
rect 2260 13218 2294 13252
rect 1448 13124 1482 13158
rect 1448 13034 1482 13068
rect 1448 12944 1482 12978
rect 1448 12854 1482 12888
rect 1448 12764 1482 12798
rect 1448 12674 1482 12708
rect 1448 12584 1482 12618
rect 1448 12494 1482 12528
rect 2338 13105 2372 13139
rect 2338 13015 2372 13049
rect 2338 12925 2372 12959
rect 2338 12835 2372 12869
rect 2338 12745 2372 12779
rect 2338 12655 2372 12689
rect 2338 12565 2372 12599
rect 2338 12475 2372 12509
rect 1448 12404 1482 12438
rect 2338 12385 2372 12419
rect 1506 12328 1540 12362
rect 1596 12328 1630 12362
rect 1686 12328 1720 12362
rect 1776 12328 1810 12362
rect 1866 12328 1900 12362
rect 1956 12328 1990 12362
rect 2046 12328 2080 12362
rect 2136 12328 2170 12362
rect 2226 12328 2260 12362
rect 2900 13218 2934 13252
rect 2990 13218 3024 13252
rect 3080 13218 3114 13252
rect 3170 13218 3204 13252
rect 3260 13218 3294 13252
rect 3350 13218 3384 13252
rect 3440 13218 3474 13252
rect 3530 13218 3564 13252
rect 3620 13218 3654 13252
rect 2808 13124 2842 13158
rect 2808 13034 2842 13068
rect 2808 12944 2842 12978
rect 2808 12854 2842 12888
rect 2808 12764 2842 12798
rect 2808 12674 2842 12708
rect 2808 12584 2842 12618
rect 2808 12494 2842 12528
rect 3698 13105 3732 13139
rect 3698 13015 3732 13049
rect 3698 12925 3732 12959
rect 3698 12835 3732 12869
rect 3698 12745 3732 12779
rect 3698 12655 3732 12689
rect 3698 12565 3732 12599
rect 3698 12475 3732 12509
rect 2808 12404 2842 12438
rect 3698 12385 3732 12419
rect 2866 12328 2900 12362
rect 2956 12328 2990 12362
rect 3046 12328 3080 12362
rect 3136 12328 3170 12362
rect 3226 12328 3260 12362
rect 3316 12328 3350 12362
rect 3406 12328 3440 12362
rect 3496 12328 3530 12362
rect 3586 12328 3620 12362
rect 4260 13218 4294 13252
rect 4350 13218 4384 13252
rect 4440 13218 4474 13252
rect 4530 13218 4564 13252
rect 4620 13218 4654 13252
rect 4710 13218 4744 13252
rect 4800 13218 4834 13252
rect 4890 13218 4924 13252
rect 4980 13218 5014 13252
rect 4168 13124 4202 13158
rect 4168 13034 4202 13068
rect 4168 12944 4202 12978
rect 4168 12854 4202 12888
rect 4168 12764 4202 12798
rect 4168 12674 4202 12708
rect 4168 12584 4202 12618
rect 4168 12494 4202 12528
rect 5058 13105 5092 13139
rect 5058 13015 5092 13049
rect 5058 12925 5092 12959
rect 5058 12835 5092 12869
rect 5058 12745 5092 12779
rect 5058 12655 5092 12689
rect 5058 12565 5092 12599
rect 5058 12475 5092 12509
rect 4168 12404 4202 12438
rect 5058 12385 5092 12419
rect 4226 12328 4260 12362
rect 4316 12328 4350 12362
rect 4406 12328 4440 12362
rect 4496 12328 4530 12362
rect 4586 12328 4620 12362
rect 4676 12328 4710 12362
rect 4766 12328 4800 12362
rect 4856 12328 4890 12362
rect 4946 12328 4980 12362
rect 1540 11858 1574 11892
rect 1630 11858 1664 11892
rect 1720 11858 1754 11892
rect 1810 11858 1844 11892
rect 1900 11858 1934 11892
rect 1990 11858 2024 11892
rect 2080 11858 2114 11892
rect 2170 11858 2204 11892
rect 2260 11858 2294 11892
rect 1448 11764 1482 11798
rect 1448 11674 1482 11708
rect 1448 11584 1482 11618
rect 1448 11494 1482 11528
rect 1448 11404 1482 11438
rect 1448 11314 1482 11348
rect 1448 11224 1482 11258
rect 1448 11134 1482 11168
rect 2338 11745 2372 11779
rect 2338 11655 2372 11689
rect 2338 11565 2372 11599
rect 2338 11475 2372 11509
rect 2338 11385 2372 11419
rect 2338 11295 2372 11329
rect 2338 11205 2372 11239
rect 2338 11115 2372 11149
rect 1448 11044 1482 11078
rect 2338 11025 2372 11059
rect 1506 10968 1540 11002
rect 1596 10968 1630 11002
rect 1686 10968 1720 11002
rect 1776 10968 1810 11002
rect 1866 10968 1900 11002
rect 1956 10968 1990 11002
rect 2046 10968 2080 11002
rect 2136 10968 2170 11002
rect 2226 10968 2260 11002
rect 2900 11858 2934 11892
rect 2990 11858 3024 11892
rect 3080 11858 3114 11892
rect 3170 11858 3204 11892
rect 3260 11858 3294 11892
rect 3350 11858 3384 11892
rect 3440 11858 3474 11892
rect 3530 11858 3564 11892
rect 3620 11858 3654 11892
rect 2808 11764 2842 11798
rect 2808 11674 2842 11708
rect 2808 11584 2842 11618
rect 2808 11494 2842 11528
rect 2808 11404 2842 11438
rect 2808 11314 2842 11348
rect 2808 11224 2842 11258
rect 2808 11134 2842 11168
rect 3698 11745 3732 11779
rect 3698 11655 3732 11689
rect 3698 11565 3732 11599
rect 3698 11475 3732 11509
rect 3698 11385 3732 11419
rect 3698 11295 3732 11329
rect 3698 11205 3732 11239
rect 3698 11115 3732 11149
rect 2808 11044 2842 11078
rect 3698 11025 3732 11059
rect 2866 10968 2900 11002
rect 2956 10968 2990 11002
rect 3046 10968 3080 11002
rect 3136 10968 3170 11002
rect 3226 10968 3260 11002
rect 3316 10968 3350 11002
rect 3406 10968 3440 11002
rect 3496 10968 3530 11002
rect 3586 10968 3620 11002
rect 4260 11858 4294 11892
rect 4350 11858 4384 11892
rect 4440 11858 4474 11892
rect 4530 11858 4564 11892
rect 4620 11858 4654 11892
rect 4710 11858 4744 11892
rect 4800 11858 4834 11892
rect 4890 11858 4924 11892
rect 4980 11858 5014 11892
rect 4168 11764 4202 11798
rect 4168 11674 4202 11708
rect 4168 11584 4202 11618
rect 4168 11494 4202 11528
rect 4168 11404 4202 11438
rect 4168 11314 4202 11348
rect 4168 11224 4202 11258
rect 4168 11134 4202 11168
rect 5058 11745 5092 11779
rect 5058 11655 5092 11689
rect 5058 11565 5092 11599
rect 5058 11475 5092 11509
rect 5058 11385 5092 11419
rect 5058 11295 5092 11329
rect 5058 11205 5092 11239
rect 5058 11115 5092 11149
rect 4168 11044 4202 11078
rect 5058 11025 5092 11059
rect 4226 10968 4260 11002
rect 4316 10968 4350 11002
rect 4406 10968 4440 11002
rect 4496 10968 4530 11002
rect 4586 10968 4620 11002
rect 4676 10968 4710 11002
rect 4766 10968 4800 11002
rect 4856 10968 4890 11002
rect 4946 10968 4980 11002
rect 450 7760 490 7800
rect 450 7660 490 7700
rect 3010 7760 3050 7800
rect 3010 7660 3050 7700
rect 3490 7760 3530 7800
rect 3490 7660 3530 7700
rect 6050 7760 6090 7800
rect 6050 7660 6090 7700
rect 9320 7280 9360 7320
rect 9320 7180 9360 7220
rect 10300 7280 10340 7320
rect 10300 7180 10340 7220
rect 10460 7280 10500 7320
rect 10460 7180 10500 7220
rect 11440 7280 11480 7320
rect 11440 7180 11480 7220
rect 1550 6600 1590 6640
rect 1550 6500 1590 6540
rect 1550 6400 1590 6440
rect 1550 6300 1590 6340
rect 1550 6200 1590 6240
rect 1550 6100 1590 6140
rect 4950 6600 4990 6640
rect 8250 6630 8290 6670
rect 4950 6500 4990 6540
rect 8250 6530 8290 6570
rect 4950 6400 4990 6440
rect 4950 6300 4990 6340
rect 5410 6400 5450 6440
rect 5410 6300 5450 6340
rect 6020 6400 6060 6440
rect 6020 6300 6060 6340
rect 8250 6430 8290 6470
rect 8250 6330 8290 6370
rect 4950 6200 4990 6240
rect 8250 6230 8290 6270
rect 10450 6630 10490 6670
rect 10450 6530 10490 6570
rect 10450 6430 10490 6470
rect 10450 6330 10490 6370
rect 10450 6230 10490 6270
rect 4950 6100 4990 6140
rect 1560 5600 1600 5640
rect 1560 5500 1600 5540
rect 3040 5600 3080 5640
rect 3040 5500 3080 5540
rect 3460 5600 3500 5640
rect 3460 5500 3500 5540
rect 4940 5600 4980 5640
rect 4940 5500 4980 5540
rect 2080 4240 2120 4280
rect 2080 4140 2120 4180
rect 2080 4040 2120 4080
rect 2080 3940 2120 3980
rect 2980 4240 3020 4280
rect 2980 4140 3020 4180
rect 2980 4040 3020 4080
rect 2980 3940 3020 3980
rect 3880 4240 3920 4280
rect 3880 4140 3920 4180
rect 3880 4040 3920 4080
rect 3880 3940 3920 3980
rect 4020 4240 4060 4280
rect 4020 4140 4060 4180
rect 4020 4040 4060 4080
rect 4020 3940 4060 3980
rect 4460 4240 4500 4280
rect 4460 4140 4500 4180
rect 4460 4040 4500 4080
rect 4460 3940 4500 3980
rect 4790 4240 4830 4280
rect 4790 4140 4830 4180
rect 4790 4040 4830 4080
rect 4790 3940 4830 3980
rect 5200 4240 5240 4280
rect 5200 4140 5240 4180
rect 5200 4040 5240 4080
rect 5200 3940 5240 3980
rect 5590 4240 5630 4280
rect 5590 4140 5630 4180
rect 5590 4040 5630 4080
rect 5590 3940 5630 3980
rect 5980 4240 6020 4280
rect 5980 4140 6020 4180
rect 5980 4040 6020 4080
rect 5980 3940 6020 3980
rect 6660 4240 6700 4280
rect 6660 4140 6700 4180
rect 6660 4040 6700 4080
rect 6660 3940 6700 3980
rect 8070 4290 8110 4330
rect 8070 4190 8110 4230
rect 8070 4090 8110 4130
rect 8070 3990 8110 4030
rect 9590 4290 9630 4330
rect 9590 4190 9630 4230
rect 9590 4090 9630 4130
rect 9590 3990 9630 4030
rect 11110 4290 11150 4330
rect 11110 4190 11150 4230
rect 11110 4090 11150 4130
rect 11110 3990 11150 4030
rect 2080 3480 2120 3520
rect 2080 3380 2120 3420
rect 2080 3280 2120 3320
rect 2080 3180 2120 3220
rect 2980 3480 3020 3520
rect 2980 3380 3020 3420
rect 2980 3280 3020 3320
rect 2980 3180 3020 3220
rect 3880 3480 3920 3520
rect 3880 3380 3920 3420
rect 3880 3280 3920 3320
rect 3880 3180 3920 3220
rect 4280 3480 4320 3520
rect 4280 3380 4320 3420
rect 4280 3280 4320 3320
rect 4280 3180 4320 3220
rect 4610 3480 4650 3520
rect 4610 3380 4650 3420
rect 4610 3280 4650 3320
rect 4610 3180 4650 3220
rect 4940 3480 4980 3520
rect 4940 3380 4980 3420
rect 4940 3280 4980 3320
rect 4940 3180 4980 3220
rect 5200 3480 5240 3520
rect 5200 3380 5240 3420
rect 5200 3280 5240 3320
rect 5200 3180 5240 3220
rect 5980 3480 6020 3520
rect 5980 3380 6020 3420
rect 5980 3280 6020 3320
rect 5980 3180 6020 3220
rect 2200 1050 2240 1090
rect 4570 1050 4610 1090
rect 7440 1050 7480 1090
rect 8740 1050 8780 1090
rect 10040 1050 10080 1090
rect 11340 1050 11380 1090
rect 12610 810 12650 850
rect 12610 710 12650 750
rect 13210 810 13250 850
rect 13210 710 13250 750
rect 13810 810 13850 850
rect 13810 710 13850 750
rect 12880 460 12920 500
rect 12880 360 12920 400
rect 12880 260 12920 300
rect 12880 160 12920 200
rect 13480 460 13520 500
rect 13480 360 13520 400
rect 13480 260 13520 300
rect 13480 160 13520 200
rect 14080 460 14120 500
rect 14080 360 14120 400
rect 14080 260 14120 300
rect 14080 160 14120 200
<< poly >>
rect 1230 10290 3230 10320
rect 3310 10290 5310 10320
rect 1230 10060 3230 10090
rect 3310 10060 5310 10090
rect 1310 10040 1390 10060
rect 1310 10000 1330 10040
rect 1370 10000 1390 10040
rect 1310 9980 1390 10000
rect 1470 10040 1550 10060
rect 1470 10000 1490 10040
rect 1530 10000 1550 10040
rect 1470 9980 1550 10000
rect 1630 10040 1710 10060
rect 1630 10000 1650 10040
rect 1690 10000 1710 10040
rect 1630 9980 1710 10000
rect 1790 10040 1870 10060
rect 1790 10000 1810 10040
rect 1850 10000 1870 10040
rect 1790 9980 1870 10000
rect 1950 10040 2030 10060
rect 1950 10000 1970 10040
rect 2010 10000 2030 10040
rect 1950 9980 2030 10000
rect 2110 10040 2190 10060
rect 2110 10000 2130 10040
rect 2170 10000 2190 10040
rect 2110 9980 2190 10000
rect 2270 10040 2350 10060
rect 2270 10000 2290 10040
rect 2330 10000 2350 10040
rect 2270 9980 2350 10000
rect 2430 10040 2510 10060
rect 2430 10000 2450 10040
rect 2490 10000 2510 10040
rect 2430 9980 2510 10000
rect 2590 10040 2670 10060
rect 2590 10000 2610 10040
rect 2650 10000 2670 10040
rect 2590 9980 2670 10000
rect 2750 10040 2830 10060
rect 2750 10000 2770 10040
rect 2810 10000 2830 10040
rect 2750 9980 2830 10000
rect 2910 10040 2990 10060
rect 2910 10000 2930 10040
rect 2970 10000 2990 10040
rect 2910 9980 2990 10000
rect 3070 10040 3150 10060
rect 3070 10000 3090 10040
rect 3130 10000 3150 10040
rect 3070 9980 3150 10000
rect 3390 10040 3470 10060
rect 3390 10000 3410 10040
rect 3450 10000 3470 10040
rect 3390 9980 3470 10000
rect 3550 10040 3630 10060
rect 3550 10000 3570 10040
rect 3610 10000 3630 10040
rect 3550 9980 3630 10000
rect 3710 10040 3790 10060
rect 3710 10000 3730 10040
rect 3770 10000 3790 10040
rect 3710 9980 3790 10000
rect 3870 10040 3950 10060
rect 3870 10000 3890 10040
rect 3930 10000 3950 10040
rect 3870 9980 3950 10000
rect 4030 10040 4110 10060
rect 4030 10000 4050 10040
rect 4090 10000 4110 10040
rect 4030 9980 4110 10000
rect 4190 10040 4270 10060
rect 4190 10000 4210 10040
rect 4250 10000 4270 10040
rect 4190 9980 4270 10000
rect 4350 10040 4430 10060
rect 4350 10000 4370 10040
rect 4410 10000 4430 10040
rect 4350 9980 4430 10000
rect 4510 10040 4590 10060
rect 4510 10000 4530 10040
rect 4570 10000 4590 10040
rect 4510 9980 4590 10000
rect 4670 10040 4750 10060
rect 4670 10000 4690 10040
rect 4730 10000 4750 10040
rect 4670 9980 4750 10000
rect 4830 10040 4910 10060
rect 4830 10000 4850 10040
rect 4890 10000 4910 10040
rect 4830 9980 4910 10000
rect 4990 10040 5070 10060
rect 4990 10000 5010 10040
rect 5050 10000 5070 10040
rect 4990 9980 5070 10000
rect 5150 10040 5230 10060
rect 5150 10000 5170 10040
rect 5210 10000 5230 10040
rect 5150 9980 5230 10000
rect 810 9680 1810 9710
rect 2050 9680 3050 9710
rect 3490 9680 4490 9710
rect 4730 9680 5730 9710
rect 810 9150 1810 9180
rect 2050 9150 3050 9180
rect 3490 9150 4490 9180
rect 4730 9150 5730 9180
rect 910 9130 990 9150
rect 910 9090 930 9130
rect 970 9090 990 9130
rect 910 9070 990 9090
rect 1150 9130 1230 9150
rect 1150 9090 1170 9130
rect 1210 9090 1230 9130
rect 1150 9070 1230 9090
rect 1390 9130 1470 9150
rect 1390 9090 1410 9130
rect 1450 9090 1470 9130
rect 1390 9070 1470 9090
rect 1630 9130 1710 9150
rect 1630 9090 1650 9130
rect 1690 9090 1710 9130
rect 1630 9070 1710 9090
rect 2270 9130 2350 9150
rect 2270 9090 2290 9130
rect 2330 9090 2350 9130
rect 2270 9070 2350 9090
rect 2510 9130 2590 9150
rect 2510 9090 2530 9130
rect 2570 9090 2590 9130
rect 2510 9070 2590 9090
rect 2750 9130 2830 9150
rect 2750 9090 2770 9130
rect 2810 9090 2830 9130
rect 2750 9070 2830 9090
rect 3710 9130 3790 9150
rect 3710 9090 3730 9130
rect 3770 9090 3790 9130
rect 3710 9070 3790 9090
rect 3950 9130 4030 9150
rect 3950 9090 3970 9130
rect 4010 9090 4030 9130
rect 3950 9070 4030 9090
rect 4190 9130 4270 9150
rect 4190 9090 4210 9130
rect 4250 9090 4270 9130
rect 4190 9070 4270 9090
rect 4830 9130 4910 9150
rect 4830 9090 4850 9130
rect 4890 9090 4910 9130
rect 4830 9070 4910 9090
rect 5070 9130 5150 9150
rect 5070 9090 5090 9130
rect 5130 9090 5150 9130
rect 5070 9070 5150 9090
rect 5310 9130 5390 9150
rect 5310 9090 5330 9130
rect 5370 9090 5390 9130
rect 5310 9070 5390 9090
rect 5550 9130 5630 9150
rect 5550 9090 5570 9130
rect 5610 9090 5630 9130
rect 5550 9070 5630 9090
rect 7840 8870 8270 8886
rect 7840 8836 7856 8870
rect 7890 8836 8270 8870
rect 7840 8820 8270 8836
rect 8750 8870 9180 8886
rect 8750 8836 9130 8870
rect 9164 8836 9180 8870
rect 8750 8820 9180 8836
rect 1421 8752 1479 8770
rect 1421 8718 1433 8752
rect 1467 8718 1479 8752
rect 1421 8700 1479 8718
rect 1781 8752 1839 8770
rect 1781 8718 1793 8752
rect 1827 8718 1839 8752
rect 1781 8700 1839 8718
rect 1901 8752 1959 8770
rect 1901 8718 1913 8752
rect 1947 8718 1959 8752
rect 1901 8700 1959 8718
rect 2261 8752 2319 8770
rect 2261 8718 2273 8752
rect 2307 8718 2319 8752
rect 2261 8700 2319 8718
rect 2381 8752 2439 8770
rect 2381 8718 2393 8752
rect 2427 8718 2439 8752
rect 2381 8700 2439 8718
rect 1430 8670 1470 8700
rect 1550 8670 1590 8700
rect 1670 8670 1710 8700
rect 1790 8670 1830 8700
rect 1910 8670 1950 8700
rect 2030 8670 2070 8700
rect 2150 8670 2190 8700
rect 2270 8670 2310 8700
rect 2390 8670 2430 8700
rect 2510 8670 2550 8700
rect 1430 8540 1470 8570
rect 1550 8540 1590 8570
rect 1522 8522 1590 8540
rect 1522 8488 1534 8522
rect 1568 8488 1590 8522
rect 1522 8470 1590 8488
rect 1670 8540 1710 8570
rect 1790 8540 1830 8570
rect 1910 8540 1950 8570
rect 2030 8540 2070 8570
rect 1670 8522 1738 8540
rect 1670 8488 1692 8522
rect 1726 8488 1738 8522
rect 1670 8470 1738 8488
rect 2004 8522 2070 8540
rect 2004 8488 2016 8522
rect 2050 8488 2070 8522
rect 2004 8470 2070 8488
rect 2150 8540 2190 8570
rect 2270 8540 2310 8570
rect 2390 8540 2430 8570
rect 2510 8540 2550 8570
rect 2150 8522 2216 8540
rect 2150 8488 2170 8522
rect 2204 8488 2216 8522
rect 2150 8470 2216 8488
rect 2482 8522 2550 8540
rect 2482 8488 2494 8522
rect 2528 8488 2550 8522
rect 4101 8752 4159 8770
rect 4101 8718 4113 8752
rect 4147 8718 4159 8752
rect 4101 8700 4159 8718
rect 4221 8752 4279 8770
rect 4221 8718 4233 8752
rect 4267 8718 4279 8752
rect 4221 8700 4279 8718
rect 4581 8752 4639 8770
rect 4581 8718 4593 8752
rect 4627 8718 4639 8752
rect 4581 8700 4639 8718
rect 4701 8752 4759 8770
rect 4701 8718 4713 8752
rect 4747 8718 4759 8752
rect 4701 8700 4759 8718
rect 5061 8752 5119 8770
rect 5061 8718 5073 8752
rect 5107 8718 5119 8752
rect 5061 8700 5119 8718
rect 9010 8700 9090 8720
rect 3990 8670 4030 8700
rect 4110 8670 4150 8700
rect 4230 8670 4270 8700
rect 4350 8670 4390 8700
rect 4470 8670 4510 8700
rect 4590 8670 4630 8700
rect 4710 8670 4750 8700
rect 4830 8670 4870 8700
rect 4950 8670 4990 8700
rect 5070 8670 5110 8700
rect 9010 8660 9030 8700
rect 9070 8660 9090 8700
rect 9410 8700 9490 8720
rect 9410 8660 9430 8700
rect 9470 8660 9490 8700
rect 8300 8610 8400 8640
rect 8500 8630 10000 8660
rect 8500 8610 8600 8630
rect 8700 8610 8800 8630
rect 8900 8610 9000 8630
rect 9100 8610 9200 8630
rect 9300 8610 9400 8630
rect 9500 8610 9600 8630
rect 9700 8610 9800 8630
rect 9900 8610 10000 8630
rect 10100 8610 10200 8640
rect 3990 8540 4030 8570
rect 4110 8540 4150 8570
rect 4230 8540 4270 8570
rect 4350 8540 4390 8570
rect 3990 8522 4058 8540
rect 2482 8470 2550 8488
rect 3990 8488 4012 8522
rect 4046 8488 4058 8522
rect 3990 8470 4058 8488
rect 4324 8522 4390 8540
rect 4324 8488 4336 8522
rect 4370 8488 4390 8522
rect 4324 8470 4390 8488
rect 4470 8540 4510 8570
rect 4590 8540 4630 8570
rect 4710 8540 4750 8570
rect 4830 8540 4870 8570
rect 4470 8522 4536 8540
rect 4470 8488 4490 8522
rect 4524 8488 4536 8522
rect 4470 8470 4536 8488
rect 4802 8522 4870 8540
rect 4802 8488 4814 8522
rect 4848 8488 4870 8522
rect 4802 8470 4870 8488
rect 4950 8540 4990 8570
rect 5070 8540 5110 8570
rect 4950 8522 5018 8540
rect 4950 8488 4972 8522
rect 5006 8488 5018 8522
rect 4950 8470 5018 8488
rect 8300 8330 8400 8360
rect 8500 8330 8600 8360
rect 8700 8330 8800 8360
rect 8900 8330 9000 8360
rect 9100 8330 9200 8360
rect 9300 8330 9400 8360
rect 9500 8330 9600 8360
rect 9700 8330 9800 8360
rect 9900 8330 10000 8360
rect 10100 8330 10200 8360
rect 8210 8310 8400 8330
rect 8210 8270 8230 8310
rect 8270 8300 8400 8310
rect 10100 8310 10290 8330
rect 10100 8300 10230 8310
rect 8270 8270 8290 8300
rect 8210 8250 8290 8270
rect 10210 8270 10230 8300
rect 10270 8270 10290 8310
rect 10210 8250 10290 8270
rect 8320 8020 8410 8040
rect 8320 7970 8340 8020
rect 8390 7970 8410 8020
rect 8320 7950 8410 7970
rect 8970 8020 9060 8040
rect 8970 7970 8990 8020
rect 9040 7970 9060 8020
rect 8970 7950 9060 7970
rect 9460 8010 9540 8030
rect 9460 7970 9480 8010
rect 9520 7970 9540 8010
rect 9460 7950 9540 7970
rect 10120 8010 10200 8030
rect 10120 7970 10140 8010
rect 10180 7970 10200 8010
rect 10120 7950 10200 7970
rect 10600 8010 10680 8030
rect 10600 7970 10620 8010
rect 10660 7970 10680 8010
rect 10600 7950 10680 7970
rect 11260 8010 11340 8030
rect 11260 7970 11280 8010
rect 11320 7970 11340 8010
rect 11260 7950 11340 7970
rect 700 7930 760 7950
rect 700 7890 710 7930
rect 750 7890 760 7930
rect 700 7870 760 7890
rect 870 7920 950 7940
rect 870 7880 890 7920
rect 930 7880 950 7920
rect 1360 7920 1420 7940
rect 1360 7880 1370 7920
rect 1410 7880 1420 7920
rect 1590 7920 1670 7940
rect 1590 7880 1610 7920
rect 1650 7880 1670 7920
rect 2080 7920 2140 7940
rect 2080 7880 2090 7920
rect 2130 7880 2140 7920
rect 2310 7920 2390 7940
rect 2310 7880 2330 7920
rect 2370 7880 2390 7920
rect 2740 7920 2800 7940
rect 2740 7880 2750 7920
rect 2790 7880 2800 7920
rect 590 7830 630 7860
rect 710 7830 750 7870
rect 830 7850 1230 7880
rect 830 7830 870 7850
rect 950 7830 990 7850
rect 1070 7830 1110 7850
rect 1190 7830 1230 7850
rect 1310 7850 1470 7880
rect 1310 7830 1350 7850
rect 1430 7830 1470 7850
rect 1550 7850 1950 7880
rect 1550 7830 1590 7850
rect 1670 7830 1710 7850
rect 1790 7830 1830 7850
rect 1910 7830 1950 7850
rect 2030 7850 2190 7880
rect 2030 7830 2070 7850
rect 2150 7830 2190 7850
rect 2270 7850 2670 7880
rect 2740 7860 2800 7880
rect 3740 7920 3800 7940
rect 3740 7880 3750 7920
rect 3790 7880 3800 7920
rect 4150 7920 4230 7940
rect 4150 7880 4170 7920
rect 4210 7880 4230 7920
rect 4400 7920 4460 7940
rect 4400 7880 4410 7920
rect 4450 7880 4460 7920
rect 4870 7920 4950 7940
rect 4870 7880 4890 7920
rect 4930 7880 4950 7920
rect 5120 7920 5180 7940
rect 5120 7880 5130 7920
rect 5170 7880 5180 7920
rect 5590 7920 5670 7940
rect 5590 7880 5610 7920
rect 5650 7880 5670 7920
rect 5780 7930 5840 7950
rect 5780 7890 5790 7930
rect 5830 7890 5840 7930
rect 8350 7920 8380 7950
rect 8480 7920 8510 7950
rect 8610 7920 8640 7950
rect 8740 7920 8770 7950
rect 8870 7920 8900 7950
rect 9000 7920 9030 7950
rect 9490 7920 9520 7950
rect 9620 7920 9650 7950
rect 9750 7920 9780 7950
rect 9880 7920 9910 7950
rect 10010 7920 10040 7950
rect 10140 7920 10170 7950
rect 10630 7920 10660 7950
rect 10760 7920 10790 7950
rect 10890 7920 10920 7950
rect 11020 7920 11050 7950
rect 11150 7920 11180 7950
rect 11280 7920 11310 7950
rect 3740 7860 3800 7880
rect 2270 7830 2310 7850
rect 2390 7830 2430 7850
rect 2510 7830 2550 7850
rect 2630 7830 2670 7850
rect 2750 7830 2790 7860
rect 2870 7830 2910 7860
rect 3630 7830 3670 7860
rect 3750 7830 3790 7860
rect 3870 7850 4270 7880
rect 3870 7830 3910 7850
rect 3990 7830 4030 7850
rect 4110 7830 4150 7850
rect 4230 7830 4270 7850
rect 4350 7850 4510 7880
rect 4350 7830 4390 7850
rect 4470 7830 4510 7850
rect 4590 7850 4990 7880
rect 4590 7830 4630 7850
rect 4710 7830 4750 7850
rect 4830 7830 4870 7850
rect 4950 7830 4990 7850
rect 5070 7850 5230 7880
rect 5070 7830 5110 7850
rect 5190 7830 5230 7850
rect 5310 7850 5710 7880
rect 5780 7870 5840 7890
rect 5310 7830 5350 7850
rect 5430 7830 5470 7850
rect 5550 7830 5590 7850
rect 5670 7830 5710 7850
rect 5790 7830 5830 7870
rect 5910 7830 5950 7860
rect 8350 7790 8380 7820
rect 8480 7800 8510 7820
rect 8610 7800 8640 7820
rect 8740 7800 8770 7820
rect 8870 7800 8900 7820
rect 8480 7770 8900 7800
rect 9000 7790 9030 7820
rect 9490 7790 9520 7820
rect 9620 7800 9650 7820
rect 9750 7800 9780 7820
rect 9620 7790 9780 7800
rect 9570 7770 9780 7790
rect 9880 7800 9910 7820
rect 10010 7800 10040 7820
rect 9880 7770 10040 7800
rect 10140 7790 10170 7820
rect 10630 7790 10660 7820
rect 8520 7730 8540 7770
rect 8580 7730 8600 7770
rect 8520 7710 8600 7730
rect 9570 7730 9590 7770
rect 9630 7730 9650 7770
rect 9570 7710 9650 7730
rect 10010 7750 10090 7770
rect 10010 7710 10030 7750
rect 10070 7710 10090 7750
rect 10010 7690 10090 7710
rect 10760 7740 10790 7820
rect 10890 7740 10920 7820
rect 11020 7740 11050 7820
rect 11150 7740 11180 7820
rect 11280 7790 11310 7820
rect 11550 7770 11630 7790
rect 11550 7740 11570 7770
rect 10760 7730 11570 7740
rect 11610 7730 11630 7770
rect 10760 7710 11630 7730
rect 10760 7670 10790 7710
rect 10710 7650 10790 7670
rect 590 7600 630 7630
rect 710 7600 750 7630
rect 830 7600 870 7630
rect 950 7600 990 7630
rect 1070 7600 1110 7630
rect 1190 7600 1230 7630
rect 1310 7600 1350 7630
rect 1430 7600 1470 7630
rect 1550 7600 1590 7630
rect 1670 7600 1710 7630
rect 1790 7600 1830 7630
rect 1910 7600 1950 7630
rect 2030 7600 2070 7630
rect 2150 7600 2190 7630
rect 2270 7600 2310 7630
rect 2390 7600 2430 7630
rect 2510 7600 2550 7630
rect 2630 7600 2670 7630
rect 2750 7600 2790 7630
rect 2870 7600 2910 7630
rect 3630 7600 3670 7630
rect 3750 7600 3790 7630
rect 3870 7600 3910 7630
rect 3990 7600 4030 7630
rect 4110 7600 4150 7630
rect 4230 7600 4270 7630
rect 4350 7600 4390 7630
rect 4470 7600 4510 7630
rect 4590 7600 4630 7630
rect 4710 7600 4750 7630
rect 4830 7600 4870 7630
rect 4950 7600 4990 7630
rect 5070 7600 5110 7630
rect 5190 7600 5230 7630
rect 5310 7600 5350 7630
rect 5430 7600 5470 7630
rect 5550 7600 5590 7630
rect 5670 7600 5710 7630
rect 5790 7600 5830 7630
rect 5910 7600 5950 7630
rect 10710 7610 10730 7650
rect 10770 7610 10790 7650
rect 520 7580 630 7600
rect 520 7540 530 7580
rect 570 7570 630 7580
rect 2870 7580 2980 7600
rect 2870 7570 2930 7580
rect 570 7540 580 7570
rect 520 7520 580 7540
rect 2920 7540 2930 7570
rect 2970 7540 2980 7580
rect 2920 7520 2980 7540
rect 3560 7580 3670 7600
rect 3560 7540 3570 7580
rect 3610 7570 3670 7580
rect 5910 7580 6020 7600
rect 10710 7590 10790 7610
rect 5910 7570 5970 7580
rect 3610 7540 3620 7570
rect 3560 7520 3620 7540
rect 5960 7540 5970 7570
rect 6010 7540 6020 7580
rect 5960 7520 6020 7540
rect 8430 7440 8510 7460
rect 8430 7400 8450 7440
rect 8490 7400 8510 7440
rect 8870 7440 8950 7460
rect 8870 7400 8890 7440
rect 8930 7400 8950 7440
rect 9660 7450 9740 7470
rect 9660 7410 9680 7450
rect 9720 7410 9740 7450
rect 10710 7440 11630 7460
rect 9660 7400 9740 7410
rect 9960 7400 10040 7420
rect 8430 7380 8640 7400
rect 8350 7350 8380 7380
rect 8480 7370 8640 7380
rect 8480 7350 8510 7370
rect 8610 7350 8640 7370
rect 8740 7380 8950 7400
rect 8740 7370 8900 7380
rect 8740 7350 8770 7370
rect 8870 7350 8900 7370
rect 9000 7350 9030 7380
rect 9490 7350 9520 7380
rect 9620 7370 10040 7400
rect 10710 7400 10730 7440
rect 10770 7430 11570 7440
rect 10770 7400 10790 7430
rect 10710 7380 10790 7400
rect 9620 7350 9650 7370
rect 9750 7350 9780 7370
rect 9880 7350 9910 7370
rect 10010 7350 10040 7370
rect 10140 7350 10170 7380
rect 10630 7350 10660 7380
rect 10760 7350 10790 7380
rect 10890 7350 10920 7430
rect 11020 7350 11050 7430
rect 11150 7350 11180 7430
rect 11550 7400 11570 7430
rect 11610 7400 11630 7440
rect 11550 7380 11630 7400
rect 11280 7350 11310 7380
rect 8350 7120 8380 7150
rect 8480 7120 8510 7150
rect 8610 7120 8640 7150
rect 8740 7120 8770 7150
rect 8870 7120 8900 7150
rect 9000 7120 9030 7150
rect 9490 7120 9520 7150
rect 9620 7120 9650 7150
rect 9750 7120 9780 7150
rect 9880 7120 9910 7150
rect 10010 7120 10040 7150
rect 10140 7120 10170 7150
rect 10630 7120 10660 7150
rect 10760 7120 10790 7150
rect 10890 7120 10920 7150
rect 11020 7120 11050 7150
rect 11150 7120 11180 7150
rect 11280 7120 11310 7150
rect 8320 7100 8400 7120
rect 8320 7060 8340 7100
rect 8380 7060 8400 7100
rect 8320 7040 8400 7060
rect 8980 7100 9060 7120
rect 8980 7060 9000 7100
rect 9040 7060 9060 7100
rect 8980 7040 9060 7060
rect 9460 7100 9540 7120
rect 9460 7060 9480 7100
rect 9520 7060 9540 7100
rect 9460 7040 9540 7060
rect 10120 7100 10200 7120
rect 10120 7060 10140 7100
rect 10180 7060 10200 7100
rect 10120 7040 10200 7060
rect 10600 7100 10680 7120
rect 10600 7060 10620 7100
rect 10660 7060 10680 7100
rect 10600 7040 10680 7060
rect 11260 7100 11340 7120
rect 11260 7060 11280 7100
rect 11320 7060 11340 7100
rect 11260 7040 11340 7060
rect 8330 6790 8410 6810
rect 1890 6760 1960 6780
rect 1890 6720 1900 6760
rect 1940 6720 1960 6760
rect 1890 6700 1960 6720
rect 2060 6760 2140 6780
rect 2060 6720 2080 6760
rect 2120 6720 2140 6760
rect 2060 6700 2140 6720
rect 2240 6760 2320 6780
rect 2240 6720 2260 6760
rect 2300 6720 2320 6760
rect 2240 6700 2320 6720
rect 2420 6760 2500 6780
rect 2420 6720 2440 6760
rect 2480 6720 2500 6760
rect 2420 6700 2500 6720
rect 2600 6760 2680 6780
rect 2600 6720 2620 6760
rect 2660 6720 2680 6760
rect 2600 6700 2680 6720
rect 2780 6760 2860 6780
rect 2780 6720 2800 6760
rect 2840 6720 2860 6760
rect 2780 6700 2860 6720
rect 2960 6760 3040 6780
rect 2960 6720 2980 6760
rect 3020 6720 3040 6760
rect 2960 6700 3040 6720
rect 3140 6760 3210 6780
rect 3140 6720 3160 6760
rect 3200 6720 3210 6760
rect 3140 6700 3210 6720
rect 3330 6760 3400 6780
rect 3330 6720 3340 6760
rect 3380 6720 3400 6760
rect 3330 6700 3400 6720
rect 3500 6760 3580 6780
rect 3500 6720 3520 6760
rect 3560 6720 3580 6760
rect 3500 6700 3580 6720
rect 3680 6760 3760 6780
rect 3680 6720 3700 6760
rect 3740 6720 3760 6760
rect 3680 6700 3760 6720
rect 3860 6760 3940 6780
rect 3860 6720 3880 6760
rect 3920 6720 3940 6760
rect 3860 6700 3940 6720
rect 4040 6760 4120 6780
rect 4040 6720 4060 6760
rect 4100 6720 4120 6760
rect 4040 6700 4120 6720
rect 4220 6760 4300 6780
rect 4220 6720 4240 6760
rect 4280 6720 4300 6760
rect 4220 6700 4300 6720
rect 4400 6760 4480 6780
rect 4400 6720 4420 6760
rect 4460 6720 4480 6760
rect 4400 6700 4480 6720
rect 4580 6760 4650 6780
rect 4580 6720 4600 6760
rect 4640 6720 4650 6760
rect 8330 6750 8350 6790
rect 8390 6760 8410 6790
rect 10330 6790 10410 6810
rect 10330 6760 10350 6790
rect 8390 6750 8520 6760
rect 8330 6730 8520 6750
rect 10220 6750 10350 6760
rect 10390 6750 10410 6790
rect 10220 6730 10410 6750
rect 4580 6710 4650 6720
rect 1690 6670 1790 6700
rect 1870 6670 1970 6700
rect 2050 6670 2150 6700
rect 2230 6670 2330 6700
rect 2410 6670 2510 6700
rect 2590 6670 2690 6700
rect 2770 6670 2870 6700
rect 2950 6670 3050 6700
rect 3130 6670 3230 6700
rect 3310 6670 3410 6700
rect 3490 6670 3590 6700
rect 3670 6670 3770 6700
rect 3850 6670 3950 6700
rect 4030 6670 4130 6700
rect 4210 6670 4310 6700
rect 4390 6670 4490 6700
rect 4570 6670 4670 6710
rect 8420 6700 8520 6730
rect 8620 6700 8720 6730
rect 8820 6700 8920 6730
rect 9020 6700 9120 6730
rect 9220 6700 9320 6730
rect 9420 6700 9520 6730
rect 9620 6700 9720 6730
rect 9820 6700 9920 6730
rect 10020 6700 10120 6730
rect 10220 6700 10320 6730
rect 4750 6670 4850 6700
rect 5700 6560 5780 6580
rect 5700 6520 5720 6560
rect 5760 6520 5780 6560
rect 5560 6470 5590 6500
rect 5670 6490 5810 6520
rect 5670 6470 5700 6490
rect 5780 6470 5810 6490
rect 5890 6470 5920 6500
rect 5560 6250 5590 6270
rect 5490 6220 5590 6250
rect 5670 6240 5700 6270
rect 5780 6240 5810 6270
rect 5890 6250 5920 6270
rect 5890 6220 5990 6250
rect 5490 6180 5500 6220
rect 5540 6180 5550 6220
rect 5490 6160 5550 6180
rect 5930 6180 5940 6220
rect 5980 6180 5990 6220
rect 5930 6160 5990 6180
rect 8420 6170 8520 6200
rect 8620 6180 8720 6200
rect 8820 6180 8920 6200
rect 9020 6180 9120 6200
rect 9220 6180 9320 6200
rect 9420 6180 9520 6200
rect 9620 6180 9720 6200
rect 9820 6180 9920 6200
rect 10020 6180 10120 6200
rect 8620 6150 10120 6180
rect 10220 6170 10320 6200
rect 9130 6110 9150 6150
rect 9190 6110 9210 6150
rect 9130 6090 9210 6110
rect 9530 6110 9550 6150
rect 9590 6110 9610 6150
rect 9530 6090 9610 6110
rect 1690 6040 1790 6070
rect 1870 6040 1970 6070
rect 2050 6040 2150 6070
rect 2230 6040 2330 6070
rect 2410 6040 2510 6070
rect 2590 6040 2690 6070
rect 2770 6040 2870 6070
rect 2950 6040 3050 6070
rect 3130 6040 3230 6070
rect 3310 6040 3410 6070
rect 3490 6040 3590 6070
rect 3670 6040 3770 6070
rect 3850 6040 3950 6070
rect 4030 6040 4130 6070
rect 4210 6040 4310 6070
rect 4390 6040 4490 6070
rect 4570 6040 4670 6070
rect 4750 6040 4850 6070
rect 1610 6020 1790 6040
rect 1610 5980 1630 6020
rect 1670 6010 1790 6020
rect 4750 6020 4930 6040
rect 4750 6010 4870 6020
rect 1670 5980 1690 6010
rect 1610 5960 1690 5980
rect 4850 5980 4870 6010
rect 4910 5980 4930 6020
rect 4850 5960 4930 5980
rect 1796 5752 1854 5770
rect 1796 5718 1808 5752
rect 1842 5718 1854 5752
rect 1796 5700 1854 5718
rect 1906 5752 1964 5770
rect 1906 5718 1918 5752
rect 1952 5718 1964 5752
rect 1906 5700 1964 5718
rect 2016 5752 2074 5770
rect 2016 5718 2028 5752
rect 2062 5718 2074 5752
rect 2016 5700 2074 5718
rect 2126 5752 2184 5770
rect 2126 5718 2138 5752
rect 2172 5718 2184 5752
rect 2126 5700 2184 5718
rect 2236 5752 2294 5770
rect 2236 5718 2248 5752
rect 2282 5718 2294 5752
rect 2236 5700 2294 5718
rect 2346 5752 2404 5770
rect 2346 5718 2358 5752
rect 2392 5718 2404 5752
rect 2346 5700 2404 5718
rect 2456 5752 2514 5770
rect 2456 5718 2468 5752
rect 2502 5718 2514 5752
rect 2456 5700 2514 5718
rect 2566 5752 2624 5770
rect 2566 5718 2578 5752
rect 2612 5718 2624 5752
rect 2566 5700 2624 5718
rect 2676 5752 2734 5770
rect 2676 5718 2688 5752
rect 2722 5718 2734 5752
rect 2676 5700 2734 5718
rect 2786 5752 2844 5770
rect 2786 5718 2798 5752
rect 2832 5718 2844 5752
rect 2786 5700 2844 5718
rect 3696 5752 3754 5770
rect 3696 5718 3708 5752
rect 3742 5718 3754 5752
rect 3696 5700 3754 5718
rect 3806 5752 3864 5770
rect 3806 5718 3818 5752
rect 3852 5718 3864 5752
rect 3806 5700 3864 5718
rect 3916 5752 3974 5770
rect 3916 5718 3928 5752
rect 3962 5718 3974 5752
rect 3916 5700 3974 5718
rect 4026 5752 4084 5770
rect 4026 5718 4038 5752
rect 4072 5718 4084 5752
rect 4026 5700 4084 5718
rect 4136 5752 4194 5770
rect 4136 5718 4148 5752
rect 4182 5718 4194 5752
rect 4136 5700 4194 5718
rect 4246 5752 4304 5770
rect 4246 5718 4258 5752
rect 4292 5718 4304 5752
rect 4246 5700 4304 5718
rect 4356 5752 4414 5770
rect 4356 5718 4368 5752
rect 4402 5718 4414 5752
rect 4356 5700 4414 5718
rect 4466 5752 4524 5770
rect 4466 5718 4478 5752
rect 4512 5718 4524 5752
rect 4466 5700 4524 5718
rect 4576 5752 4634 5770
rect 4576 5718 4588 5752
rect 4622 5718 4634 5752
rect 4576 5700 4634 5718
rect 4686 5752 4744 5770
rect 4686 5718 4698 5752
rect 4732 5718 4744 5752
rect 4686 5700 4744 5718
rect 1700 5670 1730 5700
rect 1810 5670 1840 5700
rect 1920 5670 1950 5700
rect 2030 5670 2060 5700
rect 2140 5670 2170 5700
rect 2250 5670 2280 5700
rect 2360 5670 2390 5700
rect 2470 5670 2500 5700
rect 2580 5670 2610 5700
rect 2690 5670 2720 5700
rect 2800 5670 2830 5700
rect 2910 5670 2940 5700
rect 3600 5670 3630 5700
rect 3710 5670 3740 5700
rect 3820 5670 3850 5700
rect 3930 5670 3960 5700
rect 4040 5670 4070 5700
rect 4150 5670 4180 5700
rect 4260 5670 4290 5700
rect 4370 5670 4400 5700
rect 4480 5670 4510 5700
rect 4590 5670 4620 5700
rect 4700 5670 4730 5700
rect 4810 5670 4840 5700
rect 1700 5440 1730 5470
rect 1810 5440 1840 5470
rect 1920 5440 1950 5470
rect 2030 5440 2060 5470
rect 2140 5440 2170 5470
rect 2250 5440 2280 5470
rect 2360 5440 2390 5470
rect 2470 5440 2500 5470
rect 2580 5440 2610 5470
rect 2690 5440 2720 5470
rect 2800 5440 2830 5470
rect 2910 5440 2940 5470
rect 3600 5440 3630 5470
rect 3710 5440 3740 5470
rect 3820 5440 3850 5470
rect 3930 5440 3960 5470
rect 4040 5440 4070 5470
rect 4150 5440 4180 5470
rect 4260 5440 4290 5470
rect 4370 5440 4400 5470
rect 4480 5440 4510 5470
rect 4590 5440 4620 5470
rect 4700 5440 4730 5470
rect 4810 5440 4840 5470
rect 1620 5420 1730 5440
rect 1620 5380 1640 5420
rect 1680 5410 1730 5420
rect 2910 5420 3020 5440
rect 2910 5410 2960 5420
rect 1680 5380 1700 5410
rect 1620 5360 1700 5380
rect 2940 5380 2960 5410
rect 3000 5380 3020 5420
rect 2940 5360 3020 5380
rect 3520 5420 3630 5440
rect 3520 5380 3540 5420
rect 3580 5410 3630 5420
rect 4810 5420 4920 5440
rect 4810 5410 4860 5420
rect 3580 5380 3600 5410
rect 3520 5360 3600 5380
rect 4840 5380 4860 5410
rect 4900 5380 4920 5420
rect 4840 5360 4920 5380
rect 2740 4810 3150 4840
rect 2220 4730 2250 4760
rect 2330 4730 2360 4760
rect 2740 4730 2770 4810
rect 2850 4730 2880 4760
rect 3120 4730 3150 4810
rect 4270 4820 4350 4840
rect 4270 4780 4290 4820
rect 4330 4780 4350 4820
rect 4270 4760 4350 4780
rect 3230 4730 3260 4760
rect 3640 4730 3670 4760
rect 3750 4730 3780 4760
rect 4160 4730 4190 4760
rect 4270 4730 4300 4760
rect 4600 4730 4630 4760
rect 4930 4730 4960 4760
rect 5370 4730 5400 4760
rect 5760 4730 5790 4760
rect 6150 4730 6180 4760
rect 6440 4730 6470 4760
rect 1930 4470 2010 4490
rect 1930 4430 1950 4470
rect 1990 4460 2010 4470
rect 2220 4460 2250 4530
rect 1990 4430 2250 4460
rect 1930 4410 2010 4430
rect 2220 4310 2250 4430
rect 2330 4500 2360 4530
rect 2330 4480 2430 4500
rect 2740 4490 2770 4530
rect 2330 4440 2370 4480
rect 2410 4440 2430 4480
rect 2330 4420 2430 4440
rect 2520 4460 2770 4490
rect 2330 4310 2360 4420
rect 2520 4000 2550 4460
rect 2740 4310 2770 4460
rect 2850 4420 2880 4530
rect 2850 4400 2950 4420
rect 2850 4360 2890 4400
rect 2930 4360 2950 4400
rect 2850 4340 2950 4360
rect 2850 4310 2880 4340
rect 3120 4310 3150 4530
rect 3230 4500 3260 4530
rect 3230 4480 3330 4500
rect 3640 4490 3670 4530
rect 3230 4440 3270 4480
rect 3310 4440 3330 4480
rect 3230 4420 3330 4440
rect 3420 4460 3670 4490
rect 3230 4310 3260 4420
rect 2470 3980 2550 4000
rect 2470 3940 2490 3980
rect 2530 3940 2550 3980
rect 2470 3920 2550 3940
rect 3420 4000 3450 4460
rect 3640 4310 3670 4460
rect 3750 4490 3780 4530
rect 3750 4470 3920 4490
rect 3750 4460 3860 4470
rect 3750 4310 3780 4460
rect 3840 4430 3860 4460
rect 3900 4430 3920 4470
rect 3840 4410 3920 4430
rect 4160 4310 4190 4530
rect 4270 4310 4300 4530
rect 4350 4430 4430 4450
rect 4600 4430 4630 4530
rect 4350 4390 4370 4430
rect 4410 4400 4630 4430
rect 4410 4390 4430 4400
rect 4350 4370 4430 4390
rect 4600 4310 4630 4400
rect 4680 4430 4760 4450
rect 4930 4430 4960 4530
rect 5140 4460 5220 4480
rect 4680 4390 4700 4430
rect 4740 4400 4960 4430
rect 4740 4390 4760 4400
rect 4680 4370 4760 4390
rect 4930 4310 4960 4400
rect 5010 4430 5090 4450
rect 5010 4390 5030 4430
rect 5070 4390 5090 4430
rect 5140 4420 5160 4460
rect 5200 4430 5220 4460
rect 5370 4430 5400 4530
rect 5760 4450 5790 4530
rect 6150 4500 6180 4530
rect 6440 4500 6470 4530
rect 5200 4420 5400 4430
rect 5140 4400 5400 4420
rect 5010 4370 5090 4390
rect 5370 4310 5400 4400
rect 5710 4430 5790 4450
rect 5710 4390 5730 4430
rect 5770 4390 5790 4430
rect 6100 4480 6860 4500
rect 6100 4440 6120 4480
rect 6160 4470 6860 4480
rect 6160 4440 6180 4470
rect 6100 4420 6180 4440
rect 5710 4370 5790 4390
rect 5760 4310 5790 4370
rect 6150 4310 6180 4420
rect 6230 4400 6310 4420
rect 6230 4360 6250 4400
rect 6290 4370 6310 4400
rect 6640 4400 6720 4420
rect 6640 4370 6660 4400
rect 6290 4360 6660 4370
rect 6700 4360 6720 4400
rect 6230 4340 6720 4360
rect 6440 4310 6470 4340
rect 6830 4310 6860 4470
rect 8150 4450 8230 4470
rect 8150 4410 8170 4450
rect 8210 4420 8230 4450
rect 10990 4450 11070 4470
rect 10990 4420 11010 4450
rect 8210 4410 8360 4420
rect 8150 4390 8360 4410
rect 8240 4360 8360 4390
rect 8460 4380 9240 4420
rect 8460 4360 8580 4380
rect 8680 4360 8800 4380
rect 8900 4360 9020 4380
rect 9120 4360 9240 4380
rect 9340 4360 9460 4390
rect 9760 4360 9880 4390
rect 9980 4380 10760 4420
rect 9980 4360 10100 4380
rect 10200 4360 10320 4380
rect 10420 4360 10540 4380
rect 10640 4360 10760 4380
rect 10860 4410 11010 4420
rect 11050 4410 11070 4450
rect 10860 4390 11070 4410
rect 10860 4360 10980 4390
rect 3370 3980 3450 4000
rect 3370 3940 3390 3980
rect 3430 3940 3450 3980
rect 3370 3920 3450 3940
rect 8240 3930 8360 3960
rect 8460 3940 8580 3960
rect 8680 3940 8800 3960
rect 8900 3940 9020 3960
rect 9120 3940 9240 3960
rect 2220 3880 2250 3910
rect 2330 3880 2360 3910
rect 2740 3880 2770 3910
rect 2850 3880 2880 3910
rect 3120 3880 3150 3910
rect 3230 3880 3260 3910
rect 3640 3880 3670 3910
rect 3750 3880 3780 3910
rect 4160 3880 4190 3910
rect 4270 3880 4300 3910
rect 4600 3880 4630 3910
rect 4930 3880 4960 3910
rect 5370 3880 5400 3910
rect 5760 3880 5790 3910
rect 6150 3880 6180 3910
rect 6440 3880 6470 3910
rect 6830 3880 6860 3910
rect 8460 3900 9240 3940
rect 9340 3940 9460 3960
rect 9760 3940 9880 3960
rect 9340 3910 9880 3940
rect 9980 3930 10100 3960
rect 10200 3930 10320 3960
rect 10420 3930 10540 3960
rect 10640 3930 10760 3960
rect 10860 3930 10980 3960
rect 8460 3880 8540 3900
rect 4140 3860 4220 3880
rect 4140 3820 4160 3860
rect 4200 3820 4220 3860
rect 8460 3840 8480 3880
rect 8520 3840 8540 3880
rect 9570 3870 9590 3910
rect 9630 3870 9650 3910
rect 9570 3850 9650 3870
rect 9980 3900 10760 3930
rect 9980 3880 10060 3900
rect 8460 3820 8540 3840
rect 9980 3840 10000 3880
rect 10040 3840 10060 3880
rect 9980 3820 10060 3840
rect 10680 3880 10760 3900
rect 10680 3840 10700 3880
rect 10740 3840 10760 3880
rect 10680 3820 10760 3840
rect 4140 3800 4220 3820
rect 2590 3640 2670 3660
rect 2590 3600 2610 3640
rect 2650 3600 2670 3640
rect 2590 3580 2670 3600
rect 5710 3640 5790 3660
rect 5710 3600 5730 3640
rect 5770 3600 5790 3640
rect 5710 3580 5790 3600
rect 8390 3600 8470 3620
rect 2220 3550 2250 3580
rect 2330 3550 2360 3580
rect 2740 3550 2770 3580
rect 2850 3550 2880 3580
rect 3120 3550 3150 3580
rect 3230 3550 3260 3580
rect 3640 3550 3670 3580
rect 3750 3550 3780 3580
rect 4150 3550 4180 3580
rect 4480 3550 4510 3580
rect 4810 3550 4840 3580
rect 5370 3550 5400 3580
rect 5760 3550 5790 3580
rect 6150 3550 6180 3580
rect 6440 3550 6470 3580
rect 8390 3560 8410 3600
rect 8450 3560 8470 3600
rect 2470 3520 2550 3540
rect 2470 3480 2490 3520
rect 2530 3480 2550 3520
rect 2470 3460 2550 3480
rect 2020 3030 2100 3050
rect 2220 3030 2250 3150
rect 2020 2990 2040 3030
rect 2080 3000 2250 3030
rect 2080 2990 2100 3000
rect 2020 2970 2100 2990
rect 2220 2930 2250 3000
rect 2330 3040 2360 3150
rect 2330 3020 2430 3040
rect 2330 2980 2370 3020
rect 2410 2980 2430 3020
rect 2330 2960 2430 2980
rect 2520 3000 2550 3460
rect 3370 3520 3450 3540
rect 3370 3480 3390 3520
rect 3430 3480 3450 3520
rect 3370 3460 3450 3480
rect 2740 3000 2770 3150
rect 2520 2970 2770 3000
rect 2330 2930 2360 2960
rect 2740 2930 2770 2970
rect 2850 3120 2880 3150
rect 2850 3100 2950 3120
rect 2850 3060 2890 3100
rect 2930 3060 2950 3100
rect 2850 3040 2950 3060
rect 2850 2930 2880 3040
rect 3120 2930 3150 3150
rect 3230 3040 3260 3150
rect 3230 3020 3330 3040
rect 3230 2980 3270 3020
rect 3310 2980 3330 3020
rect 3230 2960 3330 2980
rect 3420 3000 3450 3460
rect 8390 3440 8470 3560
rect 10420 3500 10500 3520
rect 8930 3470 9010 3490
rect 8040 3380 8160 3410
rect 8260 3400 8600 3440
rect 8930 3430 8950 3470
rect 8990 3430 9010 3470
rect 10010 3470 10090 3490
rect 10010 3430 10030 3470
rect 10070 3430 10090 3470
rect 10420 3460 10440 3500
rect 10480 3460 10500 3500
rect 10420 3440 10500 3460
rect 10680 3500 10760 3520
rect 10680 3460 10700 3500
rect 10740 3460 10760 3500
rect 10680 3440 10760 3460
rect 8260 3380 8380 3400
rect 8480 3380 8600 3400
rect 8700 3400 9240 3430
rect 8700 3380 8820 3400
rect 9120 3380 9240 3400
rect 9340 3400 9680 3430
rect 9340 3380 9460 3400
rect 9560 3380 9680 3400
rect 9780 3400 10320 3430
rect 9780 3380 9900 3400
rect 10200 3380 10320 3400
rect 10420 3410 10760 3440
rect 10420 3380 10540 3410
rect 10640 3380 10760 3410
rect 10860 3380 10980 3410
rect 3640 3000 3670 3150
rect 3420 2970 3670 3000
rect 3230 2930 3260 2960
rect 3640 2930 3670 2970
rect 3750 3090 3780 3150
rect 3750 3070 4100 3090
rect 3750 3060 3880 3070
rect 3750 2930 3780 3060
rect 3860 3030 3880 3060
rect 3920 3060 4040 3070
rect 3920 3030 3940 3060
rect 3860 3010 3940 3030
rect 4020 3030 4040 3060
rect 4080 3030 4100 3070
rect 4020 3010 4100 3030
rect 4150 3060 4180 3150
rect 4350 3070 4430 3090
rect 4350 3060 4370 3070
rect 4150 3030 4370 3060
rect 4410 3030 4430 3070
rect 4150 2930 4180 3030
rect 4350 3010 4430 3030
rect 4480 3060 4510 3150
rect 4680 3070 4760 3090
rect 4680 3060 4700 3070
rect 4480 3030 4700 3060
rect 4740 3030 4760 3070
rect 4480 2930 4510 3030
rect 4680 3010 4760 3030
rect 4810 3060 4840 3150
rect 4940 3070 5020 3090
rect 4940 3060 4960 3070
rect 4810 3030 4960 3060
rect 5000 3030 5020 3070
rect 4810 2930 4840 3030
rect 4940 3010 5020 3030
rect 5140 3060 5220 3080
rect 5140 3020 5160 3060
rect 5200 3030 5220 3060
rect 5370 3030 5400 3150
rect 5760 3120 5790 3150
rect 6150 3110 6180 3150
rect 6440 3110 6470 3150
rect 5840 3090 6860 3110
rect 5840 3050 5860 3090
rect 5900 3080 6860 3090
rect 5900 3050 5920 3080
rect 5840 3030 5920 3050
rect 5200 3020 5400 3030
rect 5140 3000 5400 3020
rect 5370 2930 5400 3000
rect 5760 2930 5790 2960
rect 6150 2930 6180 3080
rect 6230 3010 6310 3020
rect 6230 2970 6250 3010
rect 6290 2980 6310 3010
rect 6290 2970 6470 2980
rect 6230 2950 6470 2970
rect 6440 2930 6470 2950
rect 6830 2930 6860 3080
rect 8040 2950 8160 2980
rect 7950 2930 8160 2950
rect 7950 2890 7970 2930
rect 8010 2920 8160 2930
rect 8260 2960 8380 2980
rect 8480 2960 8600 2980
rect 8260 2920 8600 2960
rect 8700 2950 8820 2980
rect 9120 2950 9240 2980
rect 9340 2960 9460 2980
rect 9560 2960 9680 2980
rect 8010 2890 8030 2920
rect 7950 2870 8030 2890
rect 8480 2900 8600 2920
rect 9340 2920 9680 2960
rect 9780 2950 9900 2980
rect 10200 2950 10320 2980
rect 10420 2960 10540 2980
rect 10640 2960 10760 2980
rect 10420 2920 10760 2960
rect 10860 2950 10980 2980
rect 10860 2930 11070 2950
rect 10860 2920 11010 2930
rect 9340 2900 9460 2920
rect 8480 2870 9460 2900
rect 10990 2890 11010 2920
rect 11050 2890 11070 2930
rect 10990 2870 11070 2890
rect 2220 2700 2250 2730
rect 2330 2700 2360 2730
rect 2740 2650 2770 2730
rect 2850 2700 2880 2730
rect 3120 2650 3150 2730
rect 3230 2700 3260 2730
rect 3640 2700 3670 2730
rect 3750 2700 3780 2730
rect 4150 2700 4180 2730
rect 4480 2700 4510 2730
rect 4810 2700 4840 2730
rect 5370 2700 5400 2730
rect 5760 2700 5790 2730
rect 6150 2700 6180 2730
rect 6440 2700 6470 2730
rect 6830 2700 6860 2730
rect 2740 2620 3150 2650
rect 5760 2680 5870 2700
rect 5760 2640 5810 2680
rect 5850 2640 5870 2680
rect 5760 2620 5870 2640
rect 6430 2680 6510 2700
rect 6430 2640 6450 2680
rect 6490 2640 6510 2680
rect 6430 2620 6510 2640
rect 12480 2000 12510 2030
rect 13080 2000 13110 2030
rect 13680 2000 13710 2030
rect 13950 2000 13980 2030
rect 14300 1810 14380 1830
rect 12480 1780 12510 1800
rect 13080 1780 13110 1800
rect 13680 1780 13710 1800
rect 13950 1780 13980 1800
rect 14300 1780 14320 1810
rect 12480 1770 14320 1780
rect 14360 1770 14380 1810
rect 12480 1750 14380 1770
rect 12480 1670 12510 1700
rect 13080 1670 13110 1700
rect 13680 1670 13710 1700
rect 1780 1530 1860 1550
rect 1780 1490 1800 1530
rect 1840 1490 1860 1530
rect 1780 1470 1860 1490
rect 2730 1510 2810 1530
rect 2730 1470 2750 1510
rect 2790 1470 2810 1510
rect 3800 1520 3880 1540
rect 3800 1480 3820 1520
rect 3860 1480 3880 1520
rect 3800 1470 3880 1480
rect 5360 1520 5450 1540
rect 5360 1480 5380 1520
rect 5420 1480 5450 1520
rect 5360 1470 5450 1480
rect 7974 1530 8040 1550
rect 8540 1530 8570 1560
rect 8650 1530 8680 1560
rect 8760 1530 8790 1560
rect 8870 1530 8900 1560
rect 9200 1530 9230 1560
rect 9310 1530 9340 1560
rect 9420 1530 9450 1560
rect 9840 1530 9870 1560
rect 9950 1530 9980 1560
rect 10060 1530 10090 1560
rect 10170 1530 10200 1560
rect 10500 1530 10530 1560
rect 10610 1530 10640 1560
rect 10720 1530 10750 1560
rect 11140 1530 11170 1560
rect 11250 1530 11280 1560
rect 11360 1530 11390 1560
rect 11470 1530 11500 1560
rect 11800 1530 11830 1560
rect 11910 1530 11940 1560
rect 12020 1530 12050 1560
rect 12480 1540 12510 1570
rect 13080 1540 13110 1570
rect 13680 1540 13710 1570
rect 7974 1490 7984 1530
rect 8024 1490 8040 1530
rect 7974 1470 8040 1490
rect 1910 1440 1940 1470
rect 2020 1440 2050 1470
rect 2130 1440 2160 1470
rect 2240 1440 2270 1470
rect 2490 1440 2520 1470
rect 2600 1440 2630 1470
rect 2730 1450 2810 1470
rect 1910 1310 1940 1340
rect 2020 1320 2050 1340
rect 2130 1320 2160 1340
rect 2240 1320 2270 1340
rect 2490 1320 2520 1340
rect 2020 1310 2520 1320
rect 1890 1290 1970 1310
rect 2020 1290 2550 1310
rect 1890 1250 1910 1290
rect 1950 1250 1970 1290
rect 1890 1230 1970 1250
rect 2070 1120 2100 1290
rect 2470 1250 2490 1290
rect 2530 1250 2550 1290
rect 2470 1230 2550 1250
rect 2600 1210 2630 1340
rect 2730 1210 2760 1450
rect 2940 1440 2970 1470
rect 3050 1440 3080 1470
rect 3160 1440 3190 1470
rect 3270 1440 3300 1470
rect 3600 1440 3630 1470
rect 3710 1440 3740 1470
rect 3820 1440 3850 1470
rect 3930 1440 3960 1470
rect 4280 1440 4310 1470
rect 4390 1440 4420 1470
rect 4500 1440 4530 1470
rect 4610 1440 4640 1470
rect 4860 1440 4890 1470
rect 4970 1440 5000 1470
rect 5420 1440 5450 1470
rect 5780 1440 5810 1470
rect 6030 1440 6060 1470
rect 6140 1440 6170 1470
rect 6250 1440 6280 1470
rect 6360 1440 6390 1470
rect 6690 1440 6720 1470
rect 6800 1440 6830 1470
rect 6910 1440 6940 1470
rect 7240 1440 7270 1470
rect 7350 1440 7380 1470
rect 7460 1440 7490 1470
rect 7570 1440 7600 1470
rect 7900 1440 7930 1470
rect 8010 1440 8040 1470
rect 8120 1440 8150 1470
rect 12480 1520 12710 1540
rect 12480 1510 12650 1520
rect 12630 1480 12650 1510
rect 12690 1480 12710 1520
rect 13080 1520 13310 1540
rect 13080 1510 13250 1520
rect 12630 1460 12710 1480
rect 13230 1480 13250 1510
rect 13290 1480 13310 1520
rect 13680 1520 13910 1540
rect 13680 1510 13850 1520
rect 13230 1460 13310 1480
rect 13830 1480 13850 1510
rect 13890 1480 13910 1520
rect 13830 1460 13910 1480
rect 12480 1430 12510 1460
rect 13080 1430 13110 1460
rect 13680 1430 13710 1460
rect 8540 1400 8570 1430
rect 8650 1410 8680 1430
rect 8760 1410 8790 1430
rect 8870 1410 8900 1430
rect 9200 1410 9230 1430
rect 8520 1380 8600 1400
rect 8520 1340 8540 1380
rect 8580 1340 8600 1380
rect 2810 1290 2890 1310
rect 2810 1250 2830 1290
rect 2870 1250 2890 1290
rect 2810 1230 2890 1250
rect 2940 1230 2970 1340
rect 3050 1310 3080 1340
rect 3160 1310 3190 1340
rect 3270 1310 3300 1340
rect 3050 1290 3470 1310
rect 3050 1280 3410 1290
rect 2600 1180 2760 1210
rect 2940 1210 3090 1230
rect 2940 1200 3030 1210
rect 2490 1120 2520 1150
rect 2600 1120 2630 1180
rect 1760 1090 1840 1110
rect 1760 1050 1780 1090
rect 1820 1050 1840 1090
rect 1760 1030 1840 1050
rect 2070 990 2100 1020
rect 2490 990 2520 1020
rect 2600 990 2630 1020
rect 2730 1010 2760 1180
rect 3010 1170 3030 1200
rect 3070 1170 3090 1210
rect 3010 1150 3090 1170
rect 3160 1120 3190 1280
rect 3390 1250 3410 1280
rect 3450 1250 3470 1290
rect 3390 1240 3470 1250
rect 3410 1180 3490 1190
rect 3270 1170 3490 1180
rect 3270 1150 3430 1170
rect 3270 1120 3300 1150
rect 3410 1130 3430 1150
rect 3470 1130 3490 1170
rect 3410 1110 3490 1130
rect 3600 1120 3630 1340
rect 3710 1120 3740 1340
rect 3820 1120 3850 1340
rect 3930 1310 3960 1340
rect 4280 1310 4310 1340
rect 4390 1320 4420 1340
rect 4500 1320 4530 1340
rect 4610 1320 4640 1340
rect 4860 1320 4890 1340
rect 4390 1310 4890 1320
rect 3910 1290 4140 1310
rect 3910 1250 3930 1290
rect 3970 1280 4140 1290
rect 3970 1250 3990 1280
rect 3910 1240 3990 1250
rect 4110 1190 4140 1280
rect 4260 1290 4340 1310
rect 4390 1290 4920 1310
rect 4260 1250 4280 1290
rect 4320 1250 4340 1290
rect 4260 1240 4340 1250
rect 4440 1190 4470 1290
rect 4840 1250 4860 1290
rect 4900 1250 4920 1290
rect 4840 1230 4920 1250
rect 4110 1160 4470 1190
rect 4440 1120 4470 1160
rect 4970 1190 5000 1340
rect 5050 1290 5130 1310
rect 5050 1250 5070 1290
rect 5110 1280 5130 1290
rect 5290 1290 5370 1310
rect 5290 1280 5310 1290
rect 5110 1250 5310 1280
rect 5350 1250 5370 1290
rect 5050 1240 5130 1250
rect 5290 1230 5370 1250
rect 4970 1170 5190 1190
rect 5420 1170 5450 1340
rect 5630 1280 5710 1300
rect 5630 1240 5650 1280
rect 5690 1240 5710 1280
rect 5630 1220 5710 1240
rect 5780 1240 5810 1340
rect 5900 1240 5980 1260
rect 5780 1210 5920 1240
rect 5780 1170 5810 1210
rect 5900 1200 5920 1210
rect 5960 1200 5980 1240
rect 6030 1230 6060 1340
rect 6140 1310 6170 1340
rect 6250 1310 6280 1340
rect 6360 1310 6390 1340
rect 6140 1290 6610 1310
rect 6140 1280 6550 1290
rect 6030 1210 6180 1230
rect 6030 1200 6120 1210
rect 5900 1180 5980 1200
rect 4970 1160 5130 1170
rect 4860 1120 4890 1150
rect 4970 1120 5000 1160
rect 5110 1130 5130 1160
rect 5170 1130 5190 1170
rect 5110 1110 5190 1130
rect 5310 1140 5450 1170
rect 5310 1120 5340 1140
rect 5420 1120 5450 1140
rect 5670 1140 5810 1170
rect 6100 1170 6120 1200
rect 6160 1170 6180 1210
rect 6100 1150 6180 1170
rect 5670 1120 5700 1140
rect 5780 1120 5810 1140
rect 6250 1120 6280 1280
rect 6530 1250 6550 1280
rect 6590 1250 6610 1290
rect 6530 1240 6610 1250
rect 6500 1180 6580 1190
rect 6360 1170 6580 1180
rect 6360 1150 6520 1170
rect 6360 1120 6390 1150
rect 6500 1130 6520 1150
rect 6560 1130 6580 1170
rect 6500 1110 6580 1130
rect 6690 1120 6720 1340
rect 6800 1190 6830 1340
rect 6910 1310 6940 1340
rect 7240 1310 7270 1340
rect 7350 1320 7380 1340
rect 7460 1320 7490 1340
rect 7570 1320 7600 1340
rect 7900 1320 7930 1340
rect 6890 1290 7100 1310
rect 6890 1250 6910 1290
rect 6950 1280 7100 1290
rect 6950 1250 6970 1280
rect 6890 1240 6970 1250
rect 7070 1190 7100 1280
rect 7220 1290 7300 1310
rect 7220 1250 7240 1290
rect 7280 1250 7300 1290
rect 7220 1240 7300 1250
rect 7350 1290 7930 1320
rect 7350 1190 7380 1290
rect 7800 1250 7820 1290
rect 7860 1250 7880 1290
rect 7800 1230 7880 1250
rect 8010 1230 8040 1340
rect 6800 1160 6960 1190
rect 7070 1160 7380 1190
rect 7630 1210 7710 1230
rect 7630 1170 7650 1210
rect 7690 1170 7710 1210
rect 7930 1200 8040 1230
rect 8120 1260 8150 1340
rect 8520 1320 8600 1340
rect 8650 1380 9230 1410
rect 8270 1270 8350 1290
rect 8270 1260 8290 1270
rect 8120 1230 8290 1260
rect 8330 1230 8350 1270
rect 7930 1170 7960 1200
rect 6800 1120 6830 1160
rect 6930 1110 6960 1160
rect 7310 1120 7340 1160
rect 7630 1150 7710 1170
rect 7650 1120 7680 1150
rect 7760 1140 7960 1170
rect 7760 1120 7790 1140
rect 8010 1120 8040 1150
rect 8120 1120 8150 1230
rect 8270 1210 8350 1230
rect 8650 1180 8680 1380
rect 9100 1340 9120 1380
rect 9160 1340 9180 1380
rect 9100 1320 9180 1340
rect 9310 1260 9340 1430
rect 9060 1230 9340 1260
rect 9420 1260 9450 1430
rect 9840 1400 9870 1430
rect 9950 1410 9980 1430
rect 10060 1410 10090 1430
rect 10170 1410 10200 1430
rect 10500 1410 10530 1430
rect 9820 1380 9900 1400
rect 9820 1340 9840 1380
rect 9880 1340 9900 1380
rect 9820 1320 9900 1340
rect 9950 1380 10530 1410
rect 9570 1270 9650 1290
rect 9570 1260 9590 1270
rect 9420 1230 9590 1260
rect 9630 1230 9650 1270
rect 8610 1150 8680 1180
rect 8930 1210 9010 1230
rect 8930 1170 8950 1210
rect 8990 1170 9010 1210
rect 8930 1150 9010 1170
rect 8610 1120 8640 1150
rect 8950 1120 8980 1150
rect 9060 1120 9090 1230
rect 9310 1120 9340 1150
rect 9420 1120 9450 1230
rect 9570 1210 9650 1230
rect 9950 1180 9980 1380
rect 10400 1340 10420 1380
rect 10460 1340 10480 1380
rect 10400 1320 10480 1340
rect 10610 1260 10640 1430
rect 10360 1230 10640 1260
rect 10720 1260 10750 1430
rect 11140 1400 11170 1430
rect 11250 1410 11280 1430
rect 11360 1410 11390 1430
rect 11470 1410 11500 1430
rect 11800 1410 11830 1430
rect 11120 1380 11200 1400
rect 11120 1340 11140 1380
rect 11180 1340 11200 1380
rect 11120 1320 11200 1340
rect 11250 1380 11830 1410
rect 10870 1270 10950 1290
rect 10870 1260 10890 1270
rect 10720 1230 10890 1260
rect 10930 1230 10950 1270
rect 9910 1150 9980 1180
rect 10230 1210 10310 1230
rect 10230 1170 10250 1210
rect 10290 1170 10310 1210
rect 10230 1150 10310 1170
rect 9910 1120 9940 1150
rect 10250 1120 10280 1150
rect 10360 1120 10390 1230
rect 10610 1120 10640 1150
rect 10720 1120 10750 1230
rect 10870 1210 10950 1230
rect 11250 1180 11280 1380
rect 11700 1340 11720 1380
rect 11760 1340 11780 1380
rect 11700 1320 11780 1340
rect 11910 1260 11940 1430
rect 11660 1230 11940 1260
rect 12020 1260 12050 1430
rect 12290 1290 12370 1310
rect 12480 1290 12510 1330
rect 12290 1260 12310 1290
rect 12020 1250 12310 1260
rect 12350 1260 12510 1290
rect 12350 1250 12370 1260
rect 12020 1230 12370 1250
rect 11210 1150 11280 1180
rect 11530 1210 11610 1230
rect 11530 1170 11550 1210
rect 11590 1170 11610 1210
rect 11530 1150 11610 1170
rect 11210 1120 11240 1150
rect 11550 1120 11580 1150
rect 11660 1120 11690 1230
rect 11910 1120 11940 1150
rect 12020 1120 12050 1230
rect 12480 1220 12510 1260
rect 12890 1290 12970 1310
rect 13080 1290 13110 1330
rect 12890 1250 12910 1290
rect 12950 1260 13110 1290
rect 12950 1250 12970 1260
rect 12890 1230 12970 1250
rect 13080 1220 13110 1260
rect 13490 1290 13570 1310
rect 13680 1290 13710 1330
rect 13490 1250 13510 1290
rect 13550 1260 13710 1290
rect 13550 1250 13570 1260
rect 13490 1230 13570 1250
rect 13680 1220 13710 1260
rect 6930 1090 7170 1110
rect 6930 1080 7110 1090
rect 7090 1050 7110 1080
rect 7150 1050 7170 1090
rect 7090 1030 7170 1050
rect 2730 990 2810 1010
rect 3160 990 3190 1020
rect 3270 990 3300 1020
rect 3600 990 3630 1020
rect 3710 990 3740 1020
rect 3820 990 3850 1020
rect 4440 990 4470 1020
rect 4860 990 4890 1020
rect 4970 990 5000 1020
rect 5310 990 5340 1020
rect 5420 990 5450 1020
rect 5670 990 5700 1020
rect 5780 990 5810 1020
rect 6250 990 6280 1020
rect 6360 990 6390 1020
rect 2420 970 2520 990
rect 2420 930 2440 970
rect 2480 930 2520 970
rect 2730 950 2750 990
rect 2790 950 2810 990
rect 2730 930 2810 950
rect 3540 970 3630 990
rect 3540 930 3560 970
rect 3600 930 3630 970
rect 2420 910 2520 930
rect 3540 910 3630 930
rect 3680 970 3740 990
rect 3680 930 3690 970
rect 3730 930 3740 970
rect 3680 910 3740 930
rect 4800 970 4890 990
rect 6690 980 6720 1020
rect 6800 990 6830 1020
rect 7310 990 7340 1020
rect 7650 990 7680 1020
rect 7760 990 7790 1020
rect 8010 1000 8040 1020
rect 8120 1000 8150 1020
rect 4800 930 4820 970
rect 4860 930 4890 970
rect 4800 910 4890 930
rect 6560 960 6720 980
rect 8010 970 8150 1000
rect 8610 990 8640 1020
rect 8950 990 8980 1020
rect 9060 990 9090 1020
rect 9310 1000 9340 1020
rect 9420 1000 9450 1020
rect 9060 970 9170 990
rect 9310 970 9450 1000
rect 9910 990 9940 1020
rect 10250 990 10280 1020
rect 10360 990 10390 1020
rect 10610 1000 10640 1020
rect 10720 1000 10750 1020
rect 10360 970 10470 990
rect 10610 970 10750 1000
rect 11210 990 11240 1020
rect 11550 990 11580 1020
rect 11660 990 11690 1020
rect 11910 1000 11940 1020
rect 12020 1000 12050 1020
rect 11660 970 11770 990
rect 11910 970 12050 1000
rect 12480 990 12510 1020
rect 13080 990 13110 1020
rect 13680 990 13710 1020
rect 12700 970 12780 990
rect 6560 920 6580 960
rect 6620 950 6720 960
rect 6620 920 6640 950
rect 6560 910 6640 920
rect 9060 930 9110 970
rect 9150 930 9170 970
rect 9060 910 9170 930
rect 10360 930 10410 970
rect 10450 930 10470 970
rect 10360 910 10470 930
rect 11660 930 11710 970
rect 11750 930 11770 970
rect 12700 940 12720 970
rect 11660 910 11770 930
rect 12480 930 12720 940
rect 12760 930 12780 970
rect 13300 970 13380 990
rect 13300 940 13320 970
rect 12480 910 12780 930
rect 13080 930 13320 940
rect 13360 930 13380 970
rect 13900 970 13980 990
rect 13900 940 13920 970
rect 13080 910 13380 930
rect 13680 930 13920 940
rect 13960 930 13980 970
rect 13680 910 13980 930
rect 12480 880 12510 910
rect 13080 880 13110 910
rect 13680 880 13710 910
rect 12480 650 12510 680
rect 13080 650 13110 680
rect 13680 650 13710 680
rect 14220 620 14280 640
rect 14220 600 14230 620
rect 12480 580 14230 600
rect 14270 580 14280 620
rect 12480 560 14280 580
rect 14340 620 14400 640
rect 14340 580 14350 620
rect 14390 580 14400 620
rect 14340 560 14400 580
rect 14460 620 14520 640
rect 14460 580 14470 620
rect 14510 580 14520 620
rect 14460 560 14520 580
rect 12480 530 12780 560
rect 13080 530 13380 560
rect 13680 530 13980 560
rect 14220 530 14520 560
rect 12480 100 12780 130
rect 13080 100 13380 130
rect 13680 100 13980 130
rect 14220 100 14520 130
<< polycont >>
rect 1330 10000 1370 10040
rect 1490 10000 1530 10040
rect 1650 10000 1690 10040
rect 1810 10000 1850 10040
rect 1970 10000 2010 10040
rect 2130 10000 2170 10040
rect 2290 10000 2330 10040
rect 2450 10000 2490 10040
rect 2610 10000 2650 10040
rect 2770 10000 2810 10040
rect 2930 10000 2970 10040
rect 3090 10000 3130 10040
rect 3410 10000 3450 10040
rect 3570 10000 3610 10040
rect 3730 10000 3770 10040
rect 3890 10000 3930 10040
rect 4050 10000 4090 10040
rect 4210 10000 4250 10040
rect 4370 10000 4410 10040
rect 4530 10000 4570 10040
rect 4690 10000 4730 10040
rect 4850 10000 4890 10040
rect 5010 10000 5050 10040
rect 5170 10000 5210 10040
rect 930 9090 970 9130
rect 1170 9090 1210 9130
rect 1410 9090 1450 9130
rect 1650 9090 1690 9130
rect 2290 9090 2330 9130
rect 2530 9090 2570 9130
rect 2770 9090 2810 9130
rect 3730 9090 3770 9130
rect 3970 9090 4010 9130
rect 4210 9090 4250 9130
rect 4850 9090 4890 9130
rect 5090 9090 5130 9130
rect 5330 9090 5370 9130
rect 5570 9090 5610 9130
rect 7856 8836 7890 8870
rect 9130 8836 9164 8870
rect 1433 8718 1467 8752
rect 1793 8718 1827 8752
rect 1913 8718 1947 8752
rect 2273 8718 2307 8752
rect 2393 8718 2427 8752
rect 1534 8488 1568 8522
rect 1692 8488 1726 8522
rect 2016 8488 2050 8522
rect 2170 8488 2204 8522
rect 2494 8488 2528 8522
rect 4113 8718 4147 8752
rect 4233 8718 4267 8752
rect 4593 8718 4627 8752
rect 4713 8718 4747 8752
rect 5073 8718 5107 8752
rect 9030 8660 9070 8700
rect 9430 8660 9470 8700
rect 4012 8488 4046 8522
rect 4336 8488 4370 8522
rect 4490 8488 4524 8522
rect 4814 8488 4848 8522
rect 4972 8488 5006 8522
rect 8230 8270 8270 8310
rect 10230 8270 10270 8310
rect 8340 7970 8390 8020
rect 8990 7970 9040 8020
rect 9480 7970 9520 8010
rect 10140 7970 10180 8010
rect 10620 7970 10660 8010
rect 11280 7970 11320 8010
rect 710 7890 750 7930
rect 890 7880 930 7920
rect 1370 7880 1410 7920
rect 1610 7880 1650 7920
rect 2090 7880 2130 7920
rect 2330 7880 2370 7920
rect 2750 7880 2790 7920
rect 3750 7880 3790 7920
rect 4170 7880 4210 7920
rect 4410 7880 4450 7920
rect 4890 7880 4930 7920
rect 5130 7880 5170 7920
rect 5610 7880 5650 7920
rect 5790 7890 5830 7930
rect 8540 7730 8580 7770
rect 9590 7730 9630 7770
rect 10030 7710 10070 7750
rect 11570 7730 11610 7770
rect 10730 7610 10770 7650
rect 530 7540 570 7580
rect 2930 7540 2970 7580
rect 3570 7540 3610 7580
rect 5970 7540 6010 7580
rect 8450 7400 8490 7440
rect 8890 7400 8930 7440
rect 9680 7410 9720 7450
rect 10730 7400 10770 7440
rect 11570 7400 11610 7440
rect 8340 7060 8380 7100
rect 9000 7060 9040 7100
rect 9480 7060 9520 7100
rect 10140 7060 10180 7100
rect 10620 7060 10660 7100
rect 11280 7060 11320 7100
rect 1900 6720 1940 6760
rect 2080 6720 2120 6760
rect 2260 6720 2300 6760
rect 2440 6720 2480 6760
rect 2620 6720 2660 6760
rect 2800 6720 2840 6760
rect 2980 6720 3020 6760
rect 3160 6720 3200 6760
rect 3340 6720 3380 6760
rect 3520 6720 3560 6760
rect 3700 6720 3740 6760
rect 3880 6720 3920 6760
rect 4060 6720 4100 6760
rect 4240 6720 4280 6760
rect 4420 6720 4460 6760
rect 4600 6720 4640 6760
rect 8350 6750 8390 6790
rect 10350 6750 10390 6790
rect 5720 6520 5760 6560
rect 5500 6180 5540 6220
rect 5940 6180 5980 6220
rect 9150 6110 9190 6150
rect 9550 6110 9590 6150
rect 1630 5980 1670 6020
rect 4870 5980 4910 6020
rect 1808 5718 1842 5752
rect 1918 5718 1952 5752
rect 2028 5718 2062 5752
rect 2138 5718 2172 5752
rect 2248 5718 2282 5752
rect 2358 5718 2392 5752
rect 2468 5718 2502 5752
rect 2578 5718 2612 5752
rect 2688 5718 2722 5752
rect 2798 5718 2832 5752
rect 3708 5718 3742 5752
rect 3818 5718 3852 5752
rect 3928 5718 3962 5752
rect 4038 5718 4072 5752
rect 4148 5718 4182 5752
rect 4258 5718 4292 5752
rect 4368 5718 4402 5752
rect 4478 5718 4512 5752
rect 4588 5718 4622 5752
rect 4698 5718 4732 5752
rect 1640 5380 1680 5420
rect 2960 5380 3000 5420
rect 3540 5380 3580 5420
rect 4860 5380 4900 5420
rect 4290 4780 4330 4820
rect 1950 4430 1990 4470
rect 2370 4440 2410 4480
rect 2890 4360 2930 4400
rect 3270 4440 3310 4480
rect 2490 3940 2530 3980
rect 3860 4430 3900 4470
rect 4370 4390 4410 4430
rect 4700 4390 4740 4430
rect 5030 4390 5070 4430
rect 5160 4420 5200 4460
rect 5730 4390 5770 4430
rect 6120 4440 6160 4480
rect 6250 4360 6290 4400
rect 6660 4360 6700 4400
rect 8170 4410 8210 4450
rect 11010 4410 11050 4450
rect 3390 3940 3430 3980
rect 4160 3820 4200 3860
rect 8480 3840 8520 3880
rect 9590 3870 9630 3910
rect 10000 3840 10040 3880
rect 10700 3840 10740 3880
rect 2610 3600 2650 3640
rect 5730 3600 5770 3640
rect 8410 3560 8450 3600
rect 2490 3480 2530 3520
rect 2040 2990 2080 3030
rect 2370 2980 2410 3020
rect 3390 3480 3430 3520
rect 2890 3060 2930 3100
rect 3270 2980 3310 3020
rect 8950 3430 8990 3470
rect 10030 3430 10070 3470
rect 10440 3460 10480 3500
rect 10700 3460 10740 3500
rect 3880 3030 3920 3070
rect 4040 3030 4080 3070
rect 4370 3030 4410 3070
rect 4700 3030 4740 3070
rect 4960 3030 5000 3070
rect 5160 3020 5200 3060
rect 5860 3050 5900 3090
rect 6250 2970 6290 3010
rect 7970 2890 8010 2930
rect 11010 2890 11050 2930
rect 5810 2640 5850 2680
rect 6450 2640 6490 2680
rect 14320 1770 14360 1810
rect 1800 1490 1840 1530
rect 2750 1470 2790 1510
rect 3820 1480 3860 1520
rect 5380 1480 5420 1520
rect 7984 1490 8024 1530
rect 1910 1250 1950 1290
rect 2490 1250 2530 1290
rect 12650 1480 12690 1520
rect 13250 1480 13290 1520
rect 13850 1480 13890 1520
rect 8540 1340 8580 1380
rect 2830 1250 2870 1290
rect 1780 1050 1820 1090
rect 3030 1170 3070 1210
rect 3410 1250 3450 1290
rect 3430 1130 3470 1170
rect 3930 1250 3970 1290
rect 4280 1250 4320 1290
rect 4860 1250 4900 1290
rect 5070 1250 5110 1290
rect 5310 1250 5350 1290
rect 5650 1240 5690 1280
rect 5920 1200 5960 1240
rect 5130 1130 5170 1170
rect 6120 1170 6160 1210
rect 6550 1250 6590 1290
rect 6520 1130 6560 1170
rect 6910 1250 6950 1290
rect 7240 1250 7280 1290
rect 7820 1250 7860 1290
rect 7650 1170 7690 1210
rect 8290 1230 8330 1270
rect 9120 1340 9160 1380
rect 9840 1340 9880 1380
rect 9590 1230 9630 1270
rect 8950 1170 8990 1210
rect 10420 1340 10460 1380
rect 11140 1340 11180 1380
rect 10890 1230 10930 1270
rect 10250 1170 10290 1210
rect 11720 1340 11760 1380
rect 12310 1250 12350 1290
rect 11550 1170 11590 1210
rect 12910 1250 12950 1290
rect 13510 1250 13550 1290
rect 7110 1050 7150 1090
rect 2440 930 2480 970
rect 2750 950 2790 990
rect 3560 930 3600 970
rect 3690 930 3730 970
rect 4820 930 4860 970
rect 6580 920 6620 960
rect 9110 930 9150 970
rect 10410 930 10450 970
rect 11710 930 11750 970
rect 12720 930 12760 970
rect 13320 930 13360 970
rect 13920 930 13960 970
rect 14230 580 14270 620
rect 14350 580 14390 620
rect 14470 580 14510 620
<< xpolycontact >>
rect 120 13680 190 14118
rect 120 12862 190 13302
rect 240 13888 310 14328
rect 240 12810 310 13250
rect 360 13888 430 14328
rect 360 12810 430 13250
rect 480 13888 550 14328
rect 480 12810 550 13250
rect 670 14038 740 14478
rect 670 12430 740 12870
rect 790 14038 860 14478
rect 790 12430 860 12870
rect 910 14038 980 14478
rect 5440 14038 5510 14478
rect 910 12430 980 12870
rect 5440 12430 5510 12870
rect 5560 14038 5630 14478
rect 5560 12430 5630 12870
rect 5680 14038 5750 14478
rect 5800 13888 5870 14328
rect 5800 13280 5870 13720
rect 6460 13890 6530 14328
rect 6460 13072 6530 13512
rect 5680 12430 5750 12870
rect 2622 10550 3062 10620
rect 3490 10550 3930 10620
rect 11640 8960 11710 9400
rect 11640 8380 11710 8820
rect 11640 6670 11710 7110
rect 11640 6034 11710 6474
rect 23180 2440 23620 2510
rect 25092 2440 25532 2510
<< npolyres >>
rect 8270 8820 8750 8886
<< ppolyres >>
rect 120 13302 190 13680
rect 6460 13512 6530 13890
<< xpolyres >>
rect 240 13250 310 13888
rect 360 13250 430 13888
rect 480 13250 550 13888
rect 670 12870 740 14038
rect 790 12870 860 14038
rect 910 12870 980 14038
rect 5440 12870 5510 14038
rect 5560 12870 5630 14038
rect 5680 12870 5750 14038
rect 5800 13720 5870 13888
rect 3062 10550 3490 10620
rect 11640 8820 11710 8960
rect 11640 6474 11710 6670
rect 23620 2440 25092 2510
<< locali >>
rect 3230 15080 3310 15100
rect 3230 15040 3250 15080
rect 3290 15040 3310 15080
rect 3230 15000 3310 15040
rect 3230 14960 3250 15000
rect 3290 14960 3310 15000
rect 3230 14920 3310 14960
rect 3230 14880 3250 14920
rect 3290 14880 3310 14920
rect 2550 14794 2630 14800
rect 3230 14794 3310 14880
rect 3910 14794 3990 14800
rect 1266 14762 5274 14794
rect 1266 14728 1400 14762
rect 1434 14728 1490 14762
rect 1524 14728 1580 14762
rect 1614 14728 1670 14762
rect 1704 14728 1760 14762
rect 1794 14728 1850 14762
rect 1884 14728 1940 14762
rect 1974 14728 2030 14762
rect 2064 14728 2120 14762
rect 2154 14728 2210 14762
rect 2244 14728 2300 14762
rect 2334 14728 2390 14762
rect 2424 14728 2760 14762
rect 2794 14728 2850 14762
rect 2884 14728 2940 14762
rect 2974 14728 3030 14762
rect 3064 14728 3120 14762
rect 3154 14728 3210 14762
rect 3244 14728 3300 14762
rect 3334 14728 3390 14762
rect 3424 14728 3480 14762
rect 3514 14728 3570 14762
rect 3604 14728 3660 14762
rect 3694 14728 3750 14762
rect 3784 14728 4120 14762
rect 4154 14728 4210 14762
rect 4244 14728 4300 14762
rect 4334 14728 4390 14762
rect 4424 14728 4480 14762
rect 4514 14728 4570 14762
rect 4604 14728 4660 14762
rect 4694 14728 4750 14762
rect 4784 14728 4840 14762
rect 4874 14728 4930 14762
rect 4964 14728 5020 14762
rect 5054 14728 5110 14762
rect 5144 14728 5274 14762
rect 1266 14695 5274 14728
rect 1266 14678 1365 14695
rect 1266 14644 1299 14678
rect 1333 14644 1365 14678
rect 1266 14588 1365 14644
rect 2455 14678 2725 14695
rect 2455 14644 2486 14678
rect 2520 14644 2659 14678
rect 2693 14644 2725 14678
rect 910 14548 980 14568
rect 910 14498 920 14548
rect 970 14498 980 14548
rect 910 14478 980 14498
rect 480 14398 550 14418
rect 480 14348 490 14398
rect 540 14348 550 14398
rect 480 14328 550 14348
rect 120 14188 190 14208
rect 120 14138 130 14188
rect 180 14138 190 14188
rect 120 14118 190 14138
rect 310 14258 360 14328
rect 740 14408 790 14478
rect 1266 14554 1299 14588
rect 1333 14554 1365 14588
rect 1266 14498 1365 14554
rect 1266 14464 1299 14498
rect 1333 14464 1365 14498
rect 1266 14408 1365 14464
rect 1266 14374 1299 14408
rect 1333 14374 1365 14408
rect 1266 14318 1365 14374
rect 1266 14284 1299 14318
rect 1333 14284 1365 14318
rect 1266 14228 1365 14284
rect 1266 14194 1299 14228
rect 1333 14194 1365 14228
rect 1266 14138 1365 14194
rect 1266 14104 1299 14138
rect 1333 14104 1365 14138
rect 1266 14048 1365 14104
rect 1266 14014 1299 14048
rect 1333 14014 1365 14048
rect 1266 13958 1365 14014
rect 1266 13924 1299 13958
rect 1333 13924 1365 13958
rect 1266 13868 1365 13924
rect 1266 13834 1299 13868
rect 1333 13834 1365 13868
rect 1266 13778 1365 13834
rect 1266 13750 1299 13778
rect 1260 13744 1299 13750
rect 1333 13750 1365 13778
rect 1429 14612 2391 14631
rect 1429 14578 1540 14612
rect 1574 14578 1630 14612
rect 1664 14578 1720 14612
rect 1754 14578 1810 14612
rect 1844 14578 1900 14612
rect 1934 14578 1990 14612
rect 2024 14578 2080 14612
rect 2114 14578 2170 14612
rect 2204 14578 2260 14612
rect 2294 14578 2391 14612
rect 1429 14559 2391 14578
rect 1429 14518 1501 14559
rect 1429 14484 1448 14518
rect 1482 14484 1501 14518
rect 2319 14499 2391 14559
rect 1429 14428 1501 14484
rect 1429 14394 1448 14428
rect 1482 14394 1501 14428
rect 1429 14338 1501 14394
rect 1429 14304 1448 14338
rect 1482 14304 1501 14338
rect 1429 14248 1501 14304
rect 1429 14214 1448 14248
rect 1482 14214 1501 14248
rect 1429 14158 1501 14214
rect 1429 14124 1448 14158
rect 1482 14124 1501 14158
rect 1429 14068 1501 14124
rect 1429 14034 1448 14068
rect 1482 14034 1501 14068
rect 1429 13978 1501 14034
rect 1429 13944 1448 13978
rect 1482 13944 1501 13978
rect 1429 13888 1501 13944
rect 1429 13854 1448 13888
rect 1482 13854 1501 13888
rect 1429 13798 1501 13854
rect 1563 14436 2257 14497
rect 1563 14402 1622 14436
rect 1656 14424 1712 14436
rect 1684 14402 1712 14424
rect 1746 14424 1802 14436
rect 1746 14402 1750 14424
rect 1563 14390 1650 14402
rect 1684 14390 1750 14402
rect 1784 14402 1802 14424
rect 1836 14424 1892 14436
rect 1836 14402 1850 14424
rect 1784 14390 1850 14402
rect 1884 14402 1892 14424
rect 1926 14424 1982 14436
rect 2016 14424 2072 14436
rect 2106 14424 2162 14436
rect 1926 14402 1950 14424
rect 2016 14402 2050 14424
rect 2106 14402 2150 14424
rect 2196 14402 2257 14436
rect 1884 14390 1950 14402
rect 1984 14390 2050 14402
rect 2084 14390 2150 14402
rect 2184 14390 2257 14402
rect 1563 14346 2257 14390
rect 1563 14312 1622 14346
rect 1656 14324 1712 14346
rect 1684 14312 1712 14324
rect 1746 14324 1802 14346
rect 1746 14312 1750 14324
rect 1563 14290 1650 14312
rect 1684 14290 1750 14312
rect 1784 14312 1802 14324
rect 1836 14324 1892 14346
rect 1836 14312 1850 14324
rect 1784 14290 1850 14312
rect 1884 14312 1892 14324
rect 1926 14324 1982 14346
rect 2016 14324 2072 14346
rect 2106 14324 2162 14346
rect 1926 14312 1950 14324
rect 2016 14312 2050 14324
rect 2106 14312 2150 14324
rect 2196 14312 2257 14346
rect 1884 14290 1950 14312
rect 1984 14290 2050 14312
rect 2084 14290 2150 14312
rect 2184 14290 2257 14312
rect 1563 14256 2257 14290
rect 1563 14222 1622 14256
rect 1656 14224 1712 14256
rect 1684 14222 1712 14224
rect 1746 14224 1802 14256
rect 1746 14222 1750 14224
rect 1563 14190 1650 14222
rect 1684 14190 1750 14222
rect 1784 14222 1802 14224
rect 1836 14224 1892 14256
rect 1836 14222 1850 14224
rect 1784 14190 1850 14222
rect 1884 14222 1892 14224
rect 1926 14224 1982 14256
rect 2016 14224 2072 14256
rect 2106 14224 2162 14256
rect 1926 14222 1950 14224
rect 2016 14222 2050 14224
rect 2106 14222 2150 14224
rect 2196 14222 2257 14256
rect 1884 14190 1950 14222
rect 1984 14190 2050 14222
rect 2084 14190 2150 14222
rect 2184 14190 2257 14222
rect 1563 14166 2257 14190
rect 1563 14132 1622 14166
rect 1656 14132 1712 14166
rect 1746 14132 1802 14166
rect 1836 14132 1892 14166
rect 1926 14132 1982 14166
rect 2016 14132 2072 14166
rect 2106 14132 2162 14166
rect 2196 14132 2257 14166
rect 1563 14124 2257 14132
rect 1563 14090 1650 14124
rect 1684 14090 1750 14124
rect 1784 14090 1850 14124
rect 1884 14090 1950 14124
rect 1984 14090 2050 14124
rect 2084 14090 2150 14124
rect 2184 14090 2257 14124
rect 1563 14076 2257 14090
rect 1563 14042 1622 14076
rect 1656 14042 1712 14076
rect 1746 14042 1802 14076
rect 1836 14042 1892 14076
rect 1926 14042 1982 14076
rect 2016 14042 2072 14076
rect 2106 14042 2162 14076
rect 2196 14042 2257 14076
rect 1563 14024 2257 14042
rect 1563 13990 1650 14024
rect 1684 13990 1750 14024
rect 1784 13990 1850 14024
rect 1884 13990 1950 14024
rect 1984 13990 2050 14024
rect 2084 13990 2150 14024
rect 2184 13990 2257 14024
rect 1563 13986 2257 13990
rect 1563 13952 1622 13986
rect 1656 13952 1712 13986
rect 1746 13952 1802 13986
rect 1836 13952 1892 13986
rect 1926 13952 1982 13986
rect 2016 13952 2072 13986
rect 2106 13952 2162 13986
rect 2196 13952 2257 13986
rect 1563 13924 2257 13952
rect 1563 13896 1650 13924
rect 1684 13896 1750 13924
rect 1563 13862 1622 13896
rect 1684 13890 1712 13896
rect 1656 13862 1712 13890
rect 1746 13890 1750 13896
rect 1784 13896 1850 13924
rect 1784 13890 1802 13896
rect 1746 13862 1802 13890
rect 1836 13890 1850 13896
rect 1884 13896 1950 13924
rect 1984 13896 2050 13924
rect 2084 13896 2150 13924
rect 2184 13896 2257 13924
rect 1884 13890 1892 13896
rect 1836 13862 1892 13890
rect 1926 13890 1950 13896
rect 2016 13890 2050 13896
rect 2106 13890 2150 13896
rect 1926 13862 1982 13890
rect 2016 13862 2072 13890
rect 2106 13862 2162 13890
rect 2196 13862 2257 13896
rect 1563 13803 2257 13862
rect 2319 14465 2338 14499
rect 2372 14465 2391 14499
rect 2319 14409 2391 14465
rect 2319 14375 2338 14409
rect 2372 14375 2391 14409
rect 2319 14319 2391 14375
rect 2319 14285 2338 14319
rect 2372 14285 2391 14319
rect 2319 14229 2391 14285
rect 2319 14195 2338 14229
rect 2372 14195 2391 14229
rect 2319 14139 2391 14195
rect 2319 14105 2338 14139
rect 2372 14105 2391 14139
rect 2319 14049 2391 14105
rect 2319 14015 2338 14049
rect 2372 14015 2391 14049
rect 2319 13959 2391 14015
rect 2319 13925 2338 13959
rect 2372 13925 2391 13959
rect 2319 13869 2391 13925
rect 2319 13835 2338 13869
rect 2372 13835 2391 13869
rect 1429 13764 1448 13798
rect 1482 13764 1501 13798
rect 1429 13750 1501 13764
rect 2319 13779 2391 13835
rect 2319 13750 2338 13779
rect 1333 13745 2338 13750
rect 2372 13750 2391 13779
rect 2455 14588 2725 14644
rect 3815 14678 4085 14695
rect 3815 14644 3846 14678
rect 3880 14644 4019 14678
rect 4053 14644 4085 14678
rect 2455 14554 2486 14588
rect 2520 14554 2659 14588
rect 2693 14554 2725 14588
rect 2455 14498 2725 14554
rect 2455 14464 2486 14498
rect 2520 14464 2659 14498
rect 2693 14464 2725 14498
rect 2455 14408 2725 14464
rect 2455 14374 2486 14408
rect 2520 14374 2659 14408
rect 2693 14374 2725 14408
rect 2455 14318 2725 14374
rect 2455 14284 2486 14318
rect 2520 14284 2659 14318
rect 2693 14284 2725 14318
rect 2455 14228 2725 14284
rect 2455 14194 2486 14228
rect 2520 14194 2659 14228
rect 2693 14194 2725 14228
rect 2455 14138 2725 14194
rect 2455 14104 2486 14138
rect 2520 14104 2659 14138
rect 2693 14104 2725 14138
rect 2455 14048 2725 14104
rect 2455 14014 2486 14048
rect 2520 14014 2659 14048
rect 2693 14014 2725 14048
rect 2455 13958 2725 14014
rect 2455 13924 2486 13958
rect 2520 13924 2659 13958
rect 2693 13924 2725 13958
rect 2455 13868 2725 13924
rect 2455 13834 2486 13868
rect 2520 13834 2659 13868
rect 2693 13834 2725 13868
rect 2455 13778 2725 13834
rect 2455 13750 2486 13778
rect 2372 13745 2486 13750
rect 1333 13744 2486 13745
rect 2520 13744 2659 13778
rect 2693 13750 2725 13778
rect 2789 14612 3751 14631
rect 2789 14578 2900 14612
rect 2934 14578 2990 14612
rect 3024 14578 3080 14612
rect 3114 14578 3170 14612
rect 3204 14578 3260 14612
rect 3294 14578 3350 14612
rect 3384 14578 3440 14612
rect 3474 14578 3530 14612
rect 3564 14578 3620 14612
rect 3654 14578 3751 14612
rect 2789 14559 3751 14578
rect 2789 14518 2861 14559
rect 2789 14484 2808 14518
rect 2842 14484 2861 14518
rect 3679 14499 3751 14559
rect 2789 14428 2861 14484
rect 2789 14394 2808 14428
rect 2842 14394 2861 14428
rect 2789 14338 2861 14394
rect 2789 14304 2808 14338
rect 2842 14304 2861 14338
rect 2789 14248 2861 14304
rect 2789 14214 2808 14248
rect 2842 14214 2861 14248
rect 2789 14158 2861 14214
rect 2789 14124 2808 14158
rect 2842 14124 2861 14158
rect 2789 14068 2861 14124
rect 2789 14034 2808 14068
rect 2842 14034 2861 14068
rect 2789 13978 2861 14034
rect 2789 13944 2808 13978
rect 2842 13944 2861 13978
rect 2789 13888 2861 13944
rect 2789 13854 2808 13888
rect 2842 13854 2861 13888
rect 2789 13798 2861 13854
rect 2923 14436 3617 14497
rect 2923 14402 2982 14436
rect 3016 14424 3072 14436
rect 3044 14402 3072 14424
rect 3106 14424 3162 14436
rect 3106 14402 3110 14424
rect 2923 14390 3010 14402
rect 3044 14390 3110 14402
rect 3144 14402 3162 14424
rect 3196 14424 3252 14436
rect 3196 14402 3210 14424
rect 3144 14390 3210 14402
rect 3244 14402 3252 14424
rect 3286 14424 3342 14436
rect 3376 14424 3432 14436
rect 3466 14424 3522 14436
rect 3286 14402 3310 14424
rect 3376 14402 3410 14424
rect 3466 14402 3510 14424
rect 3556 14402 3617 14436
rect 3244 14390 3310 14402
rect 3344 14390 3410 14402
rect 3444 14390 3510 14402
rect 3544 14390 3617 14402
rect 2923 14346 3617 14390
rect 2923 14312 2982 14346
rect 3016 14324 3072 14346
rect 3044 14312 3072 14324
rect 3106 14324 3162 14346
rect 3106 14312 3110 14324
rect 2923 14290 3010 14312
rect 3044 14290 3110 14312
rect 3144 14312 3162 14324
rect 3196 14324 3252 14346
rect 3196 14312 3210 14324
rect 3144 14290 3210 14312
rect 3244 14312 3252 14324
rect 3286 14324 3342 14346
rect 3376 14324 3432 14346
rect 3466 14324 3522 14346
rect 3286 14312 3310 14324
rect 3376 14312 3410 14324
rect 3466 14312 3510 14324
rect 3556 14312 3617 14346
rect 3244 14290 3310 14312
rect 3344 14290 3410 14312
rect 3444 14290 3510 14312
rect 3544 14290 3617 14312
rect 2923 14256 3617 14290
rect 2923 14222 2982 14256
rect 3016 14224 3072 14256
rect 3044 14222 3072 14224
rect 3106 14224 3162 14256
rect 3106 14222 3110 14224
rect 2923 14190 3010 14222
rect 3044 14190 3110 14222
rect 3144 14222 3162 14224
rect 3196 14224 3252 14256
rect 3196 14222 3210 14224
rect 3144 14190 3210 14222
rect 3244 14222 3252 14224
rect 3286 14224 3342 14256
rect 3376 14224 3432 14256
rect 3466 14224 3522 14256
rect 3286 14222 3310 14224
rect 3376 14222 3410 14224
rect 3466 14222 3510 14224
rect 3556 14222 3617 14256
rect 3244 14190 3310 14222
rect 3344 14190 3410 14222
rect 3444 14190 3510 14222
rect 3544 14190 3617 14222
rect 2923 14166 3617 14190
rect 2923 14132 2982 14166
rect 3016 14132 3072 14166
rect 3106 14132 3162 14166
rect 3196 14132 3252 14166
rect 3286 14132 3342 14166
rect 3376 14132 3432 14166
rect 3466 14132 3522 14166
rect 3556 14132 3617 14166
rect 2923 14124 3617 14132
rect 2923 14090 3010 14124
rect 3044 14090 3110 14124
rect 3144 14090 3210 14124
rect 3244 14090 3310 14124
rect 3344 14090 3410 14124
rect 3444 14090 3510 14124
rect 3544 14090 3617 14124
rect 2923 14076 3617 14090
rect 2923 14042 2982 14076
rect 3016 14042 3072 14076
rect 3106 14042 3162 14076
rect 3196 14042 3252 14076
rect 3286 14042 3342 14076
rect 3376 14042 3432 14076
rect 3466 14042 3522 14076
rect 3556 14042 3617 14076
rect 2923 14024 3617 14042
rect 2923 13990 3010 14024
rect 3044 13990 3110 14024
rect 3144 13990 3210 14024
rect 3244 13990 3310 14024
rect 3344 13990 3410 14024
rect 3444 13990 3510 14024
rect 3544 13990 3617 14024
rect 2923 13986 3617 13990
rect 2923 13952 2982 13986
rect 3016 13952 3072 13986
rect 3106 13952 3162 13986
rect 3196 13952 3252 13986
rect 3286 13952 3342 13986
rect 3376 13952 3432 13986
rect 3466 13952 3522 13986
rect 3556 13952 3617 13986
rect 2923 13924 3617 13952
rect 2923 13896 3010 13924
rect 3044 13896 3110 13924
rect 2923 13862 2982 13896
rect 3044 13890 3072 13896
rect 3016 13862 3072 13890
rect 3106 13890 3110 13896
rect 3144 13896 3210 13924
rect 3144 13890 3162 13896
rect 3106 13862 3162 13890
rect 3196 13890 3210 13896
rect 3244 13896 3310 13924
rect 3344 13896 3410 13924
rect 3444 13896 3510 13924
rect 3544 13896 3617 13924
rect 3244 13890 3252 13896
rect 3196 13862 3252 13890
rect 3286 13890 3310 13896
rect 3376 13890 3410 13896
rect 3466 13890 3510 13896
rect 3286 13862 3342 13890
rect 3376 13862 3432 13890
rect 3466 13862 3522 13890
rect 3556 13862 3617 13896
rect 2923 13803 3617 13862
rect 3679 14465 3698 14499
rect 3732 14465 3751 14499
rect 3679 14409 3751 14465
rect 3679 14375 3698 14409
rect 3732 14375 3751 14409
rect 3679 14319 3751 14375
rect 3679 14285 3698 14319
rect 3732 14285 3751 14319
rect 3679 14229 3751 14285
rect 3679 14195 3698 14229
rect 3732 14195 3751 14229
rect 3679 14139 3751 14195
rect 3679 14105 3698 14139
rect 3732 14105 3751 14139
rect 3679 14049 3751 14105
rect 3679 14015 3698 14049
rect 3732 14015 3751 14049
rect 3679 13959 3751 14015
rect 3679 13925 3698 13959
rect 3732 13925 3751 13959
rect 3679 13869 3751 13925
rect 3679 13835 3698 13869
rect 3732 13835 3751 13869
rect 2789 13764 2808 13798
rect 2842 13764 2861 13798
rect 2789 13750 2861 13764
rect 3679 13779 3751 13835
rect 3679 13750 3698 13779
rect 2693 13745 3698 13750
rect 3732 13750 3751 13779
rect 3815 14588 4085 14644
rect 5175 14678 5274 14695
rect 5175 14644 5206 14678
rect 5240 14644 5274 14678
rect 3815 14554 3846 14588
rect 3880 14554 4019 14588
rect 4053 14554 4085 14588
rect 3815 14498 4085 14554
rect 3815 14464 3846 14498
rect 3880 14464 4019 14498
rect 4053 14464 4085 14498
rect 3815 14408 4085 14464
rect 3815 14374 3846 14408
rect 3880 14374 4019 14408
rect 4053 14374 4085 14408
rect 3815 14318 4085 14374
rect 3815 14284 3846 14318
rect 3880 14284 4019 14318
rect 4053 14284 4085 14318
rect 3815 14228 4085 14284
rect 3815 14194 3846 14228
rect 3880 14194 4019 14228
rect 4053 14194 4085 14228
rect 3815 14138 4085 14194
rect 3815 14104 3846 14138
rect 3880 14104 4019 14138
rect 4053 14104 4085 14138
rect 3815 14048 4085 14104
rect 3815 14014 3846 14048
rect 3880 14014 4019 14048
rect 4053 14014 4085 14048
rect 3815 13958 4085 14014
rect 3815 13924 3846 13958
rect 3880 13924 4019 13958
rect 4053 13924 4085 13958
rect 3815 13868 4085 13924
rect 3815 13834 3846 13868
rect 3880 13834 4019 13868
rect 4053 13834 4085 13868
rect 3815 13778 4085 13834
rect 3815 13750 3846 13778
rect 3732 13745 3846 13750
rect 2693 13744 3846 13745
rect 3880 13744 4019 13778
rect 4053 13750 4085 13778
rect 4149 14612 5111 14631
rect 4149 14578 4260 14612
rect 4294 14578 4350 14612
rect 4384 14578 4440 14612
rect 4474 14578 4530 14612
rect 4564 14578 4620 14612
rect 4654 14578 4710 14612
rect 4744 14578 4800 14612
rect 4834 14578 4890 14612
rect 4924 14578 4980 14612
rect 5014 14578 5111 14612
rect 4149 14559 5111 14578
rect 4149 14518 4221 14559
rect 4149 14484 4168 14518
rect 4202 14484 4221 14518
rect 5039 14499 5111 14559
rect 4149 14428 4221 14484
rect 4149 14394 4168 14428
rect 4202 14394 4221 14428
rect 4149 14338 4221 14394
rect 4149 14304 4168 14338
rect 4202 14304 4221 14338
rect 4149 14248 4221 14304
rect 4149 14214 4168 14248
rect 4202 14214 4221 14248
rect 4149 14158 4221 14214
rect 4149 14124 4168 14158
rect 4202 14124 4221 14158
rect 4149 14068 4221 14124
rect 4149 14034 4168 14068
rect 4202 14034 4221 14068
rect 4149 13978 4221 14034
rect 4149 13944 4168 13978
rect 4202 13944 4221 13978
rect 4149 13888 4221 13944
rect 4149 13854 4168 13888
rect 4202 13854 4221 13888
rect 4149 13798 4221 13854
rect 4283 14436 4977 14497
rect 4283 14402 4342 14436
rect 4376 14424 4432 14436
rect 4404 14402 4432 14424
rect 4466 14424 4522 14436
rect 4466 14402 4470 14424
rect 4283 14390 4370 14402
rect 4404 14390 4470 14402
rect 4504 14402 4522 14424
rect 4556 14424 4612 14436
rect 4556 14402 4570 14424
rect 4504 14390 4570 14402
rect 4604 14402 4612 14424
rect 4646 14424 4702 14436
rect 4736 14424 4792 14436
rect 4826 14424 4882 14436
rect 4646 14402 4670 14424
rect 4736 14402 4770 14424
rect 4826 14402 4870 14424
rect 4916 14402 4977 14436
rect 4604 14390 4670 14402
rect 4704 14390 4770 14402
rect 4804 14390 4870 14402
rect 4904 14390 4977 14402
rect 4283 14346 4977 14390
rect 4283 14312 4342 14346
rect 4376 14324 4432 14346
rect 4404 14312 4432 14324
rect 4466 14324 4522 14346
rect 4466 14312 4470 14324
rect 4283 14290 4370 14312
rect 4404 14290 4470 14312
rect 4504 14312 4522 14324
rect 4556 14324 4612 14346
rect 4556 14312 4570 14324
rect 4504 14290 4570 14312
rect 4604 14312 4612 14324
rect 4646 14324 4702 14346
rect 4736 14324 4792 14346
rect 4826 14324 4882 14346
rect 4646 14312 4670 14324
rect 4736 14312 4770 14324
rect 4826 14312 4870 14324
rect 4916 14312 4977 14346
rect 4604 14290 4670 14312
rect 4704 14290 4770 14312
rect 4804 14290 4870 14312
rect 4904 14290 4977 14312
rect 4283 14256 4977 14290
rect 4283 14222 4342 14256
rect 4376 14224 4432 14256
rect 4404 14222 4432 14224
rect 4466 14224 4522 14256
rect 4466 14222 4470 14224
rect 4283 14190 4370 14222
rect 4404 14190 4470 14222
rect 4504 14222 4522 14224
rect 4556 14224 4612 14256
rect 4556 14222 4570 14224
rect 4504 14190 4570 14222
rect 4604 14222 4612 14224
rect 4646 14224 4702 14256
rect 4736 14224 4792 14256
rect 4826 14224 4882 14256
rect 4646 14222 4670 14224
rect 4736 14222 4770 14224
rect 4826 14222 4870 14224
rect 4916 14222 4977 14256
rect 4604 14190 4670 14222
rect 4704 14190 4770 14222
rect 4804 14190 4870 14222
rect 4904 14190 4977 14222
rect 4283 14166 4977 14190
rect 4283 14132 4342 14166
rect 4376 14132 4432 14166
rect 4466 14132 4522 14166
rect 4556 14132 4612 14166
rect 4646 14132 4702 14166
rect 4736 14132 4792 14166
rect 4826 14132 4882 14166
rect 4916 14132 4977 14166
rect 4283 14124 4977 14132
rect 4283 14090 4370 14124
rect 4404 14090 4470 14124
rect 4504 14090 4570 14124
rect 4604 14090 4670 14124
rect 4704 14090 4770 14124
rect 4804 14090 4870 14124
rect 4904 14090 4977 14124
rect 4283 14076 4977 14090
rect 4283 14042 4342 14076
rect 4376 14042 4432 14076
rect 4466 14042 4522 14076
rect 4556 14042 4612 14076
rect 4646 14042 4702 14076
rect 4736 14042 4792 14076
rect 4826 14042 4882 14076
rect 4916 14042 4977 14076
rect 4283 14024 4977 14042
rect 4283 13990 4370 14024
rect 4404 13990 4470 14024
rect 4504 13990 4570 14024
rect 4604 13990 4670 14024
rect 4704 13990 4770 14024
rect 4804 13990 4870 14024
rect 4904 13990 4977 14024
rect 4283 13986 4977 13990
rect 4283 13952 4342 13986
rect 4376 13952 4432 13986
rect 4466 13952 4522 13986
rect 4556 13952 4612 13986
rect 4646 13952 4702 13986
rect 4736 13952 4792 13986
rect 4826 13952 4882 13986
rect 4916 13952 4977 13986
rect 4283 13924 4977 13952
rect 4283 13896 4370 13924
rect 4404 13896 4470 13924
rect 4283 13862 4342 13896
rect 4404 13890 4432 13896
rect 4376 13862 4432 13890
rect 4466 13890 4470 13896
rect 4504 13896 4570 13924
rect 4504 13890 4522 13896
rect 4466 13862 4522 13890
rect 4556 13890 4570 13896
rect 4604 13896 4670 13924
rect 4704 13896 4770 13924
rect 4804 13896 4870 13924
rect 4904 13896 4977 13924
rect 4604 13890 4612 13896
rect 4556 13862 4612 13890
rect 4646 13890 4670 13896
rect 4736 13890 4770 13896
rect 4826 13890 4870 13896
rect 4646 13862 4702 13890
rect 4736 13862 4792 13890
rect 4826 13862 4882 13890
rect 4916 13862 4977 13896
rect 4283 13803 4977 13862
rect 5039 14465 5058 14499
rect 5092 14465 5111 14499
rect 5039 14409 5111 14465
rect 5039 14375 5058 14409
rect 5092 14375 5111 14409
rect 5039 14319 5111 14375
rect 5039 14285 5058 14319
rect 5092 14285 5111 14319
rect 5039 14229 5111 14285
rect 5039 14195 5058 14229
rect 5092 14195 5111 14229
rect 5039 14139 5111 14195
rect 5039 14105 5058 14139
rect 5092 14105 5111 14139
rect 5039 14049 5111 14105
rect 5039 14015 5058 14049
rect 5092 14015 5111 14049
rect 5039 13959 5111 14015
rect 5039 13925 5058 13959
rect 5092 13925 5111 13959
rect 5039 13869 5111 13925
rect 5039 13835 5058 13869
rect 5092 13835 5111 13869
rect 4149 13764 4168 13798
rect 4202 13764 4221 13798
rect 4149 13750 4221 13764
rect 5039 13779 5111 13835
rect 5039 13750 5058 13779
rect 4053 13745 5058 13750
rect 5092 13750 5111 13779
rect 5175 14588 5274 14644
rect 5175 14554 5206 14588
rect 5240 14554 5274 14588
rect 5175 14498 5274 14554
rect 5175 14464 5206 14498
rect 5240 14464 5274 14498
rect 5175 14408 5274 14464
rect 5175 14374 5206 14408
rect 5240 14374 5274 14408
rect 5175 14318 5274 14374
rect 5175 14284 5206 14318
rect 5240 14284 5274 14318
rect 5175 14228 5274 14284
rect 5175 14194 5206 14228
rect 5240 14194 5274 14228
rect 5175 14138 5274 14194
rect 5175 14104 5206 14138
rect 5240 14104 5274 14138
rect 5175 14048 5274 14104
rect 5175 14014 5206 14048
rect 5240 14014 5274 14048
rect 5440 14548 5510 14568
rect 5440 14498 5450 14548
rect 5500 14498 5510 14548
rect 5440 14478 5510 14498
rect 5630 14408 5680 14478
rect 5800 14398 5870 14418
rect 5800 14348 5810 14398
rect 5860 14348 5870 14398
rect 5800 14328 5870 14348
rect 5175 13958 5274 14014
rect 5175 13924 5206 13958
rect 5240 13924 5274 13958
rect 5175 13868 5274 13924
rect 6460 14398 6530 14418
rect 6460 14348 6470 14398
rect 6520 14348 6530 14398
rect 6460 14328 6530 14348
rect 5175 13834 5206 13868
rect 5240 13834 5274 13868
rect 5175 13778 5274 13834
rect 5175 13750 5206 13778
rect 5092 13745 5206 13750
rect 4053 13744 5206 13745
rect 5240 13750 5274 13778
rect 5240 13744 5280 13750
rect 1260 13722 5280 13744
rect 1260 13688 1506 13722
rect 1540 13688 1596 13722
rect 1630 13688 1686 13722
rect 1720 13688 1776 13722
rect 1810 13688 1866 13722
rect 1900 13688 1956 13722
rect 1990 13688 2046 13722
rect 2080 13688 2136 13722
rect 2170 13688 2226 13722
rect 2260 13688 2866 13722
rect 2900 13688 2956 13722
rect 2990 13688 3046 13722
rect 3080 13688 3136 13722
rect 3170 13688 3226 13722
rect 3260 13688 3316 13722
rect 3350 13688 3406 13722
rect 3440 13688 3496 13722
rect 3530 13688 3586 13722
rect 3620 13688 4226 13722
rect 4260 13688 4316 13722
rect 4350 13688 4406 13722
rect 4440 13688 4496 13722
rect 4530 13688 4586 13722
rect 4620 13688 4676 13722
rect 4710 13688 4766 13722
rect 4800 13688 4856 13722
rect 4890 13688 4946 13722
rect 4980 13688 5280 13722
rect 1260 13654 1299 13688
rect 1333 13654 2486 13688
rect 2520 13654 2659 13688
rect 2693 13654 3846 13688
rect 3880 13654 4019 13688
rect 4053 13654 5206 13688
rect 5240 13654 5280 13688
rect 1260 13598 5280 13654
rect 1260 13564 1299 13598
rect 1333 13575 2486 13598
rect 1333 13564 1400 13575
rect 1260 13541 1400 13564
rect 1434 13541 1490 13575
rect 1524 13541 1580 13575
rect 1614 13541 1670 13575
rect 1704 13541 1760 13575
rect 1794 13541 1850 13575
rect 1884 13541 1940 13575
rect 1974 13541 2030 13575
rect 2064 13541 2120 13575
rect 2154 13541 2210 13575
rect 2244 13541 2300 13575
rect 2334 13541 2390 13575
rect 2424 13564 2486 13575
rect 2520 13564 2659 13598
rect 2693 13575 3846 13598
rect 2693 13564 2760 13575
rect 2424 13541 2760 13564
rect 2794 13541 2850 13575
rect 2884 13541 2940 13575
rect 2974 13541 3030 13575
rect 3064 13541 3120 13575
rect 3154 13541 3210 13575
rect 3244 13541 3300 13575
rect 3334 13541 3390 13575
rect 3424 13541 3480 13575
rect 3514 13541 3570 13575
rect 3604 13541 3660 13575
rect 3694 13541 3750 13575
rect 3784 13564 3846 13575
rect 3880 13564 4019 13598
rect 4053 13575 5206 13598
rect 4053 13564 4120 13575
rect 3784 13541 4120 13564
rect 4154 13541 4210 13575
rect 4244 13541 4300 13575
rect 4334 13541 4390 13575
rect 4424 13541 4480 13575
rect 4514 13541 4570 13575
rect 4604 13541 4660 13575
rect 4694 13541 4750 13575
rect 4784 13541 4840 13575
rect 4874 13541 4930 13575
rect 4964 13541 5020 13575
rect 5054 13541 5110 13575
rect 5144 13564 5206 13575
rect 5240 13564 5280 13598
rect 5144 13541 5280 13564
rect 1260 13500 5280 13541
rect 2550 13434 2630 13500
rect 3910 13434 3990 13500
rect 1266 13402 5274 13434
rect 1266 13368 1400 13402
rect 1434 13368 1490 13402
rect 1524 13368 1580 13402
rect 1614 13368 1670 13402
rect 1704 13368 1760 13402
rect 1794 13368 1850 13402
rect 1884 13368 1940 13402
rect 1974 13368 2030 13402
rect 2064 13368 2120 13402
rect 2154 13368 2210 13402
rect 2244 13368 2300 13402
rect 2334 13368 2390 13402
rect 2424 13368 2760 13402
rect 2794 13368 2850 13402
rect 2884 13368 2940 13402
rect 2974 13368 3030 13402
rect 3064 13368 3120 13402
rect 3154 13368 3210 13402
rect 3244 13368 3300 13402
rect 3334 13368 3390 13402
rect 3424 13368 3480 13402
rect 3514 13368 3570 13402
rect 3604 13368 3660 13402
rect 3694 13368 3750 13402
rect 3784 13368 4120 13402
rect 4154 13368 4210 13402
rect 4244 13368 4300 13402
rect 4334 13368 4390 13402
rect 4424 13368 4480 13402
rect 4514 13368 4570 13402
rect 4604 13368 4660 13402
rect 4694 13368 4750 13402
rect 4784 13368 4840 13402
rect 4874 13368 4930 13402
rect 4964 13368 5020 13402
rect 5054 13368 5110 13402
rect 5144 13368 5274 13402
rect 1266 13335 5274 13368
rect 1266 13318 1365 13335
rect 1266 13284 1299 13318
rect 1333 13284 1365 13318
rect 120 12840 190 12862
rect 120 12790 130 12840
rect 180 12790 190 12840
rect 120 12770 190 12790
rect 430 12810 480 12880
rect 1266 13228 1365 13284
rect 2455 13318 2725 13335
rect 2455 13284 2486 13318
rect 2520 13284 2659 13318
rect 2693 13284 2725 13318
rect 1266 13194 1299 13228
rect 1333 13194 1365 13228
rect 1266 13138 1365 13194
rect 1266 13104 1299 13138
rect 1333 13104 1365 13138
rect 1266 13048 1365 13104
rect 1266 13014 1299 13048
rect 1333 13014 1365 13048
rect 1266 12958 1365 13014
rect 1266 12924 1299 12958
rect 1333 12924 1365 12958
rect 240 12790 310 12810
rect 240 12740 250 12790
rect 300 12740 310 12790
rect 240 12720 310 12740
rect 860 12430 910 12500
rect 1266 12868 1365 12924
rect 1266 12834 1299 12868
rect 1333 12834 1365 12868
rect 1266 12778 1365 12834
rect 1266 12744 1299 12778
rect 1333 12744 1365 12778
rect 1266 12688 1365 12744
rect 1266 12654 1299 12688
rect 1333 12654 1365 12688
rect 1266 12598 1365 12654
rect 1266 12564 1299 12598
rect 1333 12564 1365 12598
rect 1266 12508 1365 12564
rect 1266 12474 1299 12508
rect 1333 12474 1365 12508
rect 670 12410 740 12430
rect 670 12360 680 12410
rect 730 12360 740 12410
rect 1266 12418 1365 12474
rect 1266 12390 1299 12418
rect 670 12340 740 12360
rect 1260 12384 1299 12390
rect 1333 12390 1365 12418
rect 1429 13252 2391 13271
rect 1429 13218 1540 13252
rect 1574 13218 1630 13252
rect 1664 13218 1720 13252
rect 1754 13218 1810 13252
rect 1844 13218 1900 13252
rect 1934 13218 1990 13252
rect 2024 13218 2080 13252
rect 2114 13218 2170 13252
rect 2204 13218 2260 13252
rect 2294 13218 2391 13252
rect 1429 13199 2391 13218
rect 1429 13158 1501 13199
rect 1429 13124 1448 13158
rect 1482 13124 1501 13158
rect 2319 13139 2391 13199
rect 1429 13068 1501 13124
rect 1429 13034 1448 13068
rect 1482 13034 1501 13068
rect 1429 12978 1501 13034
rect 1429 12944 1448 12978
rect 1482 12944 1501 12978
rect 1429 12888 1501 12944
rect 1429 12854 1448 12888
rect 1482 12854 1501 12888
rect 1429 12798 1501 12854
rect 1429 12764 1448 12798
rect 1482 12764 1501 12798
rect 1429 12708 1501 12764
rect 1429 12674 1448 12708
rect 1482 12674 1501 12708
rect 1429 12618 1501 12674
rect 1429 12584 1448 12618
rect 1482 12584 1501 12618
rect 1429 12528 1501 12584
rect 1429 12494 1448 12528
rect 1482 12494 1501 12528
rect 1429 12438 1501 12494
rect 1563 13076 2257 13137
rect 1563 13042 1622 13076
rect 1656 13064 1712 13076
rect 1684 13042 1712 13064
rect 1746 13064 1802 13076
rect 1746 13042 1750 13064
rect 1563 13030 1650 13042
rect 1684 13030 1750 13042
rect 1784 13042 1802 13064
rect 1836 13064 1892 13076
rect 1836 13042 1850 13064
rect 1784 13030 1850 13042
rect 1884 13042 1892 13064
rect 1926 13064 1982 13076
rect 2016 13064 2072 13076
rect 2106 13064 2162 13076
rect 1926 13042 1950 13064
rect 2016 13042 2050 13064
rect 2106 13042 2150 13064
rect 2196 13042 2257 13076
rect 1884 13030 1950 13042
rect 1984 13030 2050 13042
rect 2084 13030 2150 13042
rect 2184 13030 2257 13042
rect 1563 12986 2257 13030
rect 1563 12952 1622 12986
rect 1656 12964 1712 12986
rect 1684 12952 1712 12964
rect 1746 12964 1802 12986
rect 1746 12952 1750 12964
rect 1563 12930 1650 12952
rect 1684 12930 1750 12952
rect 1784 12952 1802 12964
rect 1836 12964 1892 12986
rect 1836 12952 1850 12964
rect 1784 12930 1850 12952
rect 1884 12952 1892 12964
rect 1926 12964 1982 12986
rect 2016 12964 2072 12986
rect 2106 12964 2162 12986
rect 1926 12952 1950 12964
rect 2016 12952 2050 12964
rect 2106 12952 2150 12964
rect 2196 12952 2257 12986
rect 1884 12930 1950 12952
rect 1984 12930 2050 12952
rect 2084 12930 2150 12952
rect 2184 12930 2257 12952
rect 1563 12896 2257 12930
rect 1563 12862 1622 12896
rect 1656 12864 1712 12896
rect 1684 12862 1712 12864
rect 1746 12864 1802 12896
rect 1746 12862 1750 12864
rect 1563 12830 1650 12862
rect 1684 12830 1750 12862
rect 1784 12862 1802 12864
rect 1836 12864 1892 12896
rect 1836 12862 1850 12864
rect 1784 12830 1850 12862
rect 1884 12862 1892 12864
rect 1926 12864 1982 12896
rect 2016 12864 2072 12896
rect 2106 12864 2162 12896
rect 1926 12862 1950 12864
rect 2016 12862 2050 12864
rect 2106 12862 2150 12864
rect 2196 12862 2257 12896
rect 1884 12830 1950 12862
rect 1984 12830 2050 12862
rect 2084 12830 2150 12862
rect 2184 12830 2257 12862
rect 1563 12806 2257 12830
rect 1563 12772 1622 12806
rect 1656 12772 1712 12806
rect 1746 12772 1802 12806
rect 1836 12772 1892 12806
rect 1926 12772 1982 12806
rect 2016 12772 2072 12806
rect 2106 12772 2162 12806
rect 2196 12772 2257 12806
rect 1563 12764 2257 12772
rect 1563 12730 1650 12764
rect 1684 12730 1750 12764
rect 1784 12730 1850 12764
rect 1884 12730 1950 12764
rect 1984 12730 2050 12764
rect 2084 12730 2150 12764
rect 2184 12730 2257 12764
rect 1563 12716 2257 12730
rect 1563 12682 1622 12716
rect 1656 12682 1712 12716
rect 1746 12682 1802 12716
rect 1836 12682 1892 12716
rect 1926 12682 1982 12716
rect 2016 12682 2072 12716
rect 2106 12682 2162 12716
rect 2196 12682 2257 12716
rect 1563 12664 2257 12682
rect 1563 12630 1650 12664
rect 1684 12630 1750 12664
rect 1784 12630 1850 12664
rect 1884 12630 1950 12664
rect 1984 12630 2050 12664
rect 2084 12630 2150 12664
rect 2184 12630 2257 12664
rect 1563 12626 2257 12630
rect 1563 12592 1622 12626
rect 1656 12592 1712 12626
rect 1746 12592 1802 12626
rect 1836 12592 1892 12626
rect 1926 12592 1982 12626
rect 2016 12592 2072 12626
rect 2106 12592 2162 12626
rect 2196 12592 2257 12626
rect 1563 12564 2257 12592
rect 1563 12536 1650 12564
rect 1684 12536 1750 12564
rect 1563 12502 1622 12536
rect 1684 12530 1712 12536
rect 1656 12502 1712 12530
rect 1746 12530 1750 12536
rect 1784 12536 1850 12564
rect 1784 12530 1802 12536
rect 1746 12502 1802 12530
rect 1836 12530 1850 12536
rect 1884 12536 1950 12564
rect 1984 12536 2050 12564
rect 2084 12536 2150 12564
rect 2184 12536 2257 12564
rect 1884 12530 1892 12536
rect 1836 12502 1892 12530
rect 1926 12530 1950 12536
rect 2016 12530 2050 12536
rect 2106 12530 2150 12536
rect 1926 12502 1982 12530
rect 2016 12502 2072 12530
rect 2106 12502 2162 12530
rect 2196 12502 2257 12536
rect 1563 12443 2257 12502
rect 2319 13105 2338 13139
rect 2372 13105 2391 13139
rect 2319 13049 2391 13105
rect 2319 13015 2338 13049
rect 2372 13015 2391 13049
rect 2319 12959 2391 13015
rect 2319 12925 2338 12959
rect 2372 12925 2391 12959
rect 2319 12869 2391 12925
rect 2319 12835 2338 12869
rect 2372 12835 2391 12869
rect 2319 12779 2391 12835
rect 2319 12745 2338 12779
rect 2372 12745 2391 12779
rect 2319 12689 2391 12745
rect 2319 12655 2338 12689
rect 2372 12655 2391 12689
rect 2319 12599 2391 12655
rect 2319 12565 2338 12599
rect 2372 12565 2391 12599
rect 2319 12509 2391 12565
rect 2319 12475 2338 12509
rect 2372 12475 2391 12509
rect 1429 12404 1448 12438
rect 1482 12404 1501 12438
rect 1429 12390 1501 12404
rect 2319 12419 2391 12475
rect 2319 12390 2338 12419
rect 1333 12385 2338 12390
rect 2372 12390 2391 12419
rect 2455 13228 2725 13284
rect 3815 13318 4085 13335
rect 3815 13284 3846 13318
rect 3880 13284 4019 13318
rect 4053 13284 4085 13318
rect 2455 13194 2486 13228
rect 2520 13194 2659 13228
rect 2693 13194 2725 13228
rect 2455 13138 2725 13194
rect 2455 13104 2486 13138
rect 2520 13104 2659 13138
rect 2693 13104 2725 13138
rect 2455 13048 2725 13104
rect 2455 13014 2486 13048
rect 2520 13014 2659 13048
rect 2693 13014 2725 13048
rect 2455 12958 2725 13014
rect 2455 12924 2486 12958
rect 2520 12924 2659 12958
rect 2693 12924 2725 12958
rect 2455 12868 2725 12924
rect 2455 12834 2486 12868
rect 2520 12834 2659 12868
rect 2693 12834 2725 12868
rect 2455 12778 2725 12834
rect 2455 12744 2486 12778
rect 2520 12744 2659 12778
rect 2693 12744 2725 12778
rect 2455 12688 2725 12744
rect 2455 12654 2486 12688
rect 2520 12654 2659 12688
rect 2693 12654 2725 12688
rect 2455 12598 2725 12654
rect 2455 12564 2486 12598
rect 2520 12564 2659 12598
rect 2693 12564 2725 12598
rect 2455 12508 2725 12564
rect 2455 12474 2486 12508
rect 2520 12474 2659 12508
rect 2693 12474 2725 12508
rect 2455 12418 2725 12474
rect 2455 12390 2486 12418
rect 2372 12385 2486 12390
rect 1333 12384 2486 12385
rect 2520 12384 2659 12418
rect 2693 12390 2725 12418
rect 2789 13252 3751 13271
rect 2789 13218 2900 13252
rect 2934 13218 2990 13252
rect 3024 13218 3080 13252
rect 3114 13218 3170 13252
rect 3204 13218 3260 13252
rect 3294 13218 3350 13252
rect 3384 13218 3440 13252
rect 3474 13218 3530 13252
rect 3564 13218 3620 13252
rect 3654 13218 3751 13252
rect 2789 13199 3751 13218
rect 2789 13158 2861 13199
rect 2789 13124 2808 13158
rect 2842 13124 2861 13158
rect 3679 13139 3751 13199
rect 2789 13068 2861 13124
rect 2789 13034 2808 13068
rect 2842 13034 2861 13068
rect 2789 12978 2861 13034
rect 2789 12944 2808 12978
rect 2842 12944 2861 12978
rect 2789 12888 2861 12944
rect 2789 12854 2808 12888
rect 2842 12854 2861 12888
rect 2789 12798 2861 12854
rect 2789 12764 2808 12798
rect 2842 12764 2861 12798
rect 2789 12708 2861 12764
rect 2789 12674 2808 12708
rect 2842 12674 2861 12708
rect 2789 12618 2861 12674
rect 2789 12584 2808 12618
rect 2842 12584 2861 12618
rect 2789 12528 2861 12584
rect 2789 12494 2808 12528
rect 2842 12494 2861 12528
rect 2789 12438 2861 12494
rect 2923 13076 3617 13137
rect 2923 13042 2982 13076
rect 3016 13064 3072 13076
rect 3044 13042 3072 13064
rect 3106 13064 3162 13076
rect 3106 13042 3110 13064
rect 2923 13030 3010 13042
rect 3044 13030 3110 13042
rect 3144 13042 3162 13064
rect 3196 13064 3252 13076
rect 3196 13042 3210 13064
rect 3144 13030 3210 13042
rect 3244 13042 3252 13064
rect 3286 13064 3342 13076
rect 3376 13064 3432 13076
rect 3466 13064 3522 13076
rect 3286 13042 3310 13064
rect 3376 13042 3410 13064
rect 3466 13042 3510 13064
rect 3556 13042 3617 13076
rect 3244 13030 3310 13042
rect 3344 13030 3410 13042
rect 3444 13030 3510 13042
rect 3544 13030 3617 13042
rect 2923 12986 3617 13030
rect 2923 12952 2982 12986
rect 3016 12964 3072 12986
rect 3044 12952 3072 12964
rect 3106 12964 3162 12986
rect 3106 12952 3110 12964
rect 2923 12930 3010 12952
rect 3044 12930 3110 12952
rect 3144 12952 3162 12964
rect 3196 12964 3252 12986
rect 3196 12952 3210 12964
rect 3144 12930 3210 12952
rect 3244 12952 3252 12964
rect 3286 12964 3342 12986
rect 3376 12964 3432 12986
rect 3466 12964 3522 12986
rect 3286 12952 3310 12964
rect 3376 12952 3410 12964
rect 3466 12952 3510 12964
rect 3556 12952 3617 12986
rect 3244 12930 3310 12952
rect 3344 12930 3410 12952
rect 3444 12930 3510 12952
rect 3544 12930 3617 12952
rect 2923 12896 3617 12930
rect 2923 12862 2982 12896
rect 3016 12864 3072 12896
rect 3044 12862 3072 12864
rect 3106 12864 3162 12896
rect 3106 12862 3110 12864
rect 2923 12830 3010 12862
rect 3044 12830 3110 12862
rect 3144 12862 3162 12864
rect 3196 12864 3252 12896
rect 3196 12862 3210 12864
rect 3144 12830 3210 12862
rect 3244 12862 3252 12864
rect 3286 12864 3342 12896
rect 3376 12864 3432 12896
rect 3466 12864 3522 12896
rect 3286 12862 3310 12864
rect 3376 12862 3410 12864
rect 3466 12862 3510 12864
rect 3556 12862 3617 12896
rect 3244 12830 3310 12862
rect 3344 12830 3410 12862
rect 3444 12830 3510 12862
rect 3544 12830 3617 12862
rect 2923 12806 3617 12830
rect 2923 12772 2982 12806
rect 3016 12772 3072 12806
rect 3106 12772 3162 12806
rect 3196 12772 3252 12806
rect 3286 12772 3342 12806
rect 3376 12772 3432 12806
rect 3466 12772 3522 12806
rect 3556 12772 3617 12806
rect 2923 12764 3617 12772
rect 2923 12730 3010 12764
rect 3044 12730 3110 12764
rect 3144 12730 3210 12764
rect 3244 12730 3310 12764
rect 3344 12730 3410 12764
rect 3444 12730 3510 12764
rect 3544 12730 3617 12764
rect 2923 12716 3617 12730
rect 2923 12682 2982 12716
rect 3016 12682 3072 12716
rect 3106 12682 3162 12716
rect 3196 12682 3252 12716
rect 3286 12682 3342 12716
rect 3376 12682 3432 12716
rect 3466 12682 3522 12716
rect 3556 12682 3617 12716
rect 2923 12664 3617 12682
rect 2923 12630 3010 12664
rect 3044 12630 3110 12664
rect 3144 12630 3210 12664
rect 3244 12630 3310 12664
rect 3344 12630 3410 12664
rect 3444 12630 3510 12664
rect 3544 12630 3617 12664
rect 2923 12626 3617 12630
rect 2923 12592 2982 12626
rect 3016 12592 3072 12626
rect 3106 12592 3162 12626
rect 3196 12592 3252 12626
rect 3286 12592 3342 12626
rect 3376 12592 3432 12626
rect 3466 12592 3522 12626
rect 3556 12592 3617 12626
rect 2923 12564 3617 12592
rect 2923 12536 3010 12564
rect 3044 12536 3110 12564
rect 2923 12502 2982 12536
rect 3044 12530 3072 12536
rect 3016 12502 3072 12530
rect 3106 12530 3110 12536
rect 3144 12536 3210 12564
rect 3144 12530 3162 12536
rect 3106 12502 3162 12530
rect 3196 12530 3210 12536
rect 3244 12536 3310 12564
rect 3344 12536 3410 12564
rect 3444 12536 3510 12564
rect 3544 12536 3617 12564
rect 3244 12530 3252 12536
rect 3196 12502 3252 12530
rect 3286 12530 3310 12536
rect 3376 12530 3410 12536
rect 3466 12530 3510 12536
rect 3286 12502 3342 12530
rect 3376 12502 3432 12530
rect 3466 12502 3522 12530
rect 3556 12502 3617 12536
rect 2923 12443 3617 12502
rect 3679 13105 3698 13139
rect 3732 13105 3751 13139
rect 3679 13049 3751 13105
rect 3679 13015 3698 13049
rect 3732 13015 3751 13049
rect 3679 12959 3751 13015
rect 3679 12925 3698 12959
rect 3732 12925 3751 12959
rect 3679 12869 3751 12925
rect 3679 12835 3698 12869
rect 3732 12835 3751 12869
rect 3679 12779 3751 12835
rect 3679 12745 3698 12779
rect 3732 12745 3751 12779
rect 3679 12689 3751 12745
rect 3679 12655 3698 12689
rect 3732 12655 3751 12689
rect 3679 12599 3751 12655
rect 3679 12565 3698 12599
rect 3732 12565 3751 12599
rect 3679 12509 3751 12565
rect 3679 12475 3698 12509
rect 3732 12475 3751 12509
rect 2789 12404 2808 12438
rect 2842 12404 2861 12438
rect 2789 12390 2861 12404
rect 3679 12419 3751 12475
rect 3679 12390 3698 12419
rect 2693 12385 3698 12390
rect 3732 12390 3751 12419
rect 3815 13228 4085 13284
rect 5175 13318 5274 13335
rect 5175 13284 5206 13318
rect 5240 13284 5274 13318
rect 3815 13194 3846 13228
rect 3880 13194 4019 13228
rect 4053 13194 4085 13228
rect 3815 13138 4085 13194
rect 3815 13104 3846 13138
rect 3880 13104 4019 13138
rect 4053 13104 4085 13138
rect 3815 13048 4085 13104
rect 3815 13014 3846 13048
rect 3880 13014 4019 13048
rect 4053 13014 4085 13048
rect 3815 12958 4085 13014
rect 3815 12924 3846 12958
rect 3880 12924 4019 12958
rect 4053 12924 4085 12958
rect 3815 12868 4085 12924
rect 3815 12834 3846 12868
rect 3880 12834 4019 12868
rect 4053 12834 4085 12868
rect 3815 12778 4085 12834
rect 3815 12744 3846 12778
rect 3880 12744 4019 12778
rect 4053 12744 4085 12778
rect 3815 12688 4085 12744
rect 3815 12654 3846 12688
rect 3880 12654 4019 12688
rect 4053 12654 4085 12688
rect 3815 12598 4085 12654
rect 3815 12564 3846 12598
rect 3880 12564 4019 12598
rect 4053 12564 4085 12598
rect 3815 12508 4085 12564
rect 3815 12474 3846 12508
rect 3880 12474 4019 12508
rect 4053 12474 4085 12508
rect 3815 12418 4085 12474
rect 3815 12390 3846 12418
rect 3732 12385 3846 12390
rect 2693 12384 3846 12385
rect 3880 12384 4019 12418
rect 4053 12390 4085 12418
rect 4149 13252 5111 13271
rect 4149 13218 4260 13252
rect 4294 13218 4350 13252
rect 4384 13218 4440 13252
rect 4474 13218 4530 13252
rect 4564 13218 4620 13252
rect 4654 13218 4710 13252
rect 4744 13218 4800 13252
rect 4834 13218 4890 13252
rect 4924 13218 4980 13252
rect 5014 13218 5111 13252
rect 4149 13199 5111 13218
rect 4149 13158 4221 13199
rect 4149 13124 4168 13158
rect 4202 13124 4221 13158
rect 5039 13139 5111 13199
rect 4149 13068 4221 13124
rect 4149 13034 4168 13068
rect 4202 13034 4221 13068
rect 4149 12978 4221 13034
rect 4149 12944 4168 12978
rect 4202 12944 4221 12978
rect 4149 12888 4221 12944
rect 4149 12854 4168 12888
rect 4202 12854 4221 12888
rect 4149 12798 4221 12854
rect 4149 12764 4168 12798
rect 4202 12764 4221 12798
rect 4149 12708 4221 12764
rect 4149 12674 4168 12708
rect 4202 12674 4221 12708
rect 4149 12618 4221 12674
rect 4149 12584 4168 12618
rect 4202 12584 4221 12618
rect 4149 12528 4221 12584
rect 4149 12494 4168 12528
rect 4202 12494 4221 12528
rect 4149 12438 4221 12494
rect 4283 13076 4977 13137
rect 4283 13042 4342 13076
rect 4376 13064 4432 13076
rect 4404 13042 4432 13064
rect 4466 13064 4522 13076
rect 4466 13042 4470 13064
rect 4283 13030 4370 13042
rect 4404 13030 4470 13042
rect 4504 13042 4522 13064
rect 4556 13064 4612 13076
rect 4556 13042 4570 13064
rect 4504 13030 4570 13042
rect 4604 13042 4612 13064
rect 4646 13064 4702 13076
rect 4736 13064 4792 13076
rect 4826 13064 4882 13076
rect 4646 13042 4670 13064
rect 4736 13042 4770 13064
rect 4826 13042 4870 13064
rect 4916 13042 4977 13076
rect 4604 13030 4670 13042
rect 4704 13030 4770 13042
rect 4804 13030 4870 13042
rect 4904 13030 4977 13042
rect 4283 12986 4977 13030
rect 4283 12952 4342 12986
rect 4376 12964 4432 12986
rect 4404 12952 4432 12964
rect 4466 12964 4522 12986
rect 4466 12952 4470 12964
rect 4283 12930 4370 12952
rect 4404 12930 4470 12952
rect 4504 12952 4522 12964
rect 4556 12964 4612 12986
rect 4556 12952 4570 12964
rect 4504 12930 4570 12952
rect 4604 12952 4612 12964
rect 4646 12964 4702 12986
rect 4736 12964 4792 12986
rect 4826 12964 4882 12986
rect 4646 12952 4670 12964
rect 4736 12952 4770 12964
rect 4826 12952 4870 12964
rect 4916 12952 4977 12986
rect 4604 12930 4670 12952
rect 4704 12930 4770 12952
rect 4804 12930 4870 12952
rect 4904 12930 4977 12952
rect 4283 12896 4977 12930
rect 4283 12862 4342 12896
rect 4376 12864 4432 12896
rect 4404 12862 4432 12864
rect 4466 12864 4522 12896
rect 4466 12862 4470 12864
rect 4283 12830 4370 12862
rect 4404 12830 4470 12862
rect 4504 12862 4522 12864
rect 4556 12864 4612 12896
rect 4556 12862 4570 12864
rect 4504 12830 4570 12862
rect 4604 12862 4612 12864
rect 4646 12864 4702 12896
rect 4736 12864 4792 12896
rect 4826 12864 4882 12896
rect 4646 12862 4670 12864
rect 4736 12862 4770 12864
rect 4826 12862 4870 12864
rect 4916 12862 4977 12896
rect 4604 12830 4670 12862
rect 4704 12830 4770 12862
rect 4804 12830 4870 12862
rect 4904 12830 4977 12862
rect 4283 12806 4977 12830
rect 4283 12772 4342 12806
rect 4376 12772 4432 12806
rect 4466 12772 4522 12806
rect 4556 12772 4612 12806
rect 4646 12772 4702 12806
rect 4736 12772 4792 12806
rect 4826 12772 4882 12806
rect 4916 12772 4977 12806
rect 4283 12764 4977 12772
rect 4283 12730 4370 12764
rect 4404 12730 4470 12764
rect 4504 12730 4570 12764
rect 4604 12730 4670 12764
rect 4704 12730 4770 12764
rect 4804 12730 4870 12764
rect 4904 12730 4977 12764
rect 4283 12716 4977 12730
rect 4283 12682 4342 12716
rect 4376 12682 4432 12716
rect 4466 12682 4522 12716
rect 4556 12682 4612 12716
rect 4646 12682 4702 12716
rect 4736 12682 4792 12716
rect 4826 12682 4882 12716
rect 4916 12682 4977 12716
rect 4283 12664 4977 12682
rect 4283 12630 4370 12664
rect 4404 12630 4470 12664
rect 4504 12630 4570 12664
rect 4604 12630 4670 12664
rect 4704 12630 4770 12664
rect 4804 12630 4870 12664
rect 4904 12630 4977 12664
rect 4283 12626 4977 12630
rect 4283 12592 4342 12626
rect 4376 12592 4432 12626
rect 4466 12592 4522 12626
rect 4556 12592 4612 12626
rect 4646 12592 4702 12626
rect 4736 12592 4792 12626
rect 4826 12592 4882 12626
rect 4916 12592 4977 12626
rect 4283 12564 4977 12592
rect 4283 12536 4370 12564
rect 4404 12536 4470 12564
rect 4283 12502 4342 12536
rect 4404 12530 4432 12536
rect 4376 12502 4432 12530
rect 4466 12530 4470 12536
rect 4504 12536 4570 12564
rect 4504 12530 4522 12536
rect 4466 12502 4522 12530
rect 4556 12530 4570 12536
rect 4604 12536 4670 12564
rect 4704 12536 4770 12564
rect 4804 12536 4870 12564
rect 4904 12536 4977 12564
rect 4604 12530 4612 12536
rect 4556 12502 4612 12530
rect 4646 12530 4670 12536
rect 4736 12530 4770 12536
rect 4826 12530 4870 12536
rect 4646 12502 4702 12530
rect 4736 12502 4792 12530
rect 4826 12502 4882 12530
rect 4916 12502 4977 12536
rect 4283 12443 4977 12502
rect 5039 13105 5058 13139
rect 5092 13105 5111 13139
rect 5039 13049 5111 13105
rect 5039 13015 5058 13049
rect 5092 13015 5111 13049
rect 5039 12959 5111 13015
rect 5039 12925 5058 12959
rect 5092 12925 5111 12959
rect 5039 12869 5111 12925
rect 5039 12835 5058 12869
rect 5092 12835 5111 12869
rect 5039 12779 5111 12835
rect 5039 12745 5058 12779
rect 5092 12745 5111 12779
rect 5039 12689 5111 12745
rect 5039 12655 5058 12689
rect 5092 12655 5111 12689
rect 5039 12599 5111 12655
rect 5039 12565 5058 12599
rect 5092 12565 5111 12599
rect 5039 12509 5111 12565
rect 5039 12475 5058 12509
rect 5092 12475 5111 12509
rect 4149 12404 4168 12438
rect 4202 12404 4221 12438
rect 4149 12390 4221 12404
rect 5039 12419 5111 12475
rect 5039 12390 5058 12419
rect 4053 12385 5058 12390
rect 5092 12390 5111 12419
rect 5175 13228 5274 13284
rect 5175 13194 5206 13228
rect 5240 13194 5274 13228
rect 5175 13138 5274 13194
rect 5800 13260 5870 13280
rect 5800 13210 5810 13260
rect 5860 13210 5870 13260
rect 5800 13190 5870 13210
rect 5175 13104 5206 13138
rect 5240 13104 5274 13138
rect 5175 13048 5274 13104
rect 5175 13014 5206 13048
rect 5240 13014 5274 13048
rect 5175 12958 5274 13014
rect 6460 13052 6530 13072
rect 6460 13002 6470 13052
rect 6520 13002 6530 13052
rect 6460 12980 6530 13002
rect 5175 12924 5206 12958
rect 5240 12924 5274 12958
rect 5175 12868 5274 12924
rect 5175 12834 5206 12868
rect 5240 12834 5274 12868
rect 5175 12778 5274 12834
rect 5175 12744 5206 12778
rect 5240 12744 5274 12778
rect 5175 12688 5274 12744
rect 5175 12654 5206 12688
rect 5240 12654 5274 12688
rect 5175 12598 5274 12654
rect 5175 12564 5206 12598
rect 5240 12564 5274 12598
rect 5175 12508 5274 12564
rect 5175 12474 5206 12508
rect 5240 12474 5274 12508
rect 5175 12418 5274 12474
rect 5510 12430 5560 12500
rect 5175 12390 5206 12418
rect 5092 12385 5206 12390
rect 4053 12384 5206 12385
rect 5240 12390 5274 12418
rect 5680 12410 5750 12430
rect 5240 12384 5280 12390
rect 1260 12362 5280 12384
rect 1260 12328 1506 12362
rect 1540 12328 1596 12362
rect 1630 12328 1686 12362
rect 1720 12328 1776 12362
rect 1810 12328 1866 12362
rect 1900 12328 1956 12362
rect 1990 12328 2046 12362
rect 2080 12328 2136 12362
rect 2170 12328 2226 12362
rect 2260 12328 2866 12362
rect 2900 12328 2956 12362
rect 2990 12328 3046 12362
rect 3080 12328 3136 12362
rect 3170 12328 3226 12362
rect 3260 12328 3316 12362
rect 3350 12328 3406 12362
rect 3440 12328 3496 12362
rect 3530 12328 3586 12362
rect 3620 12328 4226 12362
rect 4260 12328 4316 12362
rect 4350 12328 4406 12362
rect 4440 12328 4496 12362
rect 4530 12328 4586 12362
rect 4620 12328 4676 12362
rect 4710 12328 4766 12362
rect 4800 12328 4856 12362
rect 4890 12328 4946 12362
rect 4980 12328 5280 12362
rect 5680 12360 5690 12410
rect 5740 12360 5750 12410
rect 5680 12340 5750 12360
rect 1260 12294 1299 12328
rect 1333 12294 2486 12328
rect 2520 12294 2659 12328
rect 2693 12294 3846 12328
rect 3880 12294 4019 12328
rect 4053 12294 5206 12328
rect 5240 12294 5280 12328
rect 1260 12238 5280 12294
rect 1260 12204 1299 12238
rect 1333 12215 2486 12238
rect 1333 12204 1400 12215
rect 1260 12181 1400 12204
rect 1434 12181 1490 12215
rect 1524 12181 1580 12215
rect 1614 12181 1670 12215
rect 1704 12181 1760 12215
rect 1794 12181 1850 12215
rect 1884 12181 1940 12215
rect 1974 12181 2030 12215
rect 2064 12181 2120 12215
rect 2154 12181 2210 12215
rect 2244 12181 2300 12215
rect 2334 12181 2390 12215
rect 2424 12204 2486 12215
rect 2520 12204 2659 12238
rect 2693 12215 3846 12238
rect 2693 12204 2760 12215
rect 2424 12181 2760 12204
rect 2794 12181 2850 12215
rect 2884 12181 2940 12215
rect 2974 12181 3030 12215
rect 3064 12181 3120 12215
rect 3154 12181 3210 12215
rect 3244 12181 3300 12215
rect 3334 12181 3390 12215
rect 3424 12181 3480 12215
rect 3514 12181 3570 12215
rect 3604 12181 3660 12215
rect 3694 12181 3750 12215
rect 3784 12204 3846 12215
rect 3880 12204 4019 12238
rect 4053 12215 5206 12238
rect 4053 12204 4120 12215
rect 3784 12181 4120 12204
rect 4154 12181 4210 12215
rect 4244 12181 4300 12215
rect 4334 12181 4390 12215
rect 4424 12181 4480 12215
rect 4514 12181 4570 12215
rect 4604 12181 4660 12215
rect 4694 12181 4750 12215
rect 4784 12181 4840 12215
rect 4874 12181 4930 12215
rect 4964 12181 5020 12215
rect 5054 12181 5110 12215
rect 5144 12204 5206 12215
rect 5240 12204 5280 12238
rect 5144 12181 5280 12204
rect 1260 12140 5280 12181
rect 2550 12074 2630 12140
rect 3910 12074 3990 12140
rect 1266 12042 5274 12074
rect 1266 12008 1400 12042
rect 1434 12008 1490 12042
rect 1524 12008 1580 12042
rect 1614 12008 1670 12042
rect 1704 12008 1760 12042
rect 1794 12008 1850 12042
rect 1884 12008 1940 12042
rect 1974 12008 2030 12042
rect 2064 12008 2120 12042
rect 2154 12008 2210 12042
rect 2244 12008 2300 12042
rect 2334 12008 2390 12042
rect 2424 12008 2760 12042
rect 2794 12008 2850 12042
rect 2884 12008 2940 12042
rect 2974 12008 3030 12042
rect 3064 12008 3120 12042
rect 3154 12008 3210 12042
rect 3244 12008 3300 12042
rect 3334 12008 3390 12042
rect 3424 12008 3480 12042
rect 3514 12008 3570 12042
rect 3604 12008 3660 12042
rect 3694 12008 3750 12042
rect 3784 12008 4120 12042
rect 4154 12008 4210 12042
rect 4244 12008 4300 12042
rect 4334 12008 4390 12042
rect 4424 12008 4480 12042
rect 4514 12008 4570 12042
rect 4604 12008 4660 12042
rect 4694 12008 4750 12042
rect 4784 12008 4840 12042
rect 4874 12008 4930 12042
rect 4964 12008 5020 12042
rect 5054 12008 5110 12042
rect 5144 12008 5274 12042
rect 1266 11975 5274 12008
rect 1266 11958 1365 11975
rect 1266 11924 1299 11958
rect 1333 11924 1365 11958
rect 1266 11868 1365 11924
rect 2455 11958 2725 11975
rect 2455 11924 2486 11958
rect 2520 11924 2659 11958
rect 2693 11924 2725 11958
rect 1266 11834 1299 11868
rect 1333 11834 1365 11868
rect 1266 11778 1365 11834
rect 1266 11744 1299 11778
rect 1333 11744 1365 11778
rect 1266 11688 1365 11744
rect 1266 11654 1299 11688
rect 1333 11654 1365 11688
rect 1266 11598 1365 11654
rect 1266 11564 1299 11598
rect 1333 11564 1365 11598
rect 1266 11508 1365 11564
rect 1266 11474 1299 11508
rect 1333 11474 1365 11508
rect 1266 11418 1365 11474
rect 1266 11384 1299 11418
rect 1333 11384 1365 11418
rect 1266 11328 1365 11384
rect 1266 11294 1299 11328
rect 1333 11294 1365 11328
rect 1266 11238 1365 11294
rect 1266 11204 1299 11238
rect 1333 11204 1365 11238
rect 1266 11148 1365 11204
rect 1266 11114 1299 11148
rect 1333 11114 1365 11148
rect 1266 11058 1365 11114
rect 1266 11030 1299 11058
rect 1260 11024 1299 11030
rect 1333 11030 1365 11058
rect 1429 11892 2391 11911
rect 1429 11858 1540 11892
rect 1574 11858 1630 11892
rect 1664 11858 1720 11892
rect 1754 11858 1810 11892
rect 1844 11858 1900 11892
rect 1934 11858 1990 11892
rect 2024 11858 2080 11892
rect 2114 11858 2170 11892
rect 2204 11858 2260 11892
rect 2294 11858 2391 11892
rect 1429 11839 2391 11858
rect 1429 11798 1501 11839
rect 1429 11764 1448 11798
rect 1482 11764 1501 11798
rect 2319 11779 2391 11839
rect 1429 11708 1501 11764
rect 1429 11674 1448 11708
rect 1482 11674 1501 11708
rect 1429 11618 1501 11674
rect 1429 11584 1448 11618
rect 1482 11584 1501 11618
rect 1429 11528 1501 11584
rect 1429 11494 1448 11528
rect 1482 11494 1501 11528
rect 1429 11438 1501 11494
rect 1429 11404 1448 11438
rect 1482 11404 1501 11438
rect 1429 11348 1501 11404
rect 1429 11314 1448 11348
rect 1482 11314 1501 11348
rect 1429 11258 1501 11314
rect 1429 11224 1448 11258
rect 1482 11224 1501 11258
rect 1429 11168 1501 11224
rect 1429 11134 1448 11168
rect 1482 11134 1501 11168
rect 1429 11078 1501 11134
rect 1563 11716 2257 11777
rect 1563 11682 1622 11716
rect 1656 11704 1712 11716
rect 1684 11682 1712 11704
rect 1746 11704 1802 11716
rect 1746 11682 1750 11704
rect 1563 11670 1650 11682
rect 1684 11670 1750 11682
rect 1784 11682 1802 11704
rect 1836 11704 1892 11716
rect 1836 11682 1850 11704
rect 1784 11670 1850 11682
rect 1884 11682 1892 11704
rect 1926 11704 1982 11716
rect 2016 11704 2072 11716
rect 2106 11704 2162 11716
rect 1926 11682 1950 11704
rect 2016 11682 2050 11704
rect 2106 11682 2150 11704
rect 2196 11682 2257 11716
rect 1884 11670 1950 11682
rect 1984 11670 2050 11682
rect 2084 11670 2150 11682
rect 2184 11670 2257 11682
rect 1563 11626 2257 11670
rect 1563 11592 1622 11626
rect 1656 11604 1712 11626
rect 1684 11592 1712 11604
rect 1746 11604 1802 11626
rect 1746 11592 1750 11604
rect 1563 11570 1650 11592
rect 1684 11570 1750 11592
rect 1784 11592 1802 11604
rect 1836 11604 1892 11626
rect 1836 11592 1850 11604
rect 1784 11570 1850 11592
rect 1884 11592 1892 11604
rect 1926 11604 1982 11626
rect 2016 11604 2072 11626
rect 2106 11604 2162 11626
rect 1926 11592 1950 11604
rect 2016 11592 2050 11604
rect 2106 11592 2150 11604
rect 2196 11592 2257 11626
rect 1884 11570 1950 11592
rect 1984 11570 2050 11592
rect 2084 11570 2150 11592
rect 2184 11570 2257 11592
rect 1563 11536 2257 11570
rect 1563 11502 1622 11536
rect 1656 11504 1712 11536
rect 1684 11502 1712 11504
rect 1746 11504 1802 11536
rect 1746 11502 1750 11504
rect 1563 11470 1650 11502
rect 1684 11470 1750 11502
rect 1784 11502 1802 11504
rect 1836 11504 1892 11536
rect 1836 11502 1850 11504
rect 1784 11470 1850 11502
rect 1884 11502 1892 11504
rect 1926 11504 1982 11536
rect 2016 11504 2072 11536
rect 2106 11504 2162 11536
rect 1926 11502 1950 11504
rect 2016 11502 2050 11504
rect 2106 11502 2150 11504
rect 2196 11502 2257 11536
rect 1884 11470 1950 11502
rect 1984 11470 2050 11502
rect 2084 11470 2150 11502
rect 2184 11470 2257 11502
rect 1563 11446 2257 11470
rect 1563 11412 1622 11446
rect 1656 11412 1712 11446
rect 1746 11412 1802 11446
rect 1836 11412 1892 11446
rect 1926 11412 1982 11446
rect 2016 11412 2072 11446
rect 2106 11412 2162 11446
rect 2196 11412 2257 11446
rect 1563 11404 2257 11412
rect 1563 11370 1650 11404
rect 1684 11370 1750 11404
rect 1784 11370 1850 11404
rect 1884 11370 1950 11404
rect 1984 11370 2050 11404
rect 2084 11370 2150 11404
rect 2184 11370 2257 11404
rect 1563 11356 2257 11370
rect 1563 11322 1622 11356
rect 1656 11322 1712 11356
rect 1746 11322 1802 11356
rect 1836 11322 1892 11356
rect 1926 11322 1982 11356
rect 2016 11322 2072 11356
rect 2106 11322 2162 11356
rect 2196 11322 2257 11356
rect 1563 11304 2257 11322
rect 1563 11270 1650 11304
rect 1684 11270 1750 11304
rect 1784 11270 1850 11304
rect 1884 11270 1950 11304
rect 1984 11270 2050 11304
rect 2084 11270 2150 11304
rect 2184 11270 2257 11304
rect 1563 11266 2257 11270
rect 1563 11232 1622 11266
rect 1656 11232 1712 11266
rect 1746 11232 1802 11266
rect 1836 11232 1892 11266
rect 1926 11232 1982 11266
rect 2016 11232 2072 11266
rect 2106 11232 2162 11266
rect 2196 11232 2257 11266
rect 1563 11204 2257 11232
rect 1563 11176 1650 11204
rect 1684 11176 1750 11204
rect 1563 11142 1622 11176
rect 1684 11170 1712 11176
rect 1656 11142 1712 11170
rect 1746 11170 1750 11176
rect 1784 11176 1850 11204
rect 1784 11170 1802 11176
rect 1746 11142 1802 11170
rect 1836 11170 1850 11176
rect 1884 11176 1950 11204
rect 1984 11176 2050 11204
rect 2084 11176 2150 11204
rect 2184 11176 2257 11204
rect 1884 11170 1892 11176
rect 1836 11142 1892 11170
rect 1926 11170 1950 11176
rect 2016 11170 2050 11176
rect 2106 11170 2150 11176
rect 1926 11142 1982 11170
rect 2016 11142 2072 11170
rect 2106 11142 2162 11170
rect 2196 11142 2257 11176
rect 1563 11083 2257 11142
rect 2319 11745 2338 11779
rect 2372 11745 2391 11779
rect 2319 11689 2391 11745
rect 2319 11655 2338 11689
rect 2372 11655 2391 11689
rect 2319 11599 2391 11655
rect 2319 11565 2338 11599
rect 2372 11565 2391 11599
rect 2319 11509 2391 11565
rect 2319 11475 2338 11509
rect 2372 11475 2391 11509
rect 2319 11419 2391 11475
rect 2319 11385 2338 11419
rect 2372 11385 2391 11419
rect 2319 11329 2391 11385
rect 2319 11295 2338 11329
rect 2372 11295 2391 11329
rect 2319 11239 2391 11295
rect 2319 11205 2338 11239
rect 2372 11205 2391 11239
rect 2319 11149 2391 11205
rect 2319 11115 2338 11149
rect 2372 11115 2391 11149
rect 1429 11044 1448 11078
rect 1482 11044 1501 11078
rect 1429 11030 1501 11044
rect 2319 11059 2391 11115
rect 2319 11030 2338 11059
rect 1333 11025 2338 11030
rect 2372 11030 2391 11059
rect 2455 11868 2725 11924
rect 3815 11958 4085 11975
rect 3815 11924 3846 11958
rect 3880 11924 4019 11958
rect 4053 11924 4085 11958
rect 2455 11834 2486 11868
rect 2520 11834 2659 11868
rect 2693 11834 2725 11868
rect 2455 11778 2725 11834
rect 2455 11744 2486 11778
rect 2520 11744 2659 11778
rect 2693 11744 2725 11778
rect 2455 11688 2725 11744
rect 2455 11654 2486 11688
rect 2520 11654 2659 11688
rect 2693 11654 2725 11688
rect 2455 11598 2725 11654
rect 2455 11564 2486 11598
rect 2520 11564 2659 11598
rect 2693 11564 2725 11598
rect 2455 11508 2725 11564
rect 2455 11474 2486 11508
rect 2520 11474 2659 11508
rect 2693 11474 2725 11508
rect 2455 11418 2725 11474
rect 2455 11384 2486 11418
rect 2520 11384 2659 11418
rect 2693 11384 2725 11418
rect 2455 11328 2725 11384
rect 2455 11294 2486 11328
rect 2520 11294 2659 11328
rect 2693 11294 2725 11328
rect 2455 11238 2725 11294
rect 2455 11204 2486 11238
rect 2520 11204 2659 11238
rect 2693 11204 2725 11238
rect 2455 11148 2725 11204
rect 2455 11114 2486 11148
rect 2520 11114 2659 11148
rect 2693 11114 2725 11148
rect 2455 11058 2725 11114
rect 2455 11030 2486 11058
rect 2372 11025 2486 11030
rect 1333 11024 2486 11025
rect 2520 11024 2659 11058
rect 2693 11030 2725 11058
rect 2789 11892 3751 11911
rect 2789 11858 2900 11892
rect 2934 11858 2990 11892
rect 3024 11858 3080 11892
rect 3114 11858 3170 11892
rect 3204 11858 3260 11892
rect 3294 11858 3350 11892
rect 3384 11858 3440 11892
rect 3474 11858 3530 11892
rect 3564 11858 3620 11892
rect 3654 11858 3751 11892
rect 2789 11839 3751 11858
rect 2789 11798 2861 11839
rect 2789 11764 2808 11798
rect 2842 11764 2861 11798
rect 3679 11779 3751 11839
rect 2789 11708 2861 11764
rect 2789 11674 2808 11708
rect 2842 11674 2861 11708
rect 2789 11618 2861 11674
rect 2789 11584 2808 11618
rect 2842 11584 2861 11618
rect 2789 11528 2861 11584
rect 2789 11494 2808 11528
rect 2842 11494 2861 11528
rect 2789 11438 2861 11494
rect 2789 11404 2808 11438
rect 2842 11404 2861 11438
rect 2789 11348 2861 11404
rect 2789 11314 2808 11348
rect 2842 11314 2861 11348
rect 2789 11258 2861 11314
rect 2789 11224 2808 11258
rect 2842 11224 2861 11258
rect 2789 11168 2861 11224
rect 2789 11134 2808 11168
rect 2842 11134 2861 11168
rect 2789 11078 2861 11134
rect 2923 11716 3617 11777
rect 2923 11682 2982 11716
rect 3016 11704 3072 11716
rect 3044 11682 3072 11704
rect 3106 11704 3162 11716
rect 3106 11682 3110 11704
rect 2923 11670 3010 11682
rect 3044 11670 3110 11682
rect 3144 11682 3162 11704
rect 3196 11704 3252 11716
rect 3196 11682 3210 11704
rect 3144 11670 3210 11682
rect 3244 11682 3252 11704
rect 3286 11704 3342 11716
rect 3376 11704 3432 11716
rect 3466 11704 3522 11716
rect 3286 11682 3310 11704
rect 3376 11682 3410 11704
rect 3466 11682 3510 11704
rect 3556 11682 3617 11716
rect 3244 11670 3310 11682
rect 3344 11670 3410 11682
rect 3444 11670 3510 11682
rect 3544 11670 3617 11682
rect 2923 11626 3617 11670
rect 2923 11592 2982 11626
rect 3016 11604 3072 11626
rect 3044 11592 3072 11604
rect 3106 11604 3162 11626
rect 3106 11592 3110 11604
rect 2923 11570 3010 11592
rect 3044 11570 3110 11592
rect 3144 11592 3162 11604
rect 3196 11604 3252 11626
rect 3196 11592 3210 11604
rect 3144 11570 3210 11592
rect 3244 11592 3252 11604
rect 3286 11604 3342 11626
rect 3376 11604 3432 11626
rect 3466 11604 3522 11626
rect 3286 11592 3310 11604
rect 3376 11592 3410 11604
rect 3466 11592 3510 11604
rect 3556 11592 3617 11626
rect 3244 11570 3310 11592
rect 3344 11570 3410 11592
rect 3444 11570 3510 11592
rect 3544 11570 3617 11592
rect 2923 11536 3617 11570
rect 2923 11502 2982 11536
rect 3016 11504 3072 11536
rect 3044 11502 3072 11504
rect 3106 11504 3162 11536
rect 3106 11502 3110 11504
rect 2923 11470 3010 11502
rect 3044 11470 3110 11502
rect 3144 11502 3162 11504
rect 3196 11504 3252 11536
rect 3196 11502 3210 11504
rect 3144 11470 3210 11502
rect 3244 11502 3252 11504
rect 3286 11504 3342 11536
rect 3376 11504 3432 11536
rect 3466 11504 3522 11536
rect 3286 11502 3310 11504
rect 3376 11502 3410 11504
rect 3466 11502 3510 11504
rect 3556 11502 3617 11536
rect 3244 11470 3310 11502
rect 3344 11470 3410 11502
rect 3444 11470 3510 11502
rect 3544 11470 3617 11502
rect 2923 11446 3617 11470
rect 2923 11412 2982 11446
rect 3016 11412 3072 11446
rect 3106 11412 3162 11446
rect 3196 11412 3252 11446
rect 3286 11412 3342 11446
rect 3376 11412 3432 11446
rect 3466 11412 3522 11446
rect 3556 11412 3617 11446
rect 2923 11404 3617 11412
rect 2923 11370 3010 11404
rect 3044 11370 3110 11404
rect 3144 11370 3210 11404
rect 3244 11370 3310 11404
rect 3344 11370 3410 11404
rect 3444 11370 3510 11404
rect 3544 11370 3617 11404
rect 2923 11356 3617 11370
rect 2923 11322 2982 11356
rect 3016 11322 3072 11356
rect 3106 11322 3162 11356
rect 3196 11322 3252 11356
rect 3286 11322 3342 11356
rect 3376 11322 3432 11356
rect 3466 11322 3522 11356
rect 3556 11322 3617 11356
rect 2923 11304 3617 11322
rect 2923 11270 3010 11304
rect 3044 11270 3110 11304
rect 3144 11270 3210 11304
rect 3244 11270 3310 11304
rect 3344 11270 3410 11304
rect 3444 11270 3510 11304
rect 3544 11270 3617 11304
rect 2923 11266 3617 11270
rect 2923 11232 2982 11266
rect 3016 11232 3072 11266
rect 3106 11232 3162 11266
rect 3196 11232 3252 11266
rect 3286 11232 3342 11266
rect 3376 11232 3432 11266
rect 3466 11232 3522 11266
rect 3556 11232 3617 11266
rect 2923 11204 3617 11232
rect 2923 11176 3010 11204
rect 3044 11176 3110 11204
rect 2923 11142 2982 11176
rect 3044 11170 3072 11176
rect 3016 11142 3072 11170
rect 3106 11170 3110 11176
rect 3144 11176 3210 11204
rect 3144 11170 3162 11176
rect 3106 11142 3162 11170
rect 3196 11170 3210 11176
rect 3244 11176 3310 11204
rect 3344 11176 3410 11204
rect 3444 11176 3510 11204
rect 3544 11176 3617 11204
rect 3244 11170 3252 11176
rect 3196 11142 3252 11170
rect 3286 11170 3310 11176
rect 3376 11170 3410 11176
rect 3466 11170 3510 11176
rect 3286 11142 3342 11170
rect 3376 11142 3432 11170
rect 3466 11142 3522 11170
rect 3556 11142 3617 11176
rect 2923 11083 3617 11142
rect 3679 11745 3698 11779
rect 3732 11745 3751 11779
rect 3679 11689 3751 11745
rect 3679 11655 3698 11689
rect 3732 11655 3751 11689
rect 3679 11599 3751 11655
rect 3679 11565 3698 11599
rect 3732 11565 3751 11599
rect 3679 11509 3751 11565
rect 3679 11475 3698 11509
rect 3732 11475 3751 11509
rect 3679 11419 3751 11475
rect 3679 11385 3698 11419
rect 3732 11385 3751 11419
rect 3679 11329 3751 11385
rect 3679 11295 3698 11329
rect 3732 11295 3751 11329
rect 3679 11239 3751 11295
rect 3679 11205 3698 11239
rect 3732 11205 3751 11239
rect 3679 11149 3751 11205
rect 3679 11115 3698 11149
rect 3732 11115 3751 11149
rect 2789 11044 2808 11078
rect 2842 11044 2861 11078
rect 2789 11030 2861 11044
rect 3679 11059 3751 11115
rect 3679 11030 3698 11059
rect 2693 11025 3698 11030
rect 3732 11030 3751 11059
rect 3815 11868 4085 11924
rect 5175 11958 5274 11975
rect 5175 11924 5206 11958
rect 5240 11924 5274 11958
rect 3815 11834 3846 11868
rect 3880 11834 4019 11868
rect 4053 11834 4085 11868
rect 3815 11778 4085 11834
rect 3815 11744 3846 11778
rect 3880 11744 4019 11778
rect 4053 11744 4085 11778
rect 3815 11688 4085 11744
rect 3815 11654 3846 11688
rect 3880 11654 4019 11688
rect 4053 11654 4085 11688
rect 3815 11598 4085 11654
rect 3815 11564 3846 11598
rect 3880 11564 4019 11598
rect 4053 11564 4085 11598
rect 3815 11508 4085 11564
rect 3815 11474 3846 11508
rect 3880 11474 4019 11508
rect 4053 11474 4085 11508
rect 3815 11418 4085 11474
rect 3815 11384 3846 11418
rect 3880 11384 4019 11418
rect 4053 11384 4085 11418
rect 3815 11328 4085 11384
rect 3815 11294 3846 11328
rect 3880 11294 4019 11328
rect 4053 11294 4085 11328
rect 3815 11238 4085 11294
rect 3815 11204 3846 11238
rect 3880 11204 4019 11238
rect 4053 11204 4085 11238
rect 3815 11148 4085 11204
rect 3815 11114 3846 11148
rect 3880 11114 4019 11148
rect 4053 11114 4085 11148
rect 3815 11058 4085 11114
rect 3815 11030 3846 11058
rect 3732 11025 3846 11030
rect 2693 11024 3846 11025
rect 3880 11024 4019 11058
rect 4053 11030 4085 11058
rect 4149 11892 5111 11911
rect 4149 11858 4260 11892
rect 4294 11858 4350 11892
rect 4384 11858 4440 11892
rect 4474 11858 4530 11892
rect 4564 11858 4620 11892
rect 4654 11858 4710 11892
rect 4744 11858 4800 11892
rect 4834 11858 4890 11892
rect 4924 11858 4980 11892
rect 5014 11858 5111 11892
rect 4149 11839 5111 11858
rect 4149 11798 4221 11839
rect 4149 11764 4168 11798
rect 4202 11764 4221 11798
rect 5039 11779 5111 11839
rect 4149 11708 4221 11764
rect 4149 11674 4168 11708
rect 4202 11674 4221 11708
rect 4149 11618 4221 11674
rect 4149 11584 4168 11618
rect 4202 11584 4221 11618
rect 4149 11528 4221 11584
rect 4149 11494 4168 11528
rect 4202 11494 4221 11528
rect 4149 11438 4221 11494
rect 4149 11404 4168 11438
rect 4202 11404 4221 11438
rect 4149 11348 4221 11404
rect 4149 11314 4168 11348
rect 4202 11314 4221 11348
rect 4149 11258 4221 11314
rect 4149 11224 4168 11258
rect 4202 11224 4221 11258
rect 4149 11168 4221 11224
rect 4149 11134 4168 11168
rect 4202 11134 4221 11168
rect 4149 11078 4221 11134
rect 4283 11716 4977 11777
rect 4283 11682 4342 11716
rect 4376 11704 4432 11716
rect 4404 11682 4432 11704
rect 4466 11704 4522 11716
rect 4466 11682 4470 11704
rect 4283 11670 4370 11682
rect 4404 11670 4470 11682
rect 4504 11682 4522 11704
rect 4556 11704 4612 11716
rect 4556 11682 4570 11704
rect 4504 11670 4570 11682
rect 4604 11682 4612 11704
rect 4646 11704 4702 11716
rect 4736 11704 4792 11716
rect 4826 11704 4882 11716
rect 4646 11682 4670 11704
rect 4736 11682 4770 11704
rect 4826 11682 4870 11704
rect 4916 11682 4977 11716
rect 4604 11670 4670 11682
rect 4704 11670 4770 11682
rect 4804 11670 4870 11682
rect 4904 11670 4977 11682
rect 4283 11626 4977 11670
rect 4283 11592 4342 11626
rect 4376 11604 4432 11626
rect 4404 11592 4432 11604
rect 4466 11604 4522 11626
rect 4466 11592 4470 11604
rect 4283 11570 4370 11592
rect 4404 11570 4470 11592
rect 4504 11592 4522 11604
rect 4556 11604 4612 11626
rect 4556 11592 4570 11604
rect 4504 11570 4570 11592
rect 4604 11592 4612 11604
rect 4646 11604 4702 11626
rect 4736 11604 4792 11626
rect 4826 11604 4882 11626
rect 4646 11592 4670 11604
rect 4736 11592 4770 11604
rect 4826 11592 4870 11604
rect 4916 11592 4977 11626
rect 4604 11570 4670 11592
rect 4704 11570 4770 11592
rect 4804 11570 4870 11592
rect 4904 11570 4977 11592
rect 4283 11536 4977 11570
rect 4283 11502 4342 11536
rect 4376 11504 4432 11536
rect 4404 11502 4432 11504
rect 4466 11504 4522 11536
rect 4466 11502 4470 11504
rect 4283 11470 4370 11502
rect 4404 11470 4470 11502
rect 4504 11502 4522 11504
rect 4556 11504 4612 11536
rect 4556 11502 4570 11504
rect 4504 11470 4570 11502
rect 4604 11502 4612 11504
rect 4646 11504 4702 11536
rect 4736 11504 4792 11536
rect 4826 11504 4882 11536
rect 4646 11502 4670 11504
rect 4736 11502 4770 11504
rect 4826 11502 4870 11504
rect 4916 11502 4977 11536
rect 4604 11470 4670 11502
rect 4704 11470 4770 11502
rect 4804 11470 4870 11502
rect 4904 11470 4977 11502
rect 4283 11446 4977 11470
rect 4283 11412 4342 11446
rect 4376 11412 4432 11446
rect 4466 11412 4522 11446
rect 4556 11412 4612 11446
rect 4646 11412 4702 11446
rect 4736 11412 4792 11446
rect 4826 11412 4882 11446
rect 4916 11412 4977 11446
rect 4283 11404 4977 11412
rect 4283 11370 4370 11404
rect 4404 11370 4470 11404
rect 4504 11370 4570 11404
rect 4604 11370 4670 11404
rect 4704 11370 4770 11404
rect 4804 11370 4870 11404
rect 4904 11370 4977 11404
rect 4283 11356 4977 11370
rect 4283 11322 4342 11356
rect 4376 11322 4432 11356
rect 4466 11322 4522 11356
rect 4556 11322 4612 11356
rect 4646 11322 4702 11356
rect 4736 11322 4792 11356
rect 4826 11322 4882 11356
rect 4916 11322 4977 11356
rect 4283 11304 4977 11322
rect 4283 11270 4370 11304
rect 4404 11270 4470 11304
rect 4504 11270 4570 11304
rect 4604 11270 4670 11304
rect 4704 11270 4770 11304
rect 4804 11270 4870 11304
rect 4904 11270 4977 11304
rect 4283 11266 4977 11270
rect 4283 11232 4342 11266
rect 4376 11232 4432 11266
rect 4466 11232 4522 11266
rect 4556 11232 4612 11266
rect 4646 11232 4702 11266
rect 4736 11232 4792 11266
rect 4826 11232 4882 11266
rect 4916 11232 4977 11266
rect 4283 11204 4977 11232
rect 4283 11176 4370 11204
rect 4404 11176 4470 11204
rect 4283 11142 4342 11176
rect 4404 11170 4432 11176
rect 4376 11142 4432 11170
rect 4466 11170 4470 11176
rect 4504 11176 4570 11204
rect 4504 11170 4522 11176
rect 4466 11142 4522 11170
rect 4556 11170 4570 11176
rect 4604 11176 4670 11204
rect 4704 11176 4770 11204
rect 4804 11176 4870 11204
rect 4904 11176 4977 11204
rect 4604 11170 4612 11176
rect 4556 11142 4612 11170
rect 4646 11170 4670 11176
rect 4736 11170 4770 11176
rect 4826 11170 4870 11176
rect 4646 11142 4702 11170
rect 4736 11142 4792 11170
rect 4826 11142 4882 11170
rect 4916 11142 4977 11176
rect 4283 11083 4977 11142
rect 5039 11745 5058 11779
rect 5092 11745 5111 11779
rect 5039 11689 5111 11745
rect 5039 11655 5058 11689
rect 5092 11655 5111 11689
rect 5039 11599 5111 11655
rect 5039 11565 5058 11599
rect 5092 11565 5111 11599
rect 5039 11509 5111 11565
rect 5039 11475 5058 11509
rect 5092 11475 5111 11509
rect 5039 11419 5111 11475
rect 5039 11385 5058 11419
rect 5092 11385 5111 11419
rect 5039 11329 5111 11385
rect 5039 11295 5058 11329
rect 5092 11295 5111 11329
rect 5039 11239 5111 11295
rect 5039 11205 5058 11239
rect 5092 11205 5111 11239
rect 5039 11149 5111 11205
rect 5039 11115 5058 11149
rect 5092 11115 5111 11149
rect 4149 11044 4168 11078
rect 4202 11044 4221 11078
rect 4149 11030 4221 11044
rect 5039 11059 5111 11115
rect 5039 11030 5058 11059
rect 4053 11025 5058 11030
rect 5092 11030 5111 11059
rect 5175 11868 5274 11924
rect 5175 11834 5206 11868
rect 5240 11834 5274 11868
rect 5175 11778 5274 11834
rect 5175 11744 5206 11778
rect 5240 11744 5274 11778
rect 5175 11688 5274 11744
rect 5175 11654 5206 11688
rect 5240 11654 5274 11688
rect 5175 11598 5274 11654
rect 5175 11564 5206 11598
rect 5240 11564 5274 11598
rect 5175 11508 5274 11564
rect 5175 11474 5206 11508
rect 5240 11474 5274 11508
rect 5175 11418 5274 11474
rect 5175 11384 5206 11418
rect 5240 11384 5274 11418
rect 5175 11328 5274 11384
rect 5175 11294 5206 11328
rect 5240 11294 5274 11328
rect 5175 11238 5274 11294
rect 5175 11204 5206 11238
rect 5240 11204 5274 11238
rect 5175 11148 5274 11204
rect 5175 11114 5206 11148
rect 5240 11114 5274 11148
rect 5175 11058 5274 11114
rect 5175 11030 5206 11058
rect 5092 11025 5206 11030
rect 4053 11024 5206 11025
rect 5240 11030 5274 11058
rect 5240 11024 5280 11030
rect 1260 11002 5280 11024
rect 1260 10968 1506 11002
rect 1540 10968 1596 11002
rect 1630 10968 1686 11002
rect 1720 10968 1776 11002
rect 1810 10968 1866 11002
rect 1900 10968 1956 11002
rect 1990 10968 2046 11002
rect 2080 10968 2136 11002
rect 2170 10968 2226 11002
rect 2260 10968 2866 11002
rect 2900 10968 2956 11002
rect 2990 10968 3046 11002
rect 3080 10968 3136 11002
rect 3170 10968 3226 11002
rect 3260 10968 3316 11002
rect 3350 10968 3406 11002
rect 3440 10968 3496 11002
rect 3530 10968 3586 11002
rect 3620 10968 4226 11002
rect 4260 10968 4316 11002
rect 4350 10968 4406 11002
rect 4440 10968 4496 11002
rect 4530 10968 4586 11002
rect 4620 10968 4676 11002
rect 4710 10968 4766 11002
rect 4800 10968 4856 11002
rect 4890 10968 4946 11002
rect 4980 10968 5280 11002
rect 1260 10934 1299 10968
rect 1333 10934 2486 10968
rect 2520 10934 2659 10968
rect 2693 10934 3846 10968
rect 3880 10934 4019 10968
rect 4053 10934 5206 10968
rect 5240 10934 5280 10968
rect 1260 10878 5280 10934
rect 1260 10844 1299 10878
rect 1333 10855 2486 10878
rect 1333 10844 1400 10855
rect 1260 10821 1400 10844
rect 1434 10821 1490 10855
rect 1524 10821 1580 10855
rect 1614 10821 1670 10855
rect 1704 10821 1760 10855
rect 1794 10821 1850 10855
rect 1884 10821 1940 10855
rect 1974 10821 2030 10855
rect 2064 10821 2120 10855
rect 2154 10821 2210 10855
rect 2244 10821 2300 10855
rect 2334 10821 2390 10855
rect 2424 10844 2486 10855
rect 2520 10844 2659 10878
rect 2693 10855 3846 10878
rect 2693 10844 2760 10855
rect 2424 10821 2760 10844
rect 2794 10821 2850 10855
rect 2884 10821 2940 10855
rect 2974 10821 3030 10855
rect 3064 10821 3120 10855
rect 3154 10821 3210 10855
rect 3244 10821 3300 10855
rect 3334 10821 3390 10855
rect 3424 10821 3480 10855
rect 3514 10821 3570 10855
rect 3604 10821 3660 10855
rect 3694 10821 3750 10855
rect 3784 10844 3846 10855
rect 3880 10844 4019 10878
rect 4053 10855 5206 10878
rect 4053 10844 4120 10855
rect 3784 10821 4120 10844
rect 4154 10821 4210 10855
rect 4244 10821 4300 10855
rect 4334 10821 4390 10855
rect 4424 10821 4480 10855
rect 4514 10821 4570 10855
rect 4604 10821 4660 10855
rect 4694 10821 4750 10855
rect 4784 10821 4840 10855
rect 4874 10821 4930 10855
rect 4964 10821 5020 10855
rect 5054 10821 5110 10855
rect 5144 10844 5206 10855
rect 5240 10844 5280 10878
rect 5144 10821 5280 10844
rect 1260 10780 5280 10821
rect 2532 10610 2622 10620
rect 2532 10560 2552 10610
rect 2602 10560 2622 10610
rect 2532 10550 2622 10560
rect 3930 10610 4020 10620
rect 3930 10560 3950 10610
rect 4000 10560 4020 10610
rect 3930 10550 4020 10560
rect 1160 10260 1220 10280
rect 1160 10230 1170 10260
rect 1070 10220 1170 10230
rect 1210 10220 1220 10260
rect 1070 10210 1220 10220
rect 1070 10170 1090 10210
rect 1130 10170 1220 10210
rect 1070 10160 1220 10170
rect 1070 10150 1170 10160
rect 1160 10120 1170 10150
rect 1210 10120 1220 10160
rect 1160 10100 1220 10120
rect 3240 10260 3300 10280
rect 3240 10220 3250 10260
rect 3290 10220 3300 10260
rect 3240 10160 3300 10220
rect 3240 10120 3250 10160
rect 3290 10120 3300 10160
rect 3240 10100 3300 10120
rect 5320 10270 5460 10280
rect 5320 10260 5540 10270
rect 5320 10220 5330 10260
rect 5370 10220 5410 10260
rect 5450 10250 5540 10260
rect 5450 10220 5480 10250
rect 5320 10210 5480 10220
rect 5520 10210 5540 10250
rect 5320 10170 5540 10210
rect 5320 10160 5480 10170
rect 5320 10120 5330 10160
rect 5370 10120 5410 10160
rect 5450 10130 5480 10160
rect 5520 10130 5540 10170
rect 5450 10120 5540 10130
rect 5320 10110 5540 10120
rect 5320 10100 5460 10110
rect 1170 10060 1210 10100
rect 3250 10060 3290 10100
rect 1150 10040 1230 10060
rect 1150 10000 1170 10040
rect 1210 10000 1230 10040
rect 1150 9980 1230 10000
rect 1310 10040 1390 10060
rect 1310 10000 1330 10040
rect 1370 10000 1390 10040
rect 1310 9980 1390 10000
rect 1470 10040 1550 10060
rect 1470 10000 1490 10040
rect 1530 10000 1550 10040
rect 1470 9980 1550 10000
rect 1630 10040 1710 10060
rect 1630 10000 1650 10040
rect 1690 10000 1710 10040
rect 1630 9980 1710 10000
rect 1790 10040 1870 10060
rect 1790 10000 1810 10040
rect 1850 10000 1870 10040
rect 1790 9980 1870 10000
rect 1950 10040 2030 10060
rect 1950 10000 1970 10040
rect 2010 10000 2030 10040
rect 1950 9980 2030 10000
rect 2110 10040 2190 10060
rect 2110 10000 2130 10040
rect 2170 10000 2190 10040
rect 2110 9980 2190 10000
rect 2270 10040 2350 10060
rect 2270 10000 2290 10040
rect 2330 10000 2350 10040
rect 2270 9980 2350 10000
rect 2430 10040 2510 10060
rect 2430 10000 2450 10040
rect 2490 10000 2510 10040
rect 2430 9980 2510 10000
rect 2590 10040 2670 10060
rect 2590 10000 2610 10040
rect 2650 10000 2670 10040
rect 2590 9980 2670 10000
rect 2750 10040 2830 10060
rect 2750 10000 2770 10040
rect 2810 10000 2830 10040
rect 2750 9980 2830 10000
rect 2910 10040 2990 10060
rect 2910 10000 2930 10040
rect 2970 10000 2990 10040
rect 2910 9980 2990 10000
rect 3070 10040 3150 10060
rect 3070 10000 3090 10040
rect 3130 10000 3150 10040
rect 3070 9980 3150 10000
rect 3230 10040 3310 10060
rect 3230 10000 3250 10040
rect 3290 10000 3310 10040
rect 3230 9980 3310 10000
rect 3390 10040 3470 10060
rect 3390 10000 3410 10040
rect 3450 10000 3470 10040
rect 3390 9980 3470 10000
rect 3550 10040 3630 10060
rect 3550 10000 3570 10040
rect 3610 10000 3630 10040
rect 3550 9980 3630 10000
rect 3710 10040 3790 10060
rect 3710 10000 3730 10040
rect 3770 10000 3790 10040
rect 3710 9980 3790 10000
rect 3870 10040 3950 10060
rect 3870 10000 3890 10040
rect 3930 10000 3950 10040
rect 3870 9980 3950 10000
rect 4030 10040 4110 10060
rect 4030 10000 4050 10040
rect 4090 10000 4110 10040
rect 4030 9980 4110 10000
rect 4190 10040 4270 10060
rect 4190 10000 4210 10040
rect 4250 10000 4270 10040
rect 4190 9980 4270 10000
rect 4350 10040 4430 10060
rect 4350 10000 4370 10040
rect 4410 10000 4430 10040
rect 4350 9980 4430 10000
rect 4510 10040 4590 10060
rect 4510 10000 4530 10040
rect 4570 10000 4590 10040
rect 4510 9980 4590 10000
rect 4670 10040 4750 10060
rect 4670 10000 4690 10040
rect 4730 10000 4750 10040
rect 4670 9980 4750 10000
rect 4830 10040 4910 10060
rect 4830 10000 4850 10040
rect 4890 10000 4910 10040
rect 4830 9980 4910 10000
rect 4990 10040 5070 10060
rect 4990 10000 5010 10040
rect 5050 10000 5070 10040
rect 4990 9980 5070 10000
rect 5150 10040 5230 10060
rect 5150 10000 5170 10040
rect 5210 10000 5230 10040
rect 5150 9980 5230 10000
rect 11750 9810 11850 9830
rect 11750 9790 11770 9810
rect 1890 9770 1970 9790
rect 1890 9730 1910 9770
rect 1950 9730 1970 9770
rect 1890 9710 1970 9730
rect 4570 9770 4650 9790
rect 4570 9730 4590 9770
rect 4630 9730 4650 9770
rect 4570 9710 4650 9730
rect 11670 9750 11770 9790
rect 11830 9750 11850 9810
rect 1910 9670 1950 9710
rect 4590 9670 4630 9710
rect 740 9650 800 9670
rect 740 9610 750 9650
rect 790 9610 800 9650
rect 740 9550 800 9610
rect 740 9510 750 9550
rect 790 9510 800 9550
rect 740 9450 800 9510
rect 740 9410 750 9450
rect 790 9410 800 9450
rect 740 9350 800 9410
rect 740 9310 750 9350
rect 790 9310 800 9350
rect 740 9250 800 9310
rect 740 9210 750 9250
rect 790 9210 800 9250
rect 740 9190 800 9210
rect 1820 9650 2040 9670
rect 1820 9610 1830 9650
rect 1870 9610 1910 9650
rect 1950 9610 1990 9650
rect 2030 9610 2040 9650
rect 1820 9550 2040 9610
rect 1820 9510 1830 9550
rect 1870 9510 1910 9550
rect 1950 9510 1990 9550
rect 2030 9510 2040 9550
rect 1820 9450 2040 9510
rect 1820 9410 1830 9450
rect 1870 9410 1910 9450
rect 1950 9410 1990 9450
rect 2030 9410 2040 9450
rect 1820 9350 2040 9410
rect 1820 9310 1830 9350
rect 1870 9310 1910 9350
rect 1950 9310 1990 9350
rect 2030 9310 2040 9350
rect 1820 9250 2040 9310
rect 1820 9210 1830 9250
rect 1870 9210 1910 9250
rect 1950 9210 1990 9250
rect 2030 9210 2040 9250
rect 1820 9190 2040 9210
rect 3060 9650 3120 9670
rect 3060 9610 3070 9650
rect 3110 9610 3120 9650
rect 3060 9550 3120 9610
rect 3060 9510 3070 9550
rect 3110 9510 3120 9550
rect 3060 9450 3120 9510
rect 3060 9410 3070 9450
rect 3110 9410 3120 9450
rect 3060 9350 3120 9410
rect 3060 9310 3070 9350
rect 3110 9310 3120 9350
rect 3060 9250 3120 9310
rect 3060 9210 3070 9250
rect 3110 9210 3120 9250
rect 730 9170 810 9190
rect 730 9130 750 9170
rect 790 9130 810 9170
rect 3060 9160 3120 9210
rect 730 9110 810 9130
rect 910 9130 990 9150
rect 910 9090 930 9130
rect 970 9090 990 9130
rect 910 9070 990 9090
rect 1150 9130 1230 9150
rect 1150 9090 1170 9130
rect 1210 9090 1230 9130
rect 1150 9070 1230 9090
rect 1390 9130 1470 9150
rect 1390 9090 1410 9130
rect 1450 9090 1470 9130
rect 1390 9070 1470 9090
rect 1630 9130 1710 9150
rect 1630 9090 1650 9130
rect 1690 9090 1710 9130
rect 1630 9070 1710 9090
rect 2270 9130 2350 9150
rect 2270 9090 2290 9130
rect 2330 9090 2350 9130
rect 2270 9070 2350 9090
rect 2510 9130 2590 9150
rect 2510 9090 2530 9130
rect 2570 9090 2590 9130
rect 2510 9070 2590 9090
rect 2750 9130 2830 9150
rect 2750 9090 2770 9130
rect 2810 9090 2830 9130
rect 3060 9120 3070 9160
rect 3110 9120 3120 9160
rect 3060 9100 3120 9120
rect 3420 9650 3480 9670
rect 3420 9610 3430 9650
rect 3470 9610 3480 9650
rect 3420 9550 3480 9610
rect 3420 9510 3430 9550
rect 3470 9510 3480 9550
rect 3420 9450 3480 9510
rect 3420 9410 3430 9450
rect 3470 9410 3480 9450
rect 3420 9350 3480 9410
rect 3420 9310 3430 9350
rect 3470 9310 3480 9350
rect 3420 9250 3480 9310
rect 3420 9210 3430 9250
rect 3470 9210 3480 9250
rect 3420 9160 3480 9210
rect 4500 9650 4720 9670
rect 4500 9610 4510 9650
rect 4550 9610 4590 9650
rect 4630 9610 4670 9650
rect 4710 9610 4720 9650
rect 4500 9550 4720 9610
rect 4500 9510 4510 9550
rect 4550 9510 4590 9550
rect 4630 9510 4670 9550
rect 4710 9510 4720 9550
rect 4500 9450 4720 9510
rect 4500 9410 4510 9450
rect 4550 9410 4590 9450
rect 4630 9410 4670 9450
rect 4710 9410 4720 9450
rect 4500 9350 4720 9410
rect 4500 9310 4510 9350
rect 4550 9310 4590 9350
rect 4630 9310 4670 9350
rect 4710 9310 4720 9350
rect 4500 9250 4720 9310
rect 4500 9210 4510 9250
rect 4550 9210 4590 9250
rect 4630 9210 4670 9250
rect 4710 9210 4720 9250
rect 4500 9190 4720 9210
rect 5740 9650 5800 9670
rect 5740 9610 5750 9650
rect 5790 9610 5800 9650
rect 5740 9550 5800 9610
rect 5740 9510 5750 9550
rect 5790 9510 5800 9550
rect 5740 9450 5800 9510
rect 5740 9410 5750 9450
rect 5790 9410 5800 9450
rect 5740 9350 5800 9410
rect 11670 9400 11710 9750
rect 11750 9730 11850 9750
rect 5740 9310 5750 9350
rect 5790 9310 5800 9350
rect 5740 9250 5800 9310
rect 5740 9210 5750 9250
rect 5790 9210 5800 9250
rect 5740 9190 5800 9210
rect 3420 9120 3430 9160
rect 3470 9120 3480 9160
rect 3420 9100 3480 9120
rect 3710 9130 3790 9150
rect 2750 9070 2830 9090
rect 3710 9090 3730 9130
rect 3770 9090 3790 9130
rect 3710 9070 3790 9090
rect 3950 9130 4030 9150
rect 3950 9090 3970 9130
rect 4010 9090 4030 9130
rect 3950 9070 4030 9090
rect 4190 9130 4270 9150
rect 4190 9090 4210 9130
rect 4250 9090 4270 9130
rect 4190 9070 4270 9090
rect 4830 9130 4910 9150
rect 4830 9090 4850 9130
rect 4890 9090 4910 9130
rect 4830 9070 4910 9090
rect 5070 9130 5150 9150
rect 5070 9090 5090 9130
rect 5130 9090 5150 9130
rect 5070 9070 5150 9090
rect 5310 9130 5390 9150
rect 5310 9090 5330 9130
rect 5370 9090 5390 9130
rect 5310 9070 5390 9090
rect 5550 9130 5630 9150
rect 5550 9090 5570 9130
rect 5610 9090 5630 9130
rect 5550 9070 5630 9090
rect 7856 8870 7890 8886
rect 7650 8836 7856 8870
rect 7650 8830 7890 8836
rect 1421 8752 1479 8770
rect 1421 8718 1433 8752
rect 1467 8718 1479 8752
rect 1421 8700 1479 8718
rect 1781 8752 1839 8770
rect 1781 8718 1793 8752
rect 1827 8718 1839 8752
rect 1781 8700 1839 8718
rect 1901 8752 1959 8770
rect 1901 8718 1913 8752
rect 1947 8718 1959 8752
rect 1901 8700 1959 8718
rect 2261 8752 2319 8770
rect 2261 8718 2273 8752
rect 2307 8718 2319 8752
rect 2261 8700 2319 8718
rect 2381 8752 2439 8770
rect 2381 8718 2393 8752
rect 2427 8718 2439 8752
rect 4101 8752 4159 8770
rect 2381 8700 2439 8718
rect 2790 8730 2870 8750
rect 2790 8690 2810 8730
rect 2850 8690 2870 8730
rect 1360 8640 1420 8660
rect 1360 8600 1370 8640
rect 1410 8600 1420 8640
rect 1360 8580 1420 8600
rect 1480 8640 1540 8660
rect 1480 8600 1490 8640
rect 1530 8600 1540 8640
rect 1480 8580 1540 8600
rect 1600 8640 1660 8660
rect 1600 8600 1610 8640
rect 1650 8600 1660 8640
rect 1600 8580 1660 8600
rect 1720 8640 1780 8660
rect 1720 8600 1730 8640
rect 1770 8600 1780 8640
rect 1720 8580 1780 8600
rect 1840 8640 1900 8660
rect 1840 8600 1850 8640
rect 1890 8600 1900 8640
rect 1840 8580 1900 8600
rect 1960 8640 2020 8660
rect 1960 8600 1970 8640
rect 2010 8600 2020 8640
rect 1960 8580 2020 8600
rect 2080 8640 2140 8660
rect 2080 8600 2090 8640
rect 2130 8600 2140 8640
rect 2080 8580 2140 8600
rect 2200 8640 2260 8660
rect 2200 8600 2210 8640
rect 2250 8600 2260 8640
rect 2200 8580 2260 8600
rect 2320 8640 2380 8660
rect 2320 8600 2330 8640
rect 2370 8600 2380 8640
rect 2320 8580 2380 8600
rect 2440 8640 2500 8660
rect 2440 8600 2450 8640
rect 2490 8600 2500 8640
rect 2440 8580 2500 8600
rect 2560 8640 2620 8660
rect 2560 8600 2570 8640
rect 2610 8600 2620 8640
rect 2560 8580 2620 8600
rect 2790 8650 2870 8690
rect 2790 8610 2810 8650
rect 2850 8610 2870 8650
rect 2790 8570 2870 8610
rect 1522 8522 1580 8540
rect 1522 8488 1534 8522
rect 1568 8488 1580 8522
rect 1522 8470 1580 8488
rect 1680 8522 1738 8540
rect 1680 8488 1692 8522
rect 1726 8488 1738 8522
rect 1680 8470 1738 8488
rect 2004 8522 2062 8540
rect 2004 8488 2016 8522
rect 2050 8488 2062 8522
rect 2004 8470 2062 8488
rect 2158 8522 2216 8540
rect 2158 8488 2170 8522
rect 2204 8488 2216 8522
rect 2158 8470 2216 8488
rect 2482 8522 2540 8540
rect 2482 8488 2494 8522
rect 2528 8488 2540 8522
rect 2790 8530 2810 8570
rect 2850 8530 2870 8570
rect 2790 8510 2870 8530
rect 3670 8730 3750 8750
rect 3670 8690 3690 8730
rect 3730 8690 3750 8730
rect 4101 8718 4113 8752
rect 4147 8718 4159 8752
rect 4101 8700 4159 8718
rect 4221 8752 4279 8770
rect 4221 8718 4233 8752
rect 4267 8718 4279 8752
rect 4221 8700 4279 8718
rect 4581 8752 4639 8770
rect 4581 8718 4593 8752
rect 4627 8718 4639 8752
rect 4581 8700 4639 8718
rect 4701 8752 4759 8770
rect 4701 8718 4713 8752
rect 4747 8718 4759 8752
rect 4701 8700 4759 8718
rect 5061 8752 5119 8770
rect 5061 8718 5073 8752
rect 5107 8718 5119 8752
rect 5061 8700 5119 8718
rect 3670 8650 3750 8690
rect 3670 8610 3690 8650
rect 3730 8610 3750 8650
rect 3670 8570 3750 8610
rect 3920 8640 3980 8660
rect 3920 8600 3930 8640
rect 3970 8600 3980 8640
rect 3920 8580 3980 8600
rect 4040 8640 4100 8660
rect 4040 8600 4050 8640
rect 4090 8600 4100 8640
rect 4040 8580 4100 8600
rect 4160 8640 4220 8660
rect 4160 8600 4170 8640
rect 4210 8600 4220 8640
rect 4160 8580 4220 8600
rect 4280 8640 4340 8660
rect 4280 8600 4290 8640
rect 4330 8600 4340 8640
rect 4280 8580 4340 8600
rect 4400 8640 4460 8660
rect 4400 8600 4410 8640
rect 4450 8600 4460 8640
rect 4400 8580 4460 8600
rect 4520 8640 4580 8660
rect 4520 8600 4530 8640
rect 4570 8600 4580 8640
rect 4520 8580 4580 8600
rect 4640 8640 4700 8660
rect 4640 8600 4650 8640
rect 4690 8600 4700 8640
rect 4640 8580 4700 8600
rect 4760 8640 4820 8660
rect 4760 8600 4770 8640
rect 4810 8600 4820 8640
rect 4760 8580 4820 8600
rect 4880 8640 4940 8660
rect 4880 8600 4890 8640
rect 4930 8600 4940 8640
rect 4880 8580 4940 8600
rect 5000 8640 5060 8660
rect 5000 8600 5010 8640
rect 5050 8600 5060 8640
rect 5000 8580 5060 8600
rect 5120 8640 5180 8660
rect 5120 8600 5130 8640
rect 5170 8600 5180 8640
rect 5120 8580 5180 8600
rect 3670 8530 3690 8570
rect 3730 8530 3750 8570
rect 3670 8510 3750 8530
rect 4000 8522 4058 8540
rect 2482 8470 2540 8488
rect 4000 8488 4012 8522
rect 4046 8488 4058 8522
rect 4000 8470 4058 8488
rect 4324 8522 4382 8540
rect 4324 8488 4336 8522
rect 4370 8488 4382 8522
rect 4324 8470 4382 8488
rect 4478 8522 4536 8540
rect 4478 8488 4490 8522
rect 4524 8488 4536 8522
rect 4478 8470 4536 8488
rect 4802 8522 4860 8540
rect 4802 8488 4814 8522
rect 4848 8488 4860 8522
rect 4802 8470 4860 8488
rect 4960 8522 5018 8540
rect 4960 8488 4972 8522
rect 5006 8488 5018 8522
rect 4960 8470 5018 8488
rect 700 7930 760 7950
rect 700 7890 710 7930
rect 750 7890 760 7930
rect 700 7870 760 7890
rect 870 7920 950 7940
rect 870 7880 890 7920
rect 930 7880 950 7920
rect 870 7860 950 7880
rect 1360 7920 1420 7940
rect 1360 7880 1370 7920
rect 1410 7880 1420 7920
rect 1360 7860 1420 7880
rect 1590 7920 1670 7940
rect 1590 7880 1610 7920
rect 1650 7880 1670 7920
rect 1590 7860 1670 7880
rect 2080 7920 2140 7940
rect 2080 7880 2090 7920
rect 2130 7880 2140 7920
rect 2080 7860 2140 7880
rect 2310 7920 2390 7940
rect 2310 7880 2330 7920
rect 2370 7880 2390 7920
rect 2310 7860 2390 7880
rect 2740 7920 2800 7940
rect 2740 7880 2750 7920
rect 2790 7880 2800 7920
rect 2740 7860 2800 7880
rect 3740 7920 3800 7940
rect 3740 7880 3750 7920
rect 3790 7880 3800 7920
rect 3740 7860 3800 7880
rect 4150 7920 4230 7940
rect 4150 7880 4170 7920
rect 4210 7880 4230 7920
rect 4150 7860 4230 7880
rect 4400 7920 4460 7940
rect 4400 7880 4410 7920
rect 4450 7880 4460 7920
rect 4400 7860 4460 7880
rect 4870 7920 4950 7940
rect 4870 7880 4890 7920
rect 4930 7880 4950 7920
rect 4870 7860 4950 7880
rect 5120 7920 5180 7940
rect 5120 7880 5130 7920
rect 5170 7880 5180 7920
rect 5120 7860 5180 7880
rect 5590 7920 5670 7940
rect 5590 7880 5610 7920
rect 5650 7880 5670 7920
rect 5590 7860 5670 7880
rect 5780 7930 5840 7950
rect 5780 7890 5790 7930
rect 5830 7890 5840 7930
rect 5780 7870 5840 7890
rect 440 7800 580 7820
rect 440 7760 450 7800
rect 490 7760 530 7800
rect 570 7760 580 7800
rect 440 7700 580 7760
rect 440 7660 450 7700
rect 490 7660 530 7700
rect 570 7660 580 7700
rect 440 7640 580 7660
rect 640 7800 700 7820
rect 640 7760 650 7800
rect 690 7760 700 7800
rect 640 7700 700 7760
rect 640 7660 650 7700
rect 690 7660 700 7700
rect 640 7640 700 7660
rect 760 7800 820 7820
rect 760 7760 770 7800
rect 810 7760 820 7800
rect 760 7700 820 7760
rect 760 7660 770 7700
rect 810 7660 820 7700
rect 760 7640 820 7660
rect 880 7800 940 7820
rect 880 7760 890 7800
rect 930 7760 940 7800
rect 880 7700 940 7760
rect 880 7660 890 7700
rect 930 7660 940 7700
rect 880 7640 940 7660
rect 1000 7800 1060 7820
rect 1000 7760 1010 7800
rect 1050 7760 1060 7800
rect 1000 7700 1060 7760
rect 1000 7660 1010 7700
rect 1050 7660 1060 7700
rect 1000 7640 1060 7660
rect 1120 7800 1180 7820
rect 1120 7760 1130 7800
rect 1170 7760 1180 7800
rect 1120 7700 1180 7760
rect 1120 7660 1130 7700
rect 1170 7660 1180 7700
rect 1120 7640 1180 7660
rect 1240 7800 1300 7820
rect 1240 7760 1250 7800
rect 1290 7760 1300 7800
rect 1240 7700 1300 7760
rect 1240 7660 1250 7700
rect 1290 7660 1300 7700
rect 1240 7640 1300 7660
rect 1360 7800 1420 7820
rect 1360 7760 1370 7800
rect 1410 7760 1420 7800
rect 1360 7700 1420 7760
rect 1360 7660 1370 7700
rect 1410 7660 1420 7700
rect 1360 7640 1420 7660
rect 1480 7800 1540 7820
rect 1480 7760 1490 7800
rect 1530 7760 1540 7800
rect 1480 7700 1540 7760
rect 1480 7660 1490 7700
rect 1530 7660 1540 7700
rect 1480 7640 1540 7660
rect 1600 7800 1660 7820
rect 1600 7760 1610 7800
rect 1650 7760 1660 7800
rect 1600 7700 1660 7760
rect 1600 7660 1610 7700
rect 1650 7660 1660 7700
rect 1600 7640 1660 7660
rect 1720 7800 1780 7820
rect 1720 7760 1730 7800
rect 1770 7760 1780 7800
rect 1720 7700 1780 7760
rect 1720 7660 1730 7700
rect 1770 7660 1780 7700
rect 1720 7640 1780 7660
rect 1840 7800 1900 7820
rect 1840 7760 1850 7800
rect 1890 7760 1900 7800
rect 1840 7700 1900 7760
rect 1840 7660 1850 7700
rect 1890 7660 1900 7700
rect 1840 7640 1900 7660
rect 1960 7800 2020 7820
rect 1960 7760 1970 7800
rect 2010 7760 2020 7800
rect 1960 7700 2020 7760
rect 1960 7660 1970 7700
rect 2010 7660 2020 7700
rect 1960 7640 2020 7660
rect 2080 7800 2140 7820
rect 2080 7760 2090 7800
rect 2130 7760 2140 7800
rect 2080 7700 2140 7760
rect 2080 7660 2090 7700
rect 2130 7660 2140 7700
rect 2080 7640 2140 7660
rect 2200 7800 2260 7820
rect 2200 7760 2210 7800
rect 2250 7760 2260 7800
rect 2200 7700 2260 7760
rect 2200 7660 2210 7700
rect 2250 7660 2260 7700
rect 2200 7640 2260 7660
rect 2320 7800 2380 7820
rect 2320 7760 2330 7800
rect 2370 7760 2380 7800
rect 2320 7700 2380 7760
rect 2320 7660 2330 7700
rect 2370 7660 2380 7700
rect 2320 7640 2380 7660
rect 2440 7800 2500 7820
rect 2440 7760 2450 7800
rect 2490 7760 2500 7800
rect 2440 7700 2500 7760
rect 2440 7660 2450 7700
rect 2490 7660 2500 7700
rect 2440 7640 2500 7660
rect 2560 7800 2620 7820
rect 2560 7760 2570 7800
rect 2610 7760 2620 7800
rect 2560 7700 2620 7760
rect 2560 7660 2570 7700
rect 2610 7660 2620 7700
rect 2560 7640 2620 7660
rect 2680 7800 2740 7820
rect 2680 7760 2690 7800
rect 2730 7760 2740 7800
rect 2680 7700 2740 7760
rect 2680 7660 2690 7700
rect 2730 7660 2740 7700
rect 2680 7640 2740 7660
rect 2800 7800 2860 7820
rect 2800 7760 2810 7800
rect 2850 7760 2860 7800
rect 2800 7700 2860 7760
rect 2800 7660 2810 7700
rect 2850 7660 2860 7700
rect 2800 7640 2860 7660
rect 2920 7800 3060 7820
rect 2920 7760 2930 7800
rect 2970 7760 3010 7800
rect 3050 7760 3060 7800
rect 2920 7700 3060 7760
rect 2920 7660 2930 7700
rect 2970 7660 3010 7700
rect 3050 7660 3060 7700
rect 2920 7640 3060 7660
rect 3480 7800 3620 7820
rect 3480 7760 3490 7800
rect 3530 7760 3570 7800
rect 3610 7760 3620 7800
rect 3480 7700 3620 7760
rect 3480 7660 3490 7700
rect 3530 7660 3570 7700
rect 3610 7660 3620 7700
rect 3480 7640 3620 7660
rect 3680 7800 3740 7820
rect 3680 7760 3690 7800
rect 3730 7760 3740 7800
rect 3680 7700 3740 7760
rect 3680 7660 3690 7700
rect 3730 7660 3740 7700
rect 3680 7640 3740 7660
rect 3800 7800 3860 7820
rect 3800 7760 3810 7800
rect 3850 7760 3860 7800
rect 3800 7700 3860 7760
rect 3800 7660 3810 7700
rect 3850 7660 3860 7700
rect 3800 7640 3860 7660
rect 3920 7800 3980 7820
rect 3920 7760 3930 7800
rect 3970 7760 3980 7800
rect 3920 7700 3980 7760
rect 3920 7660 3930 7700
rect 3970 7660 3980 7700
rect 3920 7640 3980 7660
rect 4040 7800 4100 7820
rect 4040 7760 4050 7800
rect 4090 7760 4100 7800
rect 4040 7700 4100 7760
rect 4040 7660 4050 7700
rect 4090 7660 4100 7700
rect 4040 7640 4100 7660
rect 4160 7800 4220 7820
rect 4160 7760 4170 7800
rect 4210 7760 4220 7800
rect 4160 7700 4220 7760
rect 4160 7660 4170 7700
rect 4210 7660 4220 7700
rect 4160 7640 4220 7660
rect 4280 7800 4340 7820
rect 4280 7760 4290 7800
rect 4330 7760 4340 7800
rect 4280 7700 4340 7760
rect 4280 7660 4290 7700
rect 4330 7660 4340 7700
rect 4280 7640 4340 7660
rect 4400 7800 4460 7820
rect 4400 7760 4410 7800
rect 4450 7760 4460 7800
rect 4400 7700 4460 7760
rect 4400 7660 4410 7700
rect 4450 7660 4460 7700
rect 4400 7640 4460 7660
rect 4520 7800 4580 7820
rect 4520 7760 4530 7800
rect 4570 7760 4580 7800
rect 4520 7700 4580 7760
rect 4520 7660 4530 7700
rect 4570 7660 4580 7700
rect 4520 7640 4580 7660
rect 4640 7800 4700 7820
rect 4640 7760 4650 7800
rect 4690 7760 4700 7800
rect 4640 7700 4700 7760
rect 4640 7660 4650 7700
rect 4690 7660 4700 7700
rect 4640 7640 4700 7660
rect 4760 7800 4820 7820
rect 4760 7760 4770 7800
rect 4810 7760 4820 7800
rect 4760 7700 4820 7760
rect 4760 7660 4770 7700
rect 4810 7660 4820 7700
rect 4760 7640 4820 7660
rect 4880 7800 4940 7820
rect 4880 7760 4890 7800
rect 4930 7760 4940 7800
rect 4880 7700 4940 7760
rect 4880 7660 4890 7700
rect 4930 7660 4940 7700
rect 4880 7640 4940 7660
rect 5000 7800 5060 7820
rect 5000 7760 5010 7800
rect 5050 7760 5060 7800
rect 5000 7700 5060 7760
rect 5000 7660 5010 7700
rect 5050 7660 5060 7700
rect 5000 7640 5060 7660
rect 5120 7800 5180 7820
rect 5120 7760 5130 7800
rect 5170 7760 5180 7800
rect 5120 7700 5180 7760
rect 5120 7660 5130 7700
rect 5170 7660 5180 7700
rect 5120 7640 5180 7660
rect 5240 7800 5300 7820
rect 5240 7760 5250 7800
rect 5290 7760 5300 7800
rect 5240 7700 5300 7760
rect 5240 7660 5250 7700
rect 5290 7660 5300 7700
rect 5240 7640 5300 7660
rect 5360 7800 5420 7820
rect 5360 7760 5370 7800
rect 5410 7760 5420 7800
rect 5360 7700 5420 7760
rect 5360 7660 5370 7700
rect 5410 7660 5420 7700
rect 5360 7640 5420 7660
rect 5480 7800 5540 7820
rect 5480 7760 5490 7800
rect 5530 7760 5540 7800
rect 5480 7700 5540 7760
rect 5480 7660 5490 7700
rect 5530 7660 5540 7700
rect 5480 7640 5540 7660
rect 5600 7800 5660 7820
rect 5600 7760 5610 7800
rect 5650 7760 5660 7800
rect 5600 7700 5660 7760
rect 5600 7660 5610 7700
rect 5650 7660 5660 7700
rect 5600 7640 5660 7660
rect 5720 7800 5780 7820
rect 5720 7760 5730 7800
rect 5770 7760 5780 7800
rect 5720 7700 5780 7760
rect 5720 7660 5730 7700
rect 5770 7660 5780 7700
rect 5720 7640 5780 7660
rect 5840 7800 5900 7820
rect 5840 7760 5850 7800
rect 5890 7760 5900 7800
rect 5840 7700 5900 7760
rect 5840 7660 5850 7700
rect 5890 7660 5900 7700
rect 5840 7640 5900 7660
rect 5960 7800 6100 7820
rect 5960 7760 5970 7800
rect 6010 7760 6050 7800
rect 6090 7760 6100 7800
rect 5960 7700 6100 7760
rect 5960 7660 5970 7700
rect 6010 7660 6050 7700
rect 6090 7660 6100 7700
rect 5960 7640 6100 7660
rect 520 7580 580 7600
rect 520 7540 530 7580
rect 570 7540 580 7580
rect 520 7520 580 7540
rect 2920 7580 2980 7600
rect 2920 7540 2930 7580
rect 2970 7540 2980 7580
rect 2920 7520 2980 7540
rect 3560 7580 3620 7600
rect 3560 7540 3570 7580
rect 3610 7540 3620 7580
rect 3560 7520 3620 7540
rect 5960 7580 6020 7600
rect 5960 7540 5970 7580
rect 6010 7540 6020 7580
rect 5960 7520 6020 7540
rect 1890 6760 1960 6780
rect 1890 6720 1900 6760
rect 1940 6720 1960 6760
rect 1890 6700 1960 6720
rect 2060 6760 2140 6780
rect 2060 6720 2080 6760
rect 2120 6720 2140 6760
rect 2060 6700 2140 6720
rect 2240 6760 2320 6780
rect 2240 6720 2260 6760
rect 2300 6720 2320 6760
rect 2240 6700 2320 6720
rect 2420 6760 2500 6780
rect 2420 6720 2440 6760
rect 2480 6720 2500 6760
rect 2420 6700 2500 6720
rect 2600 6760 2680 6780
rect 2600 6720 2620 6760
rect 2660 6720 2680 6760
rect 2600 6700 2680 6720
rect 2780 6760 2860 6780
rect 2780 6720 2800 6760
rect 2840 6720 2860 6760
rect 2780 6700 2860 6720
rect 2960 6760 3040 6780
rect 2960 6720 2980 6760
rect 3020 6720 3040 6760
rect 2960 6700 3040 6720
rect 3140 6760 3210 6780
rect 3140 6720 3160 6760
rect 3200 6720 3210 6760
rect 3140 6700 3210 6720
rect 3330 6760 3400 6780
rect 3330 6720 3340 6760
rect 3380 6720 3400 6760
rect 3330 6700 3400 6720
rect 3500 6760 3580 6780
rect 3500 6720 3520 6760
rect 3560 6720 3580 6760
rect 3500 6700 3580 6720
rect 3680 6760 3760 6780
rect 3680 6720 3700 6760
rect 3740 6720 3760 6760
rect 3680 6700 3760 6720
rect 3860 6760 3940 6780
rect 3860 6720 3880 6760
rect 3920 6720 3940 6760
rect 3860 6700 3940 6720
rect 4040 6760 4120 6780
rect 4040 6720 4060 6760
rect 4100 6720 4120 6760
rect 4040 6700 4120 6720
rect 4220 6760 4300 6780
rect 4220 6720 4240 6760
rect 4280 6720 4300 6760
rect 4220 6700 4300 6720
rect 4400 6760 4480 6780
rect 4400 6720 4420 6760
rect 4460 6720 4480 6760
rect 4400 6700 4480 6720
rect 4580 6760 4650 6780
rect 4580 6720 4600 6760
rect 4640 6720 4650 6760
rect 4580 6700 4650 6720
rect 1540 6640 1680 6660
rect 1540 6600 1550 6640
rect 1590 6600 1630 6640
rect 1670 6600 1680 6640
rect 1540 6540 1680 6600
rect 1540 6500 1550 6540
rect 1590 6500 1630 6540
rect 1670 6500 1680 6540
rect 1540 6440 1680 6500
rect 1540 6400 1550 6440
rect 1590 6400 1630 6440
rect 1670 6400 1680 6440
rect 1540 6340 1680 6400
rect 1540 6300 1550 6340
rect 1590 6300 1630 6340
rect 1670 6300 1680 6340
rect 1540 6240 1680 6300
rect 1540 6200 1550 6240
rect 1590 6200 1630 6240
rect 1670 6200 1680 6240
rect 1540 6140 1680 6200
rect 1540 6100 1550 6140
rect 1590 6100 1630 6140
rect 1670 6100 1680 6140
rect 1540 6080 1680 6100
rect 1800 6640 1860 6660
rect 1800 6600 1810 6640
rect 1850 6600 1860 6640
rect 1800 6540 1860 6600
rect 1800 6500 1810 6540
rect 1850 6500 1860 6540
rect 1800 6440 1860 6500
rect 1800 6400 1810 6440
rect 1850 6400 1860 6440
rect 1800 6340 1860 6400
rect 1800 6300 1810 6340
rect 1850 6300 1860 6340
rect 1800 6240 1860 6300
rect 1800 6200 1810 6240
rect 1850 6200 1860 6240
rect 1800 6140 1860 6200
rect 1800 6100 1810 6140
rect 1850 6100 1860 6140
rect 1800 6080 1860 6100
rect 1980 6640 2040 6660
rect 1980 6600 1990 6640
rect 2030 6600 2040 6640
rect 1980 6540 2040 6600
rect 1980 6500 1990 6540
rect 2030 6500 2040 6540
rect 1980 6440 2040 6500
rect 1980 6400 1990 6440
rect 2030 6400 2040 6440
rect 1980 6340 2040 6400
rect 1980 6300 1990 6340
rect 2030 6300 2040 6340
rect 1980 6240 2040 6300
rect 1980 6200 1990 6240
rect 2030 6200 2040 6240
rect 1980 6140 2040 6200
rect 1980 6100 1990 6140
rect 2030 6100 2040 6140
rect 1980 6080 2040 6100
rect 2160 6640 2220 6660
rect 2160 6600 2170 6640
rect 2210 6600 2220 6640
rect 2160 6540 2220 6600
rect 2160 6500 2170 6540
rect 2210 6500 2220 6540
rect 2160 6440 2220 6500
rect 2160 6400 2170 6440
rect 2210 6400 2220 6440
rect 2160 6340 2220 6400
rect 2160 6300 2170 6340
rect 2210 6300 2220 6340
rect 2160 6240 2220 6300
rect 2160 6200 2170 6240
rect 2210 6200 2220 6240
rect 2160 6140 2220 6200
rect 2160 6100 2170 6140
rect 2210 6100 2220 6140
rect 2160 6080 2220 6100
rect 2340 6640 2400 6660
rect 2340 6600 2350 6640
rect 2390 6600 2400 6640
rect 2340 6540 2400 6600
rect 2340 6500 2350 6540
rect 2390 6500 2400 6540
rect 2340 6440 2400 6500
rect 2340 6400 2350 6440
rect 2390 6400 2400 6440
rect 2340 6340 2400 6400
rect 2340 6300 2350 6340
rect 2390 6300 2400 6340
rect 2340 6240 2400 6300
rect 2340 6200 2350 6240
rect 2390 6200 2400 6240
rect 2340 6140 2400 6200
rect 2340 6100 2350 6140
rect 2390 6100 2400 6140
rect 2340 6080 2400 6100
rect 2520 6640 2580 6660
rect 2520 6600 2530 6640
rect 2570 6600 2580 6640
rect 2520 6540 2580 6600
rect 2520 6500 2530 6540
rect 2570 6500 2580 6540
rect 2520 6440 2580 6500
rect 2520 6400 2530 6440
rect 2570 6400 2580 6440
rect 2520 6340 2580 6400
rect 2520 6300 2530 6340
rect 2570 6300 2580 6340
rect 2520 6240 2580 6300
rect 2520 6200 2530 6240
rect 2570 6200 2580 6240
rect 2520 6140 2580 6200
rect 2520 6100 2530 6140
rect 2570 6100 2580 6140
rect 2520 6080 2580 6100
rect 2700 6640 2760 6660
rect 2700 6600 2710 6640
rect 2750 6600 2760 6640
rect 2700 6540 2760 6600
rect 2700 6500 2710 6540
rect 2750 6500 2760 6540
rect 2700 6440 2760 6500
rect 2700 6400 2710 6440
rect 2750 6400 2760 6440
rect 2700 6340 2760 6400
rect 2700 6300 2710 6340
rect 2750 6300 2760 6340
rect 2700 6240 2760 6300
rect 2700 6200 2710 6240
rect 2750 6200 2760 6240
rect 2700 6140 2760 6200
rect 2700 6100 2710 6140
rect 2750 6100 2760 6140
rect 2700 6080 2760 6100
rect 2880 6640 2940 6660
rect 2880 6600 2890 6640
rect 2930 6600 2940 6640
rect 2880 6540 2940 6600
rect 2880 6500 2890 6540
rect 2930 6500 2940 6540
rect 2880 6440 2940 6500
rect 2880 6400 2890 6440
rect 2930 6400 2940 6440
rect 2880 6340 2940 6400
rect 2880 6300 2890 6340
rect 2930 6300 2940 6340
rect 2880 6240 2940 6300
rect 2880 6200 2890 6240
rect 2930 6200 2940 6240
rect 2880 6140 2940 6200
rect 2880 6100 2890 6140
rect 2930 6100 2940 6140
rect 2880 6080 2940 6100
rect 3060 6640 3120 6660
rect 3060 6600 3070 6640
rect 3110 6600 3120 6640
rect 3060 6540 3120 6600
rect 3060 6500 3070 6540
rect 3110 6500 3120 6540
rect 3060 6440 3120 6500
rect 3060 6400 3070 6440
rect 3110 6400 3120 6440
rect 3060 6340 3120 6400
rect 3060 6300 3070 6340
rect 3110 6300 3120 6340
rect 3060 6240 3120 6300
rect 3060 6200 3070 6240
rect 3110 6200 3120 6240
rect 3060 6140 3120 6200
rect 3060 6100 3070 6140
rect 3110 6100 3120 6140
rect 3060 6080 3120 6100
rect 3240 6640 3300 6660
rect 3240 6600 3250 6640
rect 3290 6600 3300 6640
rect 3240 6540 3300 6600
rect 3240 6500 3250 6540
rect 3290 6500 3300 6540
rect 3240 6440 3300 6500
rect 3240 6400 3250 6440
rect 3290 6400 3300 6440
rect 3240 6340 3300 6400
rect 3240 6300 3250 6340
rect 3290 6300 3300 6340
rect 3240 6240 3300 6300
rect 3240 6200 3250 6240
rect 3290 6200 3300 6240
rect 3240 6140 3300 6200
rect 3240 6100 3250 6140
rect 3290 6100 3300 6140
rect 3240 6080 3300 6100
rect 3420 6640 3480 6660
rect 3420 6600 3430 6640
rect 3470 6600 3480 6640
rect 3420 6540 3480 6600
rect 3420 6500 3430 6540
rect 3470 6500 3480 6540
rect 3420 6440 3480 6500
rect 3420 6400 3430 6440
rect 3470 6400 3480 6440
rect 3420 6340 3480 6400
rect 3420 6300 3430 6340
rect 3470 6300 3480 6340
rect 3420 6240 3480 6300
rect 3420 6200 3430 6240
rect 3470 6200 3480 6240
rect 3420 6140 3480 6200
rect 3420 6100 3430 6140
rect 3470 6100 3480 6140
rect 3420 6080 3480 6100
rect 3600 6640 3660 6660
rect 3600 6600 3610 6640
rect 3650 6600 3660 6640
rect 3600 6540 3660 6600
rect 3600 6500 3610 6540
rect 3650 6500 3660 6540
rect 3600 6440 3660 6500
rect 3600 6400 3610 6440
rect 3650 6400 3660 6440
rect 3600 6340 3660 6400
rect 3600 6300 3610 6340
rect 3650 6300 3660 6340
rect 3600 6240 3660 6300
rect 3600 6200 3610 6240
rect 3650 6200 3660 6240
rect 3600 6140 3660 6200
rect 3600 6100 3610 6140
rect 3650 6100 3660 6140
rect 3600 6080 3660 6100
rect 3780 6640 3840 6660
rect 3780 6600 3790 6640
rect 3830 6600 3840 6640
rect 3780 6540 3840 6600
rect 3780 6500 3790 6540
rect 3830 6500 3840 6540
rect 3780 6440 3840 6500
rect 3780 6400 3790 6440
rect 3830 6400 3840 6440
rect 3780 6340 3840 6400
rect 3780 6300 3790 6340
rect 3830 6300 3840 6340
rect 3780 6240 3840 6300
rect 3780 6200 3790 6240
rect 3830 6200 3840 6240
rect 3780 6140 3840 6200
rect 3780 6100 3790 6140
rect 3830 6100 3840 6140
rect 3780 6080 3840 6100
rect 3960 6640 4020 6660
rect 3960 6600 3970 6640
rect 4010 6600 4020 6640
rect 3960 6540 4020 6600
rect 3960 6500 3970 6540
rect 4010 6500 4020 6540
rect 3960 6440 4020 6500
rect 3960 6400 3970 6440
rect 4010 6400 4020 6440
rect 3960 6340 4020 6400
rect 3960 6300 3970 6340
rect 4010 6300 4020 6340
rect 3960 6240 4020 6300
rect 3960 6200 3970 6240
rect 4010 6200 4020 6240
rect 3960 6140 4020 6200
rect 3960 6100 3970 6140
rect 4010 6100 4020 6140
rect 3960 6080 4020 6100
rect 4140 6640 4200 6660
rect 4140 6600 4150 6640
rect 4190 6600 4200 6640
rect 4140 6540 4200 6600
rect 4140 6500 4150 6540
rect 4190 6500 4200 6540
rect 4140 6440 4200 6500
rect 4140 6400 4150 6440
rect 4190 6400 4200 6440
rect 4140 6340 4200 6400
rect 4140 6300 4150 6340
rect 4190 6300 4200 6340
rect 4140 6240 4200 6300
rect 4140 6200 4150 6240
rect 4190 6200 4200 6240
rect 4140 6140 4200 6200
rect 4140 6100 4150 6140
rect 4190 6100 4200 6140
rect 4140 6080 4200 6100
rect 4320 6640 4380 6660
rect 4320 6600 4330 6640
rect 4370 6600 4380 6640
rect 4320 6540 4380 6600
rect 4320 6500 4330 6540
rect 4370 6500 4380 6540
rect 4320 6440 4380 6500
rect 4320 6400 4330 6440
rect 4370 6400 4380 6440
rect 4320 6340 4380 6400
rect 4320 6300 4330 6340
rect 4370 6300 4380 6340
rect 4320 6240 4380 6300
rect 4320 6200 4330 6240
rect 4370 6200 4380 6240
rect 4320 6140 4380 6200
rect 4320 6100 4330 6140
rect 4370 6100 4380 6140
rect 4320 6080 4380 6100
rect 4500 6640 4560 6660
rect 4500 6600 4510 6640
rect 4550 6600 4560 6640
rect 4500 6540 4560 6600
rect 4500 6500 4510 6540
rect 4550 6500 4560 6540
rect 4500 6440 4560 6500
rect 4500 6400 4510 6440
rect 4550 6400 4560 6440
rect 4500 6340 4560 6400
rect 4500 6300 4510 6340
rect 4550 6300 4560 6340
rect 4500 6240 4560 6300
rect 4500 6200 4510 6240
rect 4550 6200 4560 6240
rect 4500 6140 4560 6200
rect 4500 6100 4510 6140
rect 4550 6100 4560 6140
rect 4500 6080 4560 6100
rect 4680 6640 4740 6660
rect 4680 6600 4690 6640
rect 4730 6600 4740 6640
rect 4680 6540 4740 6600
rect 4680 6500 4690 6540
rect 4730 6500 4740 6540
rect 4680 6440 4740 6500
rect 4680 6400 4690 6440
rect 4730 6400 4740 6440
rect 4680 6340 4740 6400
rect 4680 6300 4690 6340
rect 4730 6300 4740 6340
rect 4680 6240 4740 6300
rect 4680 6200 4690 6240
rect 4730 6200 4740 6240
rect 4680 6140 4740 6200
rect 4680 6100 4690 6140
rect 4730 6100 4740 6140
rect 4680 6080 4740 6100
rect 4860 6640 5000 6660
rect 4860 6600 4870 6640
rect 4910 6600 4950 6640
rect 4990 6600 5000 6640
rect 4860 6540 5000 6600
rect 4860 6500 4870 6540
rect 4910 6500 4950 6540
rect 4990 6500 5000 6540
rect 5580 6560 5660 6580
rect 5580 6520 5600 6560
rect 5640 6520 5660 6560
rect 5580 6500 5660 6520
rect 5700 6560 5780 6580
rect 5700 6520 5720 6560
rect 5760 6520 5780 6560
rect 5700 6500 5780 6520
rect 5820 6560 5900 6580
rect 5820 6520 5840 6560
rect 5880 6520 5900 6560
rect 5820 6500 5900 6520
rect 4860 6440 5000 6500
rect 4860 6400 4870 6440
rect 4910 6400 4950 6440
rect 4990 6400 5000 6440
rect 4860 6340 5000 6400
rect 4860 6300 4870 6340
rect 4910 6300 4950 6340
rect 4990 6300 5000 6340
rect 4860 6240 5000 6300
rect 5400 6440 5550 6460
rect 5400 6400 5410 6440
rect 5450 6400 5500 6440
rect 5540 6400 5550 6440
rect 5400 6340 5550 6400
rect 5400 6300 5410 6340
rect 5450 6300 5500 6340
rect 5540 6300 5550 6340
rect 5400 6280 5550 6300
rect 5600 6440 5660 6460
rect 5600 6400 5610 6440
rect 5650 6400 5660 6440
rect 5600 6340 5660 6400
rect 5600 6300 5610 6340
rect 5650 6300 5660 6340
rect 5600 6280 5660 6300
rect 5710 6440 5770 6460
rect 5710 6400 5720 6440
rect 5760 6400 5770 6440
rect 5710 6340 5770 6400
rect 5710 6300 5720 6340
rect 5760 6300 5770 6340
rect 5710 6280 5770 6300
rect 5820 6440 5880 6460
rect 5820 6400 5830 6440
rect 5870 6400 5880 6440
rect 5820 6340 5880 6400
rect 5820 6300 5830 6340
rect 5870 6300 5880 6340
rect 5820 6280 5880 6300
rect 5930 6440 6070 6460
rect 5930 6400 5940 6440
rect 5980 6400 6020 6440
rect 6060 6400 6070 6440
rect 5930 6340 6070 6400
rect 5930 6300 5940 6340
rect 5980 6300 6020 6340
rect 6060 6300 6070 6340
rect 5930 6280 6070 6300
rect 4860 6200 4870 6240
rect 4910 6200 4950 6240
rect 4990 6200 5000 6240
rect 4860 6140 5000 6200
rect 5480 6220 5560 6240
rect 5480 6180 5500 6220
rect 5540 6180 5560 6220
rect 5480 6160 5560 6180
rect 5700 6220 5780 6240
rect 5700 6180 5720 6220
rect 5760 6180 5780 6220
rect 5700 6160 5780 6180
rect 5930 6220 5990 6240
rect 5930 6180 5940 6220
rect 5980 6180 5990 6220
rect 5930 6160 5990 6180
rect 7650 6160 7690 8830
rect 7856 8820 7890 8830
rect 9130 8870 9164 8886
rect 9164 8836 9470 8870
rect 9130 8830 9470 8836
rect 9130 8820 9164 8830
rect 9430 8720 9470 8830
rect 9010 8700 9090 8720
rect 9010 8660 9030 8700
rect 9070 8680 9090 8700
rect 9410 8700 9490 8720
rect 9410 8680 9430 8700
rect 9070 8660 9430 8680
rect 9470 8660 9490 8700
rect 9010 8640 9490 8660
rect 9030 8600 9070 8640
rect 9430 8600 9470 8640
rect 8110 8580 8290 8600
rect 8110 8530 8130 8580
rect 8170 8530 8230 8580
rect 8270 8530 8290 8580
rect 8110 8440 8290 8530
rect 8110 8390 8130 8440
rect 8170 8390 8230 8440
rect 8270 8390 8290 8440
rect 8110 8370 8290 8390
rect 8410 8580 8490 8600
rect 8410 8530 8430 8580
rect 8470 8530 8490 8580
rect 8410 8440 8490 8530
rect 8410 8390 8430 8440
rect 8470 8390 8490 8440
rect 8410 8370 8490 8390
rect 8610 8580 8690 8600
rect 8610 8530 8630 8580
rect 8670 8530 8690 8580
rect 8610 8440 8690 8530
rect 8610 8390 8630 8440
rect 8670 8390 8690 8440
rect 8610 8370 8690 8390
rect 8810 8580 8890 8600
rect 8810 8530 8830 8580
rect 8870 8530 8890 8580
rect 8810 8440 8890 8530
rect 8810 8390 8830 8440
rect 8870 8390 8890 8440
rect 8810 8370 8890 8390
rect 9010 8580 9090 8600
rect 9010 8530 9030 8580
rect 9070 8530 9090 8580
rect 9010 8440 9090 8530
rect 9010 8390 9030 8440
rect 9070 8390 9090 8440
rect 9010 8370 9090 8390
rect 9210 8580 9290 8600
rect 9210 8530 9230 8580
rect 9270 8530 9290 8580
rect 9210 8440 9290 8530
rect 9210 8390 9230 8440
rect 9270 8390 9290 8440
rect 9210 8370 9290 8390
rect 9410 8580 9490 8600
rect 9410 8530 9430 8580
rect 9470 8530 9490 8580
rect 9410 8440 9490 8530
rect 9410 8390 9430 8440
rect 9470 8390 9490 8440
rect 9410 8370 9490 8390
rect 9610 8580 9690 8600
rect 9610 8530 9630 8580
rect 9670 8530 9690 8580
rect 9610 8440 9690 8530
rect 9610 8390 9630 8440
rect 9670 8390 9690 8440
rect 9610 8370 9690 8390
rect 9810 8580 9890 8600
rect 9810 8530 9830 8580
rect 9870 8530 9890 8580
rect 9810 8440 9890 8530
rect 9810 8390 9830 8440
rect 9870 8390 9890 8440
rect 9810 8370 9890 8390
rect 10010 8580 10090 8600
rect 10010 8530 10030 8580
rect 10070 8530 10090 8580
rect 10010 8440 10090 8530
rect 10010 8390 10030 8440
rect 10070 8390 10090 8440
rect 10010 8370 10090 8390
rect 10210 8580 10390 8600
rect 10210 8530 10230 8580
rect 10270 8530 10330 8580
rect 10370 8530 10390 8580
rect 10210 8440 10390 8530
rect 10210 8390 10230 8440
rect 10270 8390 10330 8440
rect 10370 8390 10390 8440
rect 10210 8370 10390 8390
rect 8230 8330 8270 8370
rect 8630 8330 8670 8370
rect 9830 8330 9870 8370
rect 10230 8330 10270 8370
rect 8210 8310 8290 8330
rect 8210 8270 8230 8310
rect 8270 8270 8290 8310
rect 8630 8290 9870 8330
rect 8210 8250 8290 8270
rect 9790 8270 9870 8290
rect 9790 8230 9810 8270
rect 9850 8230 9870 8270
rect 10210 8310 10290 8330
rect 10210 8270 10230 8310
rect 10270 8270 10290 8310
rect 10210 8250 10290 8270
rect 9790 8210 9870 8230
rect 7930 8120 7990 8160
rect 8030 8120 8090 8160
rect 8130 8120 8190 8160
rect 8230 8120 8290 8160
rect 8330 8120 8390 8160
rect 8430 8120 8490 8160
rect 8530 8120 8590 8160
rect 8630 8120 8690 8160
rect 8730 8120 8790 8160
rect 8830 8120 8890 8160
rect 8930 8120 8990 8160
rect 9030 8120 9090 8160
rect 9130 8120 9190 8160
rect 9230 8120 9290 8160
rect 9330 8120 9390 8160
rect 9430 8120 9490 8160
rect 9530 8120 9590 8160
rect 9630 8120 9690 8160
rect 9730 8120 9790 8160
rect 9830 8120 9890 8160
rect 9930 8120 9990 8160
rect 10030 8120 10090 8160
rect 10130 8120 10190 8160
rect 10230 8120 10290 8160
rect 10330 8120 10390 8160
rect 10430 8120 10490 8160
rect 10530 8120 10590 8160
rect 10630 8120 10690 8160
rect 10730 8120 10790 8160
rect 10830 8120 10890 8160
rect 10930 8120 10990 8160
rect 8320 8020 8410 8040
rect 8320 7990 8340 8020
rect 8280 7970 8340 7990
rect 8390 7990 8410 8020
rect 8670 7990 8710 8120
rect 9790 8050 9870 8070
rect 8970 8020 9060 8040
rect 8970 7990 8990 8020
rect 8390 7970 8990 7990
rect 9040 7990 9060 8020
rect 9460 8010 9540 8030
rect 9460 7990 9480 8010
rect 9040 7970 9100 7990
rect 8280 7950 9100 7970
rect 8280 7910 8320 7950
rect 8410 7910 8450 7950
rect 8670 7910 8710 7950
rect 8930 7910 8970 7950
rect 9060 7910 9100 7950
rect 9420 7970 9480 7990
rect 9520 7990 9540 8010
rect 9790 8010 9810 8050
rect 9850 8010 9870 8050
rect 9790 7990 9870 8010
rect 10120 8010 10200 8030
rect 10120 7990 10140 8010
rect 9520 7970 10140 7990
rect 10180 7990 10200 8010
rect 10600 8010 10680 8030
rect 10600 8000 10620 8010
rect 10180 7970 10240 7990
rect 9420 7950 10240 7970
rect 9420 7910 9460 7950
rect 9550 7910 9590 7950
rect 9810 7910 9850 7950
rect 10070 7910 10110 7950
rect 10200 7910 10240 7950
rect 10560 7970 10620 8000
rect 10660 8000 10680 8010
rect 10950 8000 10990 8120
rect 11260 8010 11340 8030
rect 11260 8000 11280 8010
rect 10660 7970 11280 8000
rect 11320 8000 11340 8010
rect 11320 7970 11380 8000
rect 10560 7950 11380 7970
rect 10560 7910 10600 7950
rect 10690 7910 10730 7950
rect 10950 7910 10990 7950
rect 11210 7910 11250 7950
rect 11340 7910 11380 7950
rect 8160 7890 8340 7910
rect 8160 7850 8180 7890
rect 8220 7850 8280 7890
rect 8320 7850 8340 7890
rect 8160 7830 8340 7850
rect 8390 7890 8470 7910
rect 8390 7850 8410 7890
rect 8450 7850 8470 7890
rect 8390 7830 8470 7850
rect 8520 7890 8600 7910
rect 8520 7850 8540 7890
rect 8580 7850 8600 7890
rect 8520 7830 8600 7850
rect 8650 7890 8730 7910
rect 8650 7850 8670 7890
rect 8710 7850 8730 7890
rect 8650 7830 8730 7850
rect 8780 7890 8860 7910
rect 8780 7850 8800 7890
rect 8840 7850 8860 7890
rect 8780 7830 8860 7850
rect 8910 7890 8990 7910
rect 8910 7850 8930 7890
rect 8970 7850 8990 7890
rect 8910 7830 8990 7850
rect 9040 7890 9220 7910
rect 9040 7850 9060 7890
rect 9100 7850 9160 7890
rect 9200 7850 9220 7890
rect 9040 7830 9220 7850
rect 9390 7890 9480 7910
rect 9390 7850 9420 7890
rect 9460 7850 9480 7890
rect 9390 7830 9480 7850
rect 9530 7890 9610 7910
rect 9530 7850 9550 7890
rect 9590 7850 9610 7890
rect 9530 7830 9610 7850
rect 9660 7890 9740 7910
rect 9660 7850 9680 7890
rect 9720 7850 9740 7890
rect 9660 7830 9740 7850
rect 9790 7890 9870 7910
rect 9790 7850 9810 7890
rect 9850 7850 9870 7890
rect 9790 7830 9870 7850
rect 9920 7890 10000 7910
rect 9920 7850 9940 7890
rect 9980 7850 10000 7890
rect 9920 7830 10000 7850
rect 10050 7890 10130 7910
rect 10050 7850 10070 7890
rect 10110 7850 10130 7890
rect 10050 7830 10130 7850
rect 10180 7890 10270 7910
rect 10180 7850 10200 7890
rect 10240 7850 10270 7890
rect 10180 7830 10270 7850
rect 10440 7890 10620 7910
rect 10440 7850 10460 7890
rect 10500 7850 10560 7890
rect 10600 7850 10620 7890
rect 10440 7830 10620 7850
rect 10670 7890 10750 7910
rect 10670 7850 10690 7890
rect 10730 7850 10750 7890
rect 10670 7830 10750 7850
rect 10800 7890 10880 7910
rect 10800 7850 10820 7890
rect 10860 7850 10880 7890
rect 10800 7830 10880 7850
rect 10930 7890 11010 7910
rect 10930 7850 10950 7890
rect 10990 7850 11010 7890
rect 10930 7830 11010 7850
rect 11060 7890 11140 7910
rect 11060 7850 11080 7890
rect 11120 7850 11140 7890
rect 11060 7830 11140 7850
rect 11190 7890 11270 7910
rect 11190 7850 11210 7890
rect 11250 7850 11270 7890
rect 11190 7830 11270 7850
rect 11320 7890 11500 7910
rect 11320 7850 11340 7890
rect 11380 7850 11440 7890
rect 11480 7850 11500 7890
rect 11320 7830 11500 7850
rect 8560 7790 8600 7830
rect 8520 7770 8600 7790
rect 8520 7730 8540 7770
rect 8580 7730 8600 7770
rect 8520 7710 8600 7730
rect 8430 7440 8510 7460
rect 8430 7400 8450 7440
rect 8490 7400 8510 7440
rect 8430 7380 8510 7400
rect 8560 7340 8600 7710
rect 8780 7620 8820 7830
rect 9570 7770 9650 7790
rect 9570 7730 9590 7770
rect 9630 7730 9650 7770
rect 9570 7710 9650 7730
rect 8780 7600 9410 7620
rect 8780 7580 9350 7600
rect 8780 7340 8820 7580
rect 9330 7560 9350 7580
rect 9390 7560 9410 7600
rect 9330 7550 9410 7560
rect 9700 7470 9740 7830
rect 8870 7440 8950 7460
rect 8870 7400 8890 7440
rect 8930 7400 8950 7440
rect 8870 7380 8950 7400
rect 9660 7450 9740 7470
rect 9660 7410 9680 7450
rect 9720 7410 9740 7450
rect 9660 7390 9740 7410
rect 9920 7440 9960 7830
rect 10010 7750 10090 7770
rect 10010 7710 10030 7750
rect 10070 7710 10090 7750
rect 10010 7690 10090 7710
rect 10840 7670 10880 7830
rect 11060 7670 11100 7830
rect 11550 7770 11630 7790
rect 11550 7730 11570 7770
rect 11610 7750 11630 7770
rect 11670 7750 11710 8380
rect 11610 7730 11710 7750
rect 11550 7710 11710 7730
rect 11750 7880 11860 7900
rect 11750 7810 11770 7880
rect 11840 7810 11860 7880
rect 11750 7790 11860 7810
rect 11750 7670 11790 7790
rect 10710 7650 10790 7670
rect 10710 7610 10730 7650
rect 10770 7610 10790 7650
rect 10840 7630 11960 7670
rect 10710 7590 10790 7610
rect 11920 7620 11960 7630
rect 11920 7600 12000 7620
rect 11920 7560 11940 7600
rect 11980 7560 12000 7600
rect 11920 7540 12000 7560
rect 10840 7500 11960 7540
rect 10710 7440 10790 7460
rect 9920 7400 10730 7440
rect 10770 7400 10790 7440
rect 9680 7340 9720 7390
rect 9920 7340 9960 7400
rect 10710 7380 10790 7400
rect 10840 7340 10880 7500
rect 11060 7340 11100 7500
rect 11550 7440 11710 7460
rect 11550 7400 11570 7440
rect 11610 7420 11710 7440
rect 11610 7400 11630 7420
rect 11550 7380 11630 7400
rect 8250 7320 8340 7340
rect 8250 7280 8280 7320
rect 8320 7280 8340 7320
rect 8250 7220 8340 7280
rect 8250 7180 8280 7220
rect 8320 7180 8340 7220
rect 8250 7160 8340 7180
rect 8390 7320 8470 7340
rect 8390 7280 8410 7320
rect 8450 7280 8470 7320
rect 8390 7220 8470 7280
rect 8390 7180 8410 7220
rect 8450 7180 8470 7220
rect 8390 7160 8470 7180
rect 8520 7320 8600 7340
rect 8520 7280 8540 7320
rect 8580 7280 8600 7320
rect 8520 7220 8600 7280
rect 8520 7180 8540 7220
rect 8580 7180 8600 7220
rect 8520 7160 8600 7180
rect 8650 7320 8730 7340
rect 8650 7280 8670 7320
rect 8710 7280 8730 7320
rect 8650 7220 8730 7280
rect 8650 7180 8670 7220
rect 8710 7180 8730 7220
rect 8650 7160 8730 7180
rect 8780 7320 8860 7340
rect 8780 7280 8800 7320
rect 8840 7280 8860 7320
rect 8780 7220 8860 7280
rect 8780 7180 8800 7220
rect 8840 7180 8860 7220
rect 8780 7160 8860 7180
rect 8910 7320 9000 7340
rect 8910 7280 8930 7320
rect 8970 7280 9000 7320
rect 8910 7220 9000 7280
rect 8910 7180 8930 7220
rect 8970 7180 9000 7220
rect 8910 7160 9000 7180
rect 9040 7320 9130 7340
rect 9040 7280 9060 7320
rect 9100 7280 9130 7320
rect 9040 7220 9130 7280
rect 9040 7180 9060 7220
rect 9100 7180 9130 7220
rect 9040 7160 9130 7180
rect 9300 7320 9480 7340
rect 9300 7280 9320 7320
rect 9360 7280 9420 7320
rect 9460 7280 9480 7320
rect 9300 7220 9480 7280
rect 9300 7180 9320 7220
rect 9360 7180 9420 7220
rect 9460 7180 9480 7220
rect 9300 7160 9480 7180
rect 9530 7320 9610 7340
rect 9530 7280 9550 7320
rect 9590 7280 9610 7320
rect 9530 7220 9610 7280
rect 9530 7180 9550 7220
rect 9590 7180 9610 7220
rect 9530 7160 9610 7180
rect 9660 7320 9740 7340
rect 9660 7280 9680 7320
rect 9720 7280 9740 7320
rect 9660 7220 9740 7280
rect 9660 7180 9680 7220
rect 9720 7180 9740 7220
rect 9660 7160 9740 7180
rect 9790 7320 9870 7340
rect 9790 7280 9810 7320
rect 9850 7280 9870 7320
rect 9790 7220 9870 7280
rect 9790 7180 9810 7220
rect 9850 7180 9870 7220
rect 9790 7160 9870 7180
rect 9920 7320 10000 7340
rect 9920 7280 9940 7320
rect 9980 7280 10000 7320
rect 9920 7220 10000 7280
rect 9920 7180 9940 7220
rect 9980 7180 10000 7220
rect 9920 7160 10000 7180
rect 10050 7320 10130 7340
rect 10050 7280 10070 7320
rect 10110 7280 10130 7320
rect 10050 7220 10130 7280
rect 10050 7180 10070 7220
rect 10110 7180 10130 7220
rect 10050 7160 10130 7180
rect 10180 7320 10360 7340
rect 10180 7280 10200 7320
rect 10240 7280 10300 7320
rect 10340 7280 10360 7320
rect 10180 7220 10360 7280
rect 10180 7180 10200 7220
rect 10240 7180 10300 7220
rect 10340 7180 10360 7220
rect 10180 7160 10360 7180
rect 10440 7320 10620 7340
rect 10440 7280 10460 7320
rect 10500 7280 10560 7320
rect 10600 7280 10620 7320
rect 10440 7220 10620 7280
rect 10440 7180 10460 7220
rect 10500 7180 10560 7220
rect 10600 7180 10620 7220
rect 10440 7160 10620 7180
rect 10670 7320 10750 7340
rect 10670 7280 10690 7320
rect 10730 7280 10750 7320
rect 10670 7220 10750 7280
rect 10670 7180 10690 7220
rect 10730 7180 10750 7220
rect 10670 7160 10750 7180
rect 10800 7320 10880 7340
rect 10800 7280 10820 7320
rect 10860 7280 10880 7320
rect 10800 7220 10880 7280
rect 10800 7180 10820 7220
rect 10860 7180 10880 7220
rect 10800 7160 10880 7180
rect 10930 7320 11010 7340
rect 10930 7280 10950 7320
rect 10990 7280 11010 7320
rect 10930 7220 11010 7280
rect 10930 7180 10950 7220
rect 10990 7180 11010 7220
rect 10930 7160 11010 7180
rect 11060 7320 11140 7340
rect 11060 7280 11080 7320
rect 11120 7280 11140 7320
rect 11060 7220 11140 7280
rect 11060 7180 11080 7220
rect 11120 7180 11140 7220
rect 11060 7160 11140 7180
rect 11190 7320 11270 7340
rect 11190 7280 11210 7320
rect 11250 7280 11270 7320
rect 11190 7220 11270 7280
rect 11190 7180 11210 7220
rect 11250 7180 11270 7220
rect 11190 7160 11270 7180
rect 11320 7320 11500 7340
rect 11320 7280 11340 7320
rect 11380 7280 11440 7320
rect 11480 7280 11500 7320
rect 11320 7220 11500 7280
rect 11320 7180 11340 7220
rect 11380 7180 11440 7220
rect 11480 7180 11500 7220
rect 11320 7160 11500 7180
rect 8280 7120 8320 7160
rect 8410 7120 8450 7160
rect 8670 7120 8710 7160
rect 8930 7120 8970 7160
rect 9060 7120 9100 7160
rect 8280 7100 9100 7120
rect 8280 7080 8340 7100
rect 8320 7060 8340 7080
rect 8380 7080 9000 7100
rect 8380 7060 8400 7080
rect 8320 7040 8400 7060
rect 8750 7060 8830 7080
rect 8750 7020 8770 7060
rect 8810 7020 8830 7060
rect 8980 7060 9000 7080
rect 9040 7080 9100 7100
rect 9420 7120 9460 7160
rect 9550 7120 9590 7160
rect 9810 7120 9850 7160
rect 10070 7120 10110 7160
rect 10200 7120 10240 7160
rect 9420 7100 10240 7120
rect 9420 7080 9480 7100
rect 9040 7060 9060 7080
rect 8980 7040 9060 7060
rect 9460 7060 9480 7080
rect 9520 7080 10140 7100
rect 9520 7060 9540 7080
rect 9460 7040 9540 7060
rect 8750 7000 8830 7020
rect 9810 6950 9850 7080
rect 10120 7060 10140 7080
rect 10180 7080 10240 7100
rect 10560 7120 10600 7160
rect 10690 7120 10730 7160
rect 10950 7120 10990 7160
rect 11210 7120 11250 7160
rect 11340 7120 11380 7160
rect 10560 7100 11380 7120
rect 11670 7110 11710 7420
rect 11750 7400 11790 7500
rect 11750 7380 11860 7400
rect 11750 7310 11770 7380
rect 11840 7310 11860 7380
rect 11750 7290 11860 7310
rect 10560 7080 10620 7100
rect 10180 7060 10200 7080
rect 10120 7040 10200 7060
rect 10600 7060 10620 7080
rect 10660 7080 11280 7100
rect 10660 7060 10680 7080
rect 10600 7040 10680 7060
rect 10950 6950 10990 7080
rect 11260 7060 11280 7080
rect 11320 7080 11380 7100
rect 11320 7060 11340 7080
rect 11260 7040 11340 7060
rect 7930 6910 7990 6950
rect 8030 6910 8090 6950
rect 8130 6910 8190 6950
rect 8230 6910 8290 6950
rect 8330 6910 8390 6950
rect 8430 6910 8490 6950
rect 8530 6910 8590 6950
rect 8630 6910 8690 6950
rect 8730 6910 8790 6950
rect 8830 6910 8890 6950
rect 8930 6910 8990 6950
rect 9030 6910 9090 6950
rect 9130 6910 9190 6950
rect 9230 6910 9290 6950
rect 9330 6910 9390 6950
rect 9430 6910 9490 6950
rect 9530 6910 9590 6950
rect 9630 6910 9690 6950
rect 9730 6910 9790 6950
rect 9830 6910 9890 6950
rect 9930 6910 9990 6950
rect 10030 6910 10090 6950
rect 10130 6910 10190 6950
rect 10230 6910 10290 6950
rect 10330 6910 10390 6950
rect 10430 6910 10490 6950
rect 10530 6910 10590 6950
rect 10630 6910 10690 6950
rect 10730 6910 10790 6950
rect 10830 6910 10890 6950
rect 10930 6910 10990 6950
rect 8750 6840 8830 6860
rect 8330 6790 8410 6810
rect 8330 6750 8350 6790
rect 8390 6750 8410 6790
rect 8330 6730 8410 6750
rect 8750 6800 8770 6840
rect 8810 6800 8830 6840
rect 8750 6780 8830 6800
rect 10330 6790 10410 6810
rect 8750 6740 9990 6780
rect 8350 6690 8390 6730
rect 8750 6690 8790 6740
rect 9950 6690 9990 6740
rect 10330 6750 10350 6790
rect 10390 6750 10410 6790
rect 10330 6730 10410 6750
rect 10350 6690 10390 6730
rect 8230 6670 8410 6690
rect 8230 6630 8250 6670
rect 8290 6630 8350 6670
rect 8390 6630 8410 6670
rect 8230 6570 8410 6630
rect 8230 6530 8250 6570
rect 8290 6530 8350 6570
rect 8390 6530 8410 6570
rect 8230 6470 8410 6530
rect 8230 6430 8250 6470
rect 8290 6430 8350 6470
rect 8390 6430 8410 6470
rect 8230 6370 8410 6430
rect 8230 6330 8250 6370
rect 8290 6330 8350 6370
rect 8390 6330 8410 6370
rect 8230 6270 8410 6330
rect 8230 6230 8250 6270
rect 8290 6230 8350 6270
rect 8390 6230 8410 6270
rect 8230 6210 8410 6230
rect 8530 6670 8610 6690
rect 8530 6630 8550 6670
rect 8590 6630 8610 6670
rect 8530 6570 8610 6630
rect 8530 6530 8550 6570
rect 8590 6530 8610 6570
rect 8530 6470 8610 6530
rect 8530 6430 8550 6470
rect 8590 6430 8610 6470
rect 8530 6370 8610 6430
rect 8530 6330 8550 6370
rect 8590 6330 8610 6370
rect 8530 6270 8610 6330
rect 8530 6230 8550 6270
rect 8590 6230 8610 6270
rect 8530 6210 8610 6230
rect 8730 6670 8810 6690
rect 8730 6630 8750 6670
rect 8790 6630 8810 6670
rect 8730 6570 8810 6630
rect 8730 6530 8750 6570
rect 8790 6530 8810 6570
rect 8730 6470 8810 6530
rect 8730 6430 8750 6470
rect 8790 6430 8810 6470
rect 8730 6370 8810 6430
rect 8730 6330 8750 6370
rect 8790 6330 8810 6370
rect 8730 6270 8810 6330
rect 8730 6230 8750 6270
rect 8790 6230 8810 6270
rect 8730 6210 8810 6230
rect 8930 6670 9010 6690
rect 8930 6630 8950 6670
rect 8990 6630 9010 6670
rect 8930 6570 9010 6630
rect 8930 6530 8950 6570
rect 8990 6530 9010 6570
rect 8930 6470 9010 6530
rect 8930 6430 8950 6470
rect 8990 6430 9010 6470
rect 8930 6370 9010 6430
rect 8930 6330 8950 6370
rect 8990 6330 9010 6370
rect 8930 6270 9010 6330
rect 8930 6230 8950 6270
rect 8990 6230 9010 6270
rect 8930 6210 9010 6230
rect 9130 6670 9210 6690
rect 9130 6630 9150 6670
rect 9190 6630 9210 6670
rect 9130 6570 9210 6630
rect 9130 6530 9150 6570
rect 9190 6530 9210 6570
rect 9130 6470 9210 6530
rect 9130 6430 9150 6470
rect 9190 6430 9210 6470
rect 9130 6370 9210 6430
rect 9130 6330 9150 6370
rect 9190 6330 9210 6370
rect 9130 6270 9210 6330
rect 9130 6230 9150 6270
rect 9190 6230 9210 6270
rect 9130 6210 9210 6230
rect 9330 6670 9410 6690
rect 9330 6630 9350 6670
rect 9390 6630 9410 6670
rect 9330 6570 9410 6630
rect 9330 6530 9350 6570
rect 9390 6530 9410 6570
rect 9330 6470 9410 6530
rect 9330 6430 9350 6470
rect 9390 6430 9410 6470
rect 9330 6370 9410 6430
rect 9330 6330 9350 6370
rect 9390 6330 9410 6370
rect 9330 6270 9410 6330
rect 9330 6230 9350 6270
rect 9390 6230 9410 6270
rect 9330 6210 9410 6230
rect 9530 6670 9610 6690
rect 9530 6630 9550 6670
rect 9590 6630 9610 6670
rect 9530 6570 9610 6630
rect 9530 6530 9550 6570
rect 9590 6530 9610 6570
rect 9530 6470 9610 6530
rect 9530 6430 9550 6470
rect 9590 6430 9610 6470
rect 9530 6370 9610 6430
rect 9530 6330 9550 6370
rect 9590 6330 9610 6370
rect 9530 6270 9610 6330
rect 9530 6230 9550 6270
rect 9590 6230 9610 6270
rect 9530 6210 9610 6230
rect 9730 6670 9810 6690
rect 9730 6630 9750 6670
rect 9790 6630 9810 6670
rect 9730 6570 9810 6630
rect 9730 6530 9750 6570
rect 9790 6530 9810 6570
rect 9730 6470 9810 6530
rect 9730 6430 9750 6470
rect 9790 6430 9810 6470
rect 9730 6370 9810 6430
rect 9730 6330 9750 6370
rect 9790 6330 9810 6370
rect 9730 6270 9810 6330
rect 9730 6230 9750 6270
rect 9790 6230 9810 6270
rect 9730 6210 9810 6230
rect 9930 6670 10010 6690
rect 9930 6630 9950 6670
rect 9990 6630 10010 6670
rect 9930 6570 10010 6630
rect 9930 6530 9950 6570
rect 9990 6530 10010 6570
rect 9930 6470 10010 6530
rect 9930 6430 9950 6470
rect 9990 6430 10010 6470
rect 9930 6370 10010 6430
rect 9930 6330 9950 6370
rect 9990 6330 10010 6370
rect 9930 6270 10010 6330
rect 9930 6230 9950 6270
rect 9990 6230 10010 6270
rect 9930 6210 10010 6230
rect 10130 6670 10210 6690
rect 10130 6630 10150 6670
rect 10190 6630 10210 6670
rect 10130 6570 10210 6630
rect 10130 6530 10150 6570
rect 10190 6530 10210 6570
rect 10130 6470 10210 6530
rect 10130 6430 10150 6470
rect 10190 6430 10210 6470
rect 10130 6370 10210 6430
rect 10130 6330 10150 6370
rect 10190 6330 10210 6370
rect 10130 6270 10210 6330
rect 10130 6230 10150 6270
rect 10190 6230 10210 6270
rect 10130 6210 10210 6230
rect 10330 6670 10510 6690
rect 10330 6630 10350 6670
rect 10390 6630 10450 6670
rect 10490 6630 10510 6670
rect 10330 6570 10510 6630
rect 10330 6530 10350 6570
rect 10390 6530 10450 6570
rect 10490 6530 10510 6570
rect 10330 6470 10510 6530
rect 10330 6430 10350 6470
rect 10390 6430 10450 6470
rect 10490 6430 10510 6470
rect 10330 6370 10510 6430
rect 10330 6330 10350 6370
rect 10390 6330 10450 6370
rect 10490 6330 10510 6370
rect 10330 6270 10510 6330
rect 10330 6230 10350 6270
rect 10390 6230 10450 6270
rect 10490 6230 10510 6270
rect 10330 6210 10510 6230
rect 9150 6170 9190 6210
rect 9550 6170 9590 6210
rect 9130 6160 9210 6170
rect 9530 6160 9610 6170
rect 4860 6100 4870 6140
rect 4910 6100 4950 6140
rect 4990 6100 5000 6140
rect 7650 6150 9610 6160
rect 7650 6120 9150 6150
rect 4860 6080 5000 6100
rect 9130 6110 9150 6120
rect 9190 6120 9550 6150
rect 9190 6110 9210 6120
rect 9130 6090 9210 6110
rect 9530 6110 9550 6120
rect 9590 6110 9610 6150
rect 9530 6090 9610 6110
rect 1630 6040 1670 6080
rect 1990 6040 2030 6080
rect 2350 6040 2390 6080
rect 2710 6040 2750 6080
rect 3070 6040 3110 6080
rect 3430 6040 3470 6080
rect 3790 6040 3830 6080
rect 4150 6040 4190 6080
rect 4510 6040 4550 6080
rect 4870 6040 4910 6080
rect 1610 6020 1690 6040
rect 1610 5980 1630 6020
rect 1670 5980 1690 6020
rect 1610 5960 1690 5980
rect 1970 6020 2050 6040
rect 1970 5980 1990 6020
rect 2030 5980 2050 6020
rect 1970 5960 2050 5980
rect 2330 6020 2410 6040
rect 2330 5980 2350 6020
rect 2390 5980 2410 6020
rect 2330 5960 2410 5980
rect 2690 6020 2770 6040
rect 2690 5980 2710 6020
rect 2750 5980 2770 6020
rect 2690 5960 2770 5980
rect 3050 6020 3130 6040
rect 3050 5980 3070 6020
rect 3110 5980 3130 6020
rect 3050 5960 3130 5980
rect 3410 6020 3490 6040
rect 3410 5980 3430 6020
rect 3470 5980 3490 6020
rect 3410 5960 3490 5980
rect 3770 6020 3850 6040
rect 3770 5980 3790 6020
rect 3830 5980 3850 6020
rect 3770 5960 3850 5980
rect 4130 6020 4210 6040
rect 4130 5980 4150 6020
rect 4190 5980 4210 6020
rect 4130 5960 4210 5980
rect 4490 6020 4570 6040
rect 4490 5980 4510 6020
rect 4550 5980 4570 6020
rect 4490 5960 4570 5980
rect 4850 6020 4930 6040
rect 4850 5980 4870 6020
rect 4910 5980 4930 6020
rect 4850 5960 4930 5980
rect 1796 5752 1854 5770
rect 1796 5718 1808 5752
rect 1842 5718 1854 5752
rect 1796 5700 1854 5718
rect 1906 5752 1964 5770
rect 1906 5718 1918 5752
rect 1952 5718 1964 5752
rect 1906 5700 1964 5718
rect 2016 5752 2074 5770
rect 2016 5718 2028 5752
rect 2062 5718 2074 5752
rect 2016 5700 2074 5718
rect 2126 5752 2184 5770
rect 2126 5718 2138 5752
rect 2172 5718 2184 5752
rect 2126 5700 2184 5718
rect 2236 5752 2294 5770
rect 2236 5718 2248 5752
rect 2282 5718 2294 5752
rect 2236 5700 2294 5718
rect 2346 5752 2404 5770
rect 2346 5718 2358 5752
rect 2392 5718 2404 5752
rect 2346 5700 2404 5718
rect 2456 5752 2514 5770
rect 2456 5718 2468 5752
rect 2502 5718 2514 5752
rect 2456 5700 2514 5718
rect 2566 5752 2624 5770
rect 2566 5718 2578 5752
rect 2612 5718 2624 5752
rect 2566 5700 2624 5718
rect 2676 5752 2734 5770
rect 2676 5718 2688 5752
rect 2722 5718 2734 5752
rect 2676 5700 2734 5718
rect 2786 5752 2844 5770
rect 2786 5718 2798 5752
rect 2832 5718 2844 5752
rect 2786 5700 2844 5718
rect 3696 5752 3754 5770
rect 3696 5718 3708 5752
rect 3742 5718 3754 5752
rect 3696 5700 3754 5718
rect 3806 5752 3864 5770
rect 3806 5718 3818 5752
rect 3852 5718 3864 5752
rect 3806 5700 3864 5718
rect 3916 5752 3974 5770
rect 3916 5718 3928 5752
rect 3962 5718 3974 5752
rect 3916 5700 3974 5718
rect 4026 5752 4084 5770
rect 4026 5718 4038 5752
rect 4072 5718 4084 5752
rect 4026 5700 4084 5718
rect 4136 5752 4194 5770
rect 4136 5718 4148 5752
rect 4182 5718 4194 5752
rect 4136 5700 4194 5718
rect 4246 5752 4304 5770
rect 4246 5718 4258 5752
rect 4292 5718 4304 5752
rect 4246 5700 4304 5718
rect 4356 5752 4414 5770
rect 4356 5718 4368 5752
rect 4402 5718 4414 5752
rect 4356 5700 4414 5718
rect 4466 5752 4524 5770
rect 4466 5718 4478 5752
rect 4512 5718 4524 5752
rect 4466 5700 4524 5718
rect 4576 5752 4634 5770
rect 4576 5718 4588 5752
rect 4622 5718 4634 5752
rect 4576 5700 4634 5718
rect 4686 5752 4744 5770
rect 4686 5718 4698 5752
rect 4732 5718 4744 5752
rect 4686 5700 4744 5718
rect 1550 5640 1690 5660
rect 1550 5600 1560 5640
rect 1600 5600 1640 5640
rect 1680 5600 1690 5640
rect 1550 5540 1690 5600
rect 1550 5500 1560 5540
rect 1600 5500 1640 5540
rect 1680 5500 1690 5540
rect 1550 5480 1690 5500
rect 1740 5640 1800 5660
rect 1740 5600 1750 5640
rect 1790 5600 1800 5640
rect 1740 5540 1800 5600
rect 1740 5500 1750 5540
rect 1790 5500 1800 5540
rect 1740 5480 1800 5500
rect 1850 5640 1910 5660
rect 1850 5600 1860 5640
rect 1900 5600 1910 5640
rect 1850 5540 1910 5600
rect 1850 5500 1860 5540
rect 1900 5500 1910 5540
rect 1850 5480 1910 5500
rect 1960 5640 2020 5660
rect 1960 5600 1970 5640
rect 2010 5600 2020 5640
rect 1960 5540 2020 5600
rect 1960 5500 1970 5540
rect 2010 5500 2020 5540
rect 1960 5480 2020 5500
rect 2070 5640 2130 5660
rect 2070 5600 2080 5640
rect 2120 5600 2130 5640
rect 2070 5540 2130 5600
rect 2070 5500 2080 5540
rect 2120 5500 2130 5540
rect 2070 5480 2130 5500
rect 2180 5640 2240 5660
rect 2180 5600 2190 5640
rect 2230 5600 2240 5640
rect 2180 5540 2240 5600
rect 2180 5500 2190 5540
rect 2230 5500 2240 5540
rect 2180 5480 2240 5500
rect 2290 5640 2350 5660
rect 2290 5600 2300 5640
rect 2340 5600 2350 5640
rect 2290 5540 2350 5600
rect 2290 5500 2300 5540
rect 2340 5500 2350 5540
rect 2290 5480 2350 5500
rect 2400 5640 2460 5660
rect 2400 5600 2410 5640
rect 2450 5600 2460 5640
rect 2400 5540 2460 5600
rect 2400 5500 2410 5540
rect 2450 5500 2460 5540
rect 2400 5480 2460 5500
rect 2510 5640 2570 5660
rect 2510 5600 2520 5640
rect 2560 5600 2570 5640
rect 2510 5540 2570 5600
rect 2510 5500 2520 5540
rect 2560 5500 2570 5540
rect 2510 5480 2570 5500
rect 2620 5640 2680 5660
rect 2620 5600 2630 5640
rect 2670 5600 2680 5640
rect 2620 5540 2680 5600
rect 2620 5500 2630 5540
rect 2670 5500 2680 5540
rect 2620 5480 2680 5500
rect 2730 5640 2790 5660
rect 2730 5600 2740 5640
rect 2780 5600 2790 5640
rect 2730 5540 2790 5600
rect 2730 5500 2740 5540
rect 2780 5500 2790 5540
rect 2730 5480 2790 5500
rect 2840 5640 2900 5660
rect 2840 5600 2850 5640
rect 2890 5600 2900 5640
rect 2840 5540 2900 5600
rect 2840 5500 2850 5540
rect 2890 5500 2900 5540
rect 2840 5480 2900 5500
rect 2950 5640 3090 5660
rect 2950 5600 2960 5640
rect 3000 5600 3040 5640
rect 3080 5600 3090 5640
rect 2950 5540 3090 5600
rect 2950 5500 2960 5540
rect 3000 5500 3040 5540
rect 3080 5500 3090 5540
rect 2950 5480 3090 5500
rect 3450 5640 3590 5660
rect 3450 5600 3460 5640
rect 3500 5600 3540 5640
rect 3580 5600 3590 5640
rect 3450 5540 3590 5600
rect 3450 5500 3460 5540
rect 3500 5500 3540 5540
rect 3580 5500 3590 5540
rect 3450 5480 3590 5500
rect 3640 5640 3700 5660
rect 3640 5600 3650 5640
rect 3690 5600 3700 5640
rect 3640 5540 3700 5600
rect 3640 5500 3650 5540
rect 3690 5500 3700 5540
rect 3640 5480 3700 5500
rect 3750 5640 3810 5660
rect 3750 5600 3760 5640
rect 3800 5600 3810 5640
rect 3750 5540 3810 5600
rect 3750 5500 3760 5540
rect 3800 5500 3810 5540
rect 3750 5480 3810 5500
rect 3860 5640 3920 5660
rect 3860 5600 3870 5640
rect 3910 5600 3920 5640
rect 3860 5540 3920 5600
rect 3860 5500 3870 5540
rect 3910 5500 3920 5540
rect 3860 5480 3920 5500
rect 3970 5640 4030 5660
rect 3970 5600 3980 5640
rect 4020 5600 4030 5640
rect 3970 5540 4030 5600
rect 3970 5500 3980 5540
rect 4020 5500 4030 5540
rect 3970 5480 4030 5500
rect 4080 5640 4140 5660
rect 4080 5600 4090 5640
rect 4130 5600 4140 5640
rect 4080 5540 4140 5600
rect 4080 5500 4090 5540
rect 4130 5500 4140 5540
rect 4080 5480 4140 5500
rect 4190 5640 4250 5660
rect 4190 5600 4200 5640
rect 4240 5600 4250 5640
rect 4190 5540 4250 5600
rect 4190 5500 4200 5540
rect 4240 5500 4250 5540
rect 4190 5480 4250 5500
rect 4300 5640 4360 5660
rect 4300 5600 4310 5640
rect 4350 5600 4360 5640
rect 4300 5540 4360 5600
rect 4300 5500 4310 5540
rect 4350 5500 4360 5540
rect 4300 5480 4360 5500
rect 4410 5640 4470 5660
rect 4410 5600 4420 5640
rect 4460 5600 4470 5640
rect 4410 5540 4470 5600
rect 4410 5500 4420 5540
rect 4460 5500 4470 5540
rect 4410 5480 4470 5500
rect 4520 5640 4580 5660
rect 4520 5600 4530 5640
rect 4570 5600 4580 5640
rect 4520 5540 4580 5600
rect 4520 5500 4530 5540
rect 4570 5500 4580 5540
rect 4520 5480 4580 5500
rect 4630 5640 4690 5660
rect 4630 5600 4640 5640
rect 4680 5600 4690 5640
rect 4630 5540 4690 5600
rect 4630 5500 4640 5540
rect 4680 5500 4690 5540
rect 4630 5480 4690 5500
rect 4740 5640 4800 5660
rect 4740 5600 4750 5640
rect 4790 5600 4800 5640
rect 4740 5540 4800 5600
rect 4740 5500 4750 5540
rect 4790 5500 4800 5540
rect 4740 5480 4800 5500
rect 4850 5640 4990 5660
rect 4850 5600 4860 5640
rect 4900 5600 4940 5640
rect 4980 5600 4990 5640
rect 4850 5540 4990 5600
rect 4850 5500 4860 5540
rect 4900 5500 4940 5540
rect 4980 5500 4990 5540
rect 4850 5480 4990 5500
rect 11670 5440 11710 6034
rect 11750 5440 11850 5460
rect 1620 5420 1700 5440
rect 1620 5380 1640 5420
rect 1680 5380 1700 5420
rect 1620 5360 1700 5380
rect 2940 5420 3020 5440
rect 2940 5380 2960 5420
rect 3000 5380 3020 5420
rect 2940 5360 3020 5380
rect 3520 5420 3600 5440
rect 3520 5380 3540 5420
rect 3580 5380 3600 5420
rect 3520 5360 3600 5380
rect 4840 5420 4920 5440
rect 4840 5380 4860 5420
rect 4900 5380 4920 5420
rect 11670 5400 11770 5440
rect 4840 5360 4920 5380
rect 11750 5380 11770 5400
rect 11830 5380 11850 5440
rect 11750 5360 11850 5380
rect 11590 5090 11700 5110
rect 11590 5020 11610 5090
rect 11680 5020 11700 5090
rect 11590 5000 11700 5020
rect 1720 4930 1820 4950
rect 1720 4920 1880 4930
rect 1720 4880 1750 4920
rect 1790 4890 1880 4920
rect 1920 4890 1980 4930
rect 2020 4890 2080 4930
rect 2120 4890 2180 4930
rect 2220 4890 2280 4930
rect 2320 4890 2380 4930
rect 2420 4890 2480 4930
rect 2520 4890 2580 4930
rect 2620 4890 2680 4930
rect 2720 4890 2780 4930
rect 2820 4890 2880 4930
rect 2920 4890 2980 4930
rect 3020 4890 3080 4930
rect 3120 4890 3180 4930
rect 3220 4890 3280 4930
rect 3320 4890 3380 4930
rect 3420 4890 3480 4930
rect 3520 4890 3580 4930
rect 3620 4890 3680 4930
rect 3720 4890 3780 4930
rect 3820 4890 3880 4930
rect 3920 4890 3980 4930
rect 4020 4890 4080 4930
rect 4120 4890 4180 4930
rect 4220 4890 4280 4930
rect 4320 4890 4380 4930
rect 4420 4890 4480 4930
rect 4520 4890 4580 4930
rect 4620 4890 4680 4930
rect 4720 4890 4780 4930
rect 4820 4890 4880 4930
rect 4920 4890 4980 4930
rect 5020 4890 5080 4930
rect 5120 4890 5180 4930
rect 5220 4890 5280 4930
rect 5320 4890 5380 4930
rect 5420 4890 5480 4930
rect 5520 4890 5580 4930
rect 5620 4890 5680 4930
rect 5720 4890 5780 4930
rect 5820 4890 5880 4930
rect 5920 4890 5980 4930
rect 6020 4890 6080 4930
rect 6120 4890 6180 4930
rect 6220 4890 6280 4930
rect 6320 4890 6380 4930
rect 6420 4890 6480 4930
rect 6520 4890 6580 4930
rect 6620 4890 6680 4930
rect 6720 4890 6780 4930
rect 6820 4890 6880 4930
rect 6920 4890 7040 4930
rect 1790 4880 1820 4890
rect 1720 4850 1820 4880
rect 2160 4720 2200 4890
rect 2380 4720 2420 4890
rect 2550 4820 2630 4840
rect 2550 4780 2570 4820
rect 2610 4780 2630 4820
rect 2550 4760 2630 4780
rect 2070 4700 2210 4720
rect 2070 4660 2080 4700
rect 2120 4660 2160 4700
rect 2200 4660 2210 4700
rect 2070 4600 2210 4660
rect 2070 4560 2080 4600
rect 2120 4560 2160 4600
rect 2200 4560 2210 4600
rect 2070 4540 2210 4560
rect 2260 4700 2320 4720
rect 2260 4660 2270 4700
rect 2310 4660 2320 4700
rect 2260 4600 2320 4660
rect 2260 4560 2270 4600
rect 2310 4560 2320 4600
rect 2260 4540 2320 4560
rect 2370 4700 2430 4720
rect 2370 4660 2380 4700
rect 2420 4660 2430 4700
rect 2370 4600 2430 4660
rect 2370 4560 2380 4600
rect 2420 4560 2430 4600
rect 2370 4540 2430 4560
rect 1930 4470 2010 4490
rect 1930 4430 1950 4470
rect 1990 4430 2010 4470
rect 1930 4410 2010 4430
rect 2260 4380 2300 4540
rect 2350 4480 2430 4500
rect 2350 4440 2370 4480
rect 2410 4460 2430 4480
rect 2590 4460 2630 4760
rect 2680 4720 2720 4890
rect 2900 4720 2940 4890
rect 3060 4720 3100 4890
rect 3280 4720 3320 4890
rect 3580 4720 3620 4890
rect 3800 4720 3840 4890
rect 4100 4720 4140 4890
rect 4270 4820 4350 4840
rect 4270 4780 4290 4820
rect 4330 4780 4350 4820
rect 4270 4760 4350 4780
rect 4540 4720 4580 4890
rect 4870 4720 4910 4890
rect 5300 4720 5340 4890
rect 5690 4720 5730 4890
rect 6080 4720 6120 4890
rect 6340 4820 6420 4840
rect 6340 4780 6360 4820
rect 6400 4780 6420 4820
rect 6340 4760 6420 4780
rect 6360 4720 6400 4760
rect 2670 4700 2730 4720
rect 2670 4660 2680 4700
rect 2720 4660 2730 4700
rect 2670 4600 2730 4660
rect 2670 4560 2680 4600
rect 2720 4560 2730 4600
rect 2670 4540 2730 4560
rect 2780 4700 2840 4720
rect 2780 4660 2790 4700
rect 2830 4660 2840 4700
rect 2780 4600 2840 4660
rect 2780 4560 2790 4600
rect 2830 4560 2840 4600
rect 2780 4540 2840 4560
rect 2890 4700 3110 4720
rect 2890 4660 2900 4700
rect 2940 4660 2980 4700
rect 3020 4660 3060 4700
rect 3100 4660 3110 4700
rect 2890 4600 3110 4660
rect 2890 4560 2900 4600
rect 2940 4560 2980 4600
rect 3020 4560 3060 4600
rect 3100 4560 3110 4600
rect 2890 4540 3110 4560
rect 3160 4700 3220 4720
rect 3160 4660 3170 4700
rect 3210 4660 3220 4700
rect 3160 4600 3220 4660
rect 3160 4560 3170 4600
rect 3210 4560 3220 4600
rect 3160 4540 3220 4560
rect 3270 4700 3330 4720
rect 3270 4660 3280 4700
rect 3320 4660 3330 4700
rect 3270 4600 3330 4660
rect 3270 4560 3280 4600
rect 3320 4560 3330 4600
rect 3270 4540 3330 4560
rect 3570 4700 3630 4720
rect 3570 4660 3580 4700
rect 3620 4660 3630 4700
rect 3570 4600 3630 4660
rect 3570 4560 3580 4600
rect 3620 4560 3630 4600
rect 3570 4540 3630 4560
rect 3680 4700 3740 4720
rect 3680 4660 3690 4700
rect 3730 4660 3740 4700
rect 3680 4600 3740 4660
rect 3680 4560 3690 4600
rect 3730 4560 3740 4600
rect 3680 4540 3740 4560
rect 3790 4700 3930 4720
rect 3790 4660 3800 4700
rect 3840 4660 3880 4700
rect 3920 4660 3930 4700
rect 3790 4600 3930 4660
rect 3790 4560 3800 4600
rect 3840 4560 3880 4600
rect 3920 4560 3930 4600
rect 3790 4540 3930 4560
rect 4010 4700 4150 4720
rect 4010 4660 4020 4700
rect 4060 4660 4100 4700
rect 4140 4660 4150 4700
rect 4010 4600 4150 4660
rect 4010 4560 4020 4600
rect 4060 4560 4100 4600
rect 4140 4560 4150 4600
rect 4010 4540 4150 4560
rect 4200 4700 4260 4720
rect 4200 4660 4210 4700
rect 4250 4660 4260 4700
rect 4200 4600 4260 4660
rect 4200 4560 4210 4600
rect 4250 4560 4260 4600
rect 4200 4540 4260 4560
rect 4310 4700 4370 4720
rect 4310 4660 4320 4700
rect 4360 4660 4370 4700
rect 4310 4600 4370 4660
rect 4310 4560 4320 4600
rect 4360 4560 4370 4600
rect 4310 4540 4370 4560
rect 4450 4700 4590 4720
rect 4450 4660 4460 4700
rect 4500 4660 4540 4700
rect 4580 4660 4590 4700
rect 4450 4600 4590 4660
rect 4450 4560 4460 4600
rect 4500 4560 4540 4600
rect 4580 4560 4590 4600
rect 4450 4540 4590 4560
rect 4640 4700 4700 4720
rect 4640 4660 4650 4700
rect 4690 4660 4700 4700
rect 4640 4600 4700 4660
rect 4640 4560 4650 4600
rect 4690 4560 4700 4600
rect 4640 4540 4700 4560
rect 4780 4700 4920 4720
rect 4780 4660 4790 4700
rect 4830 4660 4870 4700
rect 4910 4660 4920 4700
rect 4780 4600 4920 4660
rect 4780 4560 4790 4600
rect 4830 4560 4870 4600
rect 4910 4560 4920 4600
rect 4780 4540 4920 4560
rect 4970 4700 5030 4720
rect 4970 4660 4980 4700
rect 5020 4660 5030 4700
rect 4970 4600 5030 4660
rect 4970 4560 4980 4600
rect 5020 4560 5030 4600
rect 4970 4540 5030 4560
rect 5200 4700 5360 4720
rect 5200 4660 5210 4700
rect 5250 4660 5300 4700
rect 5340 4660 5360 4700
rect 5200 4600 5360 4660
rect 5200 4560 5210 4600
rect 5250 4560 5300 4600
rect 5340 4560 5360 4600
rect 5200 4540 5360 4560
rect 5410 4700 5490 4720
rect 5410 4660 5430 4700
rect 5470 4660 5490 4700
rect 5410 4600 5490 4660
rect 5410 4560 5430 4600
rect 5470 4560 5490 4600
rect 5410 4540 5490 4560
rect 5590 4700 5750 4720
rect 5590 4660 5600 4700
rect 5640 4660 5690 4700
rect 5730 4660 5750 4700
rect 5590 4600 5750 4660
rect 5590 4560 5600 4600
rect 5640 4560 5690 4600
rect 5730 4560 5750 4600
rect 5590 4540 5750 4560
rect 5800 4700 5880 4720
rect 5800 4660 5820 4700
rect 5860 4660 5880 4700
rect 5800 4600 5880 4660
rect 5800 4560 5820 4600
rect 5860 4560 5880 4600
rect 5800 4540 5880 4560
rect 5980 4700 6140 4720
rect 5980 4660 5990 4700
rect 6030 4660 6080 4700
rect 6120 4660 6140 4700
rect 5980 4600 6140 4660
rect 5980 4560 5990 4600
rect 6030 4560 6080 4600
rect 6120 4560 6140 4600
rect 5980 4540 6140 4560
rect 6190 4700 6270 4720
rect 6190 4660 6210 4700
rect 6250 4660 6270 4700
rect 6190 4600 6270 4660
rect 6190 4560 6210 4600
rect 6250 4560 6270 4600
rect 6190 4540 6270 4560
rect 6350 4700 6430 4720
rect 6350 4660 6370 4700
rect 6410 4660 6430 4700
rect 6350 4600 6430 4660
rect 6350 4560 6370 4600
rect 6410 4560 6430 4600
rect 6350 4540 6430 4560
rect 6480 4700 6560 4720
rect 6480 4660 6500 4700
rect 6540 4660 6560 4700
rect 6480 4600 6560 4660
rect 6480 4560 6500 4600
rect 6540 4560 6560 4600
rect 6480 4540 6560 4560
rect 2410 4440 2630 4460
rect 2350 4420 2630 4440
rect 2260 4340 2420 4380
rect 2380 4300 2420 4340
rect 2070 4280 2210 4300
rect 2070 4240 2080 4280
rect 2120 4240 2160 4280
rect 2200 4240 2210 4280
rect 2070 4180 2210 4240
rect 2070 4140 2080 4180
rect 2120 4140 2160 4180
rect 2200 4140 2210 4180
rect 2070 4080 2210 4140
rect 2070 4040 2080 4080
rect 2120 4040 2160 4080
rect 2200 4040 2210 4080
rect 2070 3980 2210 4040
rect 2070 3940 2080 3980
rect 2120 3940 2160 3980
rect 2200 3940 2210 3980
rect 2070 3920 2210 3940
rect 2260 4280 2320 4300
rect 2260 4240 2270 4280
rect 2310 4240 2320 4280
rect 2260 4180 2320 4240
rect 2260 4140 2270 4180
rect 2310 4140 2320 4180
rect 2260 4080 2320 4140
rect 2260 4040 2270 4080
rect 2310 4040 2320 4080
rect 2260 3980 2320 4040
rect 2260 3940 2270 3980
rect 2310 3940 2320 3980
rect 2260 3920 2320 3940
rect 2370 4280 2430 4300
rect 2370 4240 2380 4280
rect 2420 4240 2430 4280
rect 2370 4180 2430 4240
rect 2370 4140 2380 4180
rect 2420 4140 2430 4180
rect 2370 4080 2430 4140
rect 2370 4040 2380 4080
rect 2420 4040 2430 4080
rect 2370 3980 2430 4040
rect 2370 3940 2380 3980
rect 2420 3970 2430 3980
rect 2470 3980 2550 4000
rect 2470 3970 2490 3980
rect 2420 3940 2490 3970
rect 2530 3940 2550 3980
rect 2370 3920 2550 3940
rect 2590 3960 2630 4420
rect 2790 4380 2830 4540
rect 2680 4340 2830 4380
rect 2870 4400 2950 4420
rect 2870 4360 2890 4400
rect 2930 4380 2950 4400
rect 3160 4380 3200 4540
rect 3250 4480 3330 4500
rect 3250 4440 3270 4480
rect 3310 4460 3330 4480
rect 3310 4440 3530 4460
rect 3250 4420 3530 4440
rect 2930 4360 3320 4380
rect 2870 4340 3320 4360
rect 2680 4300 2720 4340
rect 3280 4300 3320 4340
rect 2670 4280 2730 4300
rect 2670 4240 2680 4280
rect 2720 4240 2730 4280
rect 2670 4180 2730 4240
rect 2670 4140 2680 4180
rect 2720 4140 2730 4180
rect 2670 4080 2730 4140
rect 2670 4040 2680 4080
rect 2720 4040 2730 4080
rect 2670 3980 2730 4040
rect 2670 3960 2680 3980
rect 2590 3940 2680 3960
rect 2720 3940 2730 3980
rect 2590 3920 2730 3940
rect 2780 4280 2840 4300
rect 2780 4240 2790 4280
rect 2830 4240 2840 4280
rect 2780 4180 2840 4240
rect 2780 4140 2790 4180
rect 2830 4140 2840 4180
rect 2780 4080 2840 4140
rect 2780 4040 2790 4080
rect 2830 4040 2840 4080
rect 2780 3980 2840 4040
rect 2780 3940 2790 3980
rect 2830 3940 2840 3980
rect 2780 3920 2840 3940
rect 2890 4280 3110 4300
rect 2890 4240 2900 4280
rect 2940 4240 2980 4280
rect 3020 4240 3060 4280
rect 3100 4240 3110 4280
rect 2890 4180 3110 4240
rect 2890 4140 2900 4180
rect 2940 4140 2980 4180
rect 3020 4140 3060 4180
rect 3100 4140 3110 4180
rect 2890 4080 3110 4140
rect 2890 4040 2900 4080
rect 2940 4040 2980 4080
rect 3020 4040 3060 4080
rect 3100 4040 3110 4080
rect 2890 3980 3110 4040
rect 2890 3940 2900 3980
rect 2940 3940 2980 3980
rect 3020 3940 3060 3980
rect 3100 3940 3110 3980
rect 2890 3920 3110 3940
rect 3160 4280 3220 4300
rect 3160 4240 3170 4280
rect 3210 4240 3220 4280
rect 3160 4180 3220 4240
rect 3160 4140 3170 4180
rect 3210 4140 3220 4180
rect 3160 4080 3220 4140
rect 3160 4040 3170 4080
rect 3210 4040 3220 4080
rect 3160 3980 3220 4040
rect 3160 3940 3170 3980
rect 3210 3940 3220 3980
rect 3160 3920 3220 3940
rect 3270 4280 3330 4300
rect 3270 4240 3280 4280
rect 3320 4240 3330 4280
rect 3270 4180 3330 4240
rect 3270 4140 3280 4180
rect 3320 4140 3330 4180
rect 3270 4080 3330 4140
rect 3270 4040 3280 4080
rect 3320 4040 3330 4080
rect 3270 3980 3330 4040
rect 3270 3940 3280 3980
rect 3320 3970 3330 3980
rect 3370 3980 3450 4000
rect 3370 3970 3390 3980
rect 3320 3940 3390 3970
rect 3430 3940 3450 3980
rect 3270 3920 3450 3940
rect 3490 3960 3530 4420
rect 3690 4380 3730 4540
rect 3840 4470 3920 4490
rect 3840 4430 3860 4470
rect 3900 4430 3920 4470
rect 3840 4410 3920 4430
rect 4320 4450 4360 4540
rect 4660 4450 4700 4540
rect 4990 4450 5030 4540
rect 5140 4460 5220 4480
rect 4320 4430 4430 4450
rect 4320 4410 4370 4430
rect 3580 4340 3730 4380
rect 4210 4390 4370 4410
rect 4410 4390 4430 4430
rect 4210 4370 4430 4390
rect 4660 4430 4760 4450
rect 4660 4390 4700 4430
rect 4740 4390 4760 4430
rect 4660 4370 4760 4390
rect 4990 4430 5090 4450
rect 4990 4390 5030 4430
rect 5070 4390 5090 4430
rect 5140 4420 5160 4460
rect 5200 4420 5220 4460
rect 5140 4400 5220 4420
rect 5450 4430 5490 4540
rect 5840 4460 5880 4540
rect 6100 4480 6180 4500
rect 6100 4460 6120 4480
rect 5710 4430 5790 4450
rect 4990 4370 5090 4390
rect 5450 4390 5730 4430
rect 5770 4390 5790 4430
rect 3580 4300 3620 4340
rect 4210 4300 4250 4370
rect 4660 4300 4700 4370
rect 4990 4300 5030 4370
rect 5450 4300 5490 4390
rect 5710 4370 5790 4390
rect 5840 4440 6120 4460
rect 6160 4440 6180 4480
rect 5840 4420 6180 4440
rect 6230 4420 6270 4540
rect 5840 4300 5880 4420
rect 6230 4400 6310 4420
rect 6230 4360 6250 4400
rect 6290 4360 6310 4400
rect 6230 4340 6310 4360
rect 6230 4300 6270 4340
rect 6370 4300 6410 4540
rect 6500 4500 6540 4540
rect 7850 4520 7900 4560
rect 7940 4520 8000 4560
rect 8040 4520 8100 4560
rect 8140 4520 8200 4560
rect 8240 4520 8300 4560
rect 8340 4520 8400 4560
rect 8440 4520 8500 4560
rect 8540 4520 8600 4560
rect 8640 4520 8700 4560
rect 8740 4520 8800 4560
rect 8840 4520 8900 4560
rect 8940 4520 9000 4560
rect 9040 4520 9100 4560
rect 9140 4520 9200 4560
rect 9240 4520 9300 4560
rect 9340 4520 9400 4560
rect 9440 4520 9500 4560
rect 9540 4520 9600 4560
rect 9640 4520 9700 4560
rect 9740 4520 9800 4560
rect 9840 4520 9900 4560
rect 9940 4520 10000 4560
rect 10040 4520 10100 4560
rect 10140 4520 10200 4560
rect 10240 4520 10300 4560
rect 10340 4520 10400 4560
rect 10440 4520 10500 4560
rect 10540 4520 10600 4560
rect 10640 4520 10700 4560
rect 10740 4520 10800 4560
rect 10840 4520 10900 4560
rect 10940 4520 11000 4560
rect 11040 4520 11070 4560
rect 6500 4460 6930 4500
rect 6500 4300 6540 4460
rect 6890 4420 6930 4460
rect 8150 4450 8230 4520
rect 6640 4400 6720 4420
rect 6640 4360 6660 4400
rect 6700 4360 6720 4400
rect 6640 4340 6720 4360
rect 6880 4400 6960 4420
rect 6880 4360 6900 4400
rect 6940 4360 6960 4400
rect 6880 4340 6960 4360
rect 8150 4410 8170 4450
rect 8210 4410 8230 4450
rect 8150 4350 8230 4410
rect 6890 4300 6930 4340
rect 8050 4330 8230 4350
rect 3570 4280 3630 4300
rect 3570 4240 3580 4280
rect 3620 4240 3630 4280
rect 3570 4180 3630 4240
rect 3570 4140 3580 4180
rect 3620 4140 3630 4180
rect 3570 4080 3630 4140
rect 3570 4040 3580 4080
rect 3620 4040 3630 4080
rect 3570 3980 3630 4040
rect 3570 3960 3580 3980
rect 3490 3940 3580 3960
rect 3620 3940 3630 3980
rect 3490 3920 3630 3940
rect 3680 4280 3740 4300
rect 3680 4240 3690 4280
rect 3730 4240 3740 4280
rect 3680 4180 3740 4240
rect 3680 4140 3690 4180
rect 3730 4140 3740 4180
rect 3680 4080 3740 4140
rect 3680 4040 3690 4080
rect 3730 4040 3740 4080
rect 3680 3980 3740 4040
rect 3680 3940 3690 3980
rect 3730 3940 3740 3980
rect 3680 3920 3740 3940
rect 3790 4280 3930 4300
rect 3790 4240 3800 4280
rect 3840 4240 3880 4280
rect 3920 4240 3930 4280
rect 3790 4180 3930 4240
rect 3790 4140 3800 4180
rect 3840 4140 3880 4180
rect 3920 4140 3930 4180
rect 3790 4080 3930 4140
rect 3790 4040 3800 4080
rect 3840 4040 3880 4080
rect 3920 4040 3930 4080
rect 3790 3980 3930 4040
rect 3790 3940 3800 3980
rect 3840 3940 3880 3980
rect 3920 3940 3930 3980
rect 3790 3920 3930 3940
rect 4010 4280 4150 4300
rect 4010 4240 4020 4280
rect 4060 4240 4100 4280
rect 4140 4240 4150 4280
rect 4010 4180 4150 4240
rect 4010 4140 4020 4180
rect 4060 4140 4100 4180
rect 4140 4140 4150 4180
rect 4010 4080 4150 4140
rect 4010 4040 4020 4080
rect 4060 4040 4100 4080
rect 4140 4040 4150 4080
rect 4010 3980 4150 4040
rect 4010 3940 4020 3980
rect 4060 3940 4100 3980
rect 4140 3940 4150 3980
rect 4010 3920 4150 3940
rect 4200 4280 4260 4300
rect 4200 4240 4210 4280
rect 4250 4240 4260 4280
rect 4200 4180 4260 4240
rect 4200 4140 4210 4180
rect 4250 4140 4260 4180
rect 4200 4080 4260 4140
rect 4200 4040 4210 4080
rect 4250 4040 4260 4080
rect 4200 3980 4260 4040
rect 4200 3940 4210 3980
rect 4250 3940 4260 3980
rect 4200 3920 4260 3940
rect 4310 4280 4370 4300
rect 4310 4240 4320 4280
rect 4360 4240 4370 4280
rect 4310 4180 4370 4240
rect 4310 4140 4320 4180
rect 4360 4140 4370 4180
rect 4310 4080 4370 4140
rect 4310 4040 4320 4080
rect 4360 4040 4370 4080
rect 4310 3980 4370 4040
rect 4310 3940 4320 3980
rect 4360 3940 4370 3980
rect 4310 3920 4370 3940
rect 4450 4280 4590 4300
rect 4450 4240 4460 4280
rect 4500 4240 4540 4280
rect 4580 4240 4590 4280
rect 4450 4180 4590 4240
rect 4450 4140 4460 4180
rect 4500 4140 4540 4180
rect 4580 4140 4590 4180
rect 4450 4080 4590 4140
rect 4450 4040 4460 4080
rect 4500 4040 4540 4080
rect 4580 4040 4590 4080
rect 4450 3980 4590 4040
rect 4450 3940 4460 3980
rect 4500 3940 4540 3980
rect 4580 3940 4590 3980
rect 4450 3920 4590 3940
rect 4640 4280 4700 4300
rect 4640 4240 4650 4280
rect 4690 4240 4700 4280
rect 4640 4180 4700 4240
rect 4640 4140 4650 4180
rect 4690 4140 4700 4180
rect 4640 4080 4700 4140
rect 4640 4040 4650 4080
rect 4690 4040 4700 4080
rect 4640 3980 4700 4040
rect 4640 3940 4650 3980
rect 4690 3940 4700 3980
rect 4640 3920 4700 3940
rect 4780 4280 4920 4300
rect 4780 4240 4790 4280
rect 4830 4240 4870 4280
rect 4910 4240 4920 4280
rect 4780 4180 4920 4240
rect 4780 4140 4790 4180
rect 4830 4140 4870 4180
rect 4910 4140 4920 4180
rect 4780 4080 4920 4140
rect 4780 4040 4790 4080
rect 4830 4040 4870 4080
rect 4910 4040 4920 4080
rect 4780 3980 4920 4040
rect 4780 3940 4790 3980
rect 4830 3940 4870 3980
rect 4910 3940 4920 3980
rect 4780 3920 4920 3940
rect 4970 4280 5030 4300
rect 4970 4240 4980 4280
rect 5020 4240 5030 4280
rect 4970 4180 5030 4240
rect 4970 4140 4980 4180
rect 5020 4140 5030 4180
rect 4970 4080 5030 4140
rect 4970 4040 4980 4080
rect 5020 4040 5030 4080
rect 4970 3980 5030 4040
rect 4970 3940 4980 3980
rect 5020 3940 5030 3980
rect 4970 3920 5030 3940
rect 5180 4280 5360 4300
rect 5180 4240 5200 4280
rect 5240 4240 5300 4280
rect 5340 4240 5360 4280
rect 5180 4180 5360 4240
rect 5180 4140 5200 4180
rect 5240 4140 5300 4180
rect 5340 4140 5360 4180
rect 5180 4080 5360 4140
rect 5180 4040 5200 4080
rect 5240 4040 5300 4080
rect 5340 4040 5360 4080
rect 5180 3980 5360 4040
rect 5180 3940 5200 3980
rect 5240 3940 5300 3980
rect 5340 3940 5360 3980
rect 5180 3920 5360 3940
rect 5410 4280 5490 4300
rect 5410 4240 5430 4280
rect 5470 4240 5490 4280
rect 5410 4180 5490 4240
rect 5410 4140 5430 4180
rect 5470 4140 5490 4180
rect 5410 4080 5490 4140
rect 5410 4040 5430 4080
rect 5470 4040 5490 4080
rect 5410 3980 5490 4040
rect 5410 3940 5430 3980
rect 5470 3940 5490 3980
rect 5410 3920 5490 3940
rect 5570 4280 5750 4300
rect 5570 4240 5590 4280
rect 5630 4240 5690 4280
rect 5730 4240 5750 4280
rect 5570 4180 5750 4240
rect 5570 4140 5590 4180
rect 5630 4140 5690 4180
rect 5730 4140 5750 4180
rect 5570 4080 5750 4140
rect 5570 4040 5590 4080
rect 5630 4040 5690 4080
rect 5730 4040 5750 4080
rect 5570 3980 5750 4040
rect 5570 3940 5590 3980
rect 5630 3940 5690 3980
rect 5730 3940 5750 3980
rect 5570 3920 5750 3940
rect 5800 4280 5880 4300
rect 5800 4240 5820 4280
rect 5860 4240 5880 4280
rect 5800 4180 5880 4240
rect 5800 4140 5820 4180
rect 5860 4140 5880 4180
rect 5800 4080 5880 4140
rect 5800 4040 5820 4080
rect 5860 4040 5880 4080
rect 5800 3980 5880 4040
rect 5800 3940 5820 3980
rect 5860 3940 5880 3980
rect 5800 3920 5880 3940
rect 5960 4280 6140 4300
rect 5960 4240 5980 4280
rect 6020 4240 6080 4280
rect 6120 4240 6140 4280
rect 5960 4180 6140 4240
rect 5960 4140 5980 4180
rect 6020 4140 6080 4180
rect 6120 4140 6140 4180
rect 5960 4080 6140 4140
rect 5960 4040 5980 4080
rect 6020 4040 6080 4080
rect 6120 4040 6140 4080
rect 5960 3980 6140 4040
rect 5960 3940 5980 3980
rect 6020 3940 6080 3980
rect 6120 3940 6140 3980
rect 5960 3920 6140 3940
rect 6190 4280 6270 4300
rect 6190 4240 6210 4280
rect 6250 4240 6270 4280
rect 6190 4180 6270 4240
rect 6190 4140 6210 4180
rect 6250 4140 6270 4180
rect 6190 4080 6270 4140
rect 6190 4040 6210 4080
rect 6250 4040 6270 4080
rect 6190 3980 6270 4040
rect 6190 3940 6210 3980
rect 6250 3940 6270 3980
rect 6190 3920 6270 3940
rect 6350 4280 6430 4300
rect 6350 4240 6370 4280
rect 6410 4240 6430 4280
rect 6350 4180 6430 4240
rect 6350 4140 6370 4180
rect 6410 4140 6430 4180
rect 6350 4080 6430 4140
rect 6350 4040 6370 4080
rect 6410 4040 6430 4080
rect 6350 3980 6430 4040
rect 6350 3940 6370 3980
rect 6410 3940 6430 3980
rect 6350 3920 6430 3940
rect 6480 4280 6560 4300
rect 6480 4240 6500 4280
rect 6540 4240 6560 4280
rect 6480 4180 6560 4240
rect 6480 4140 6500 4180
rect 6540 4140 6560 4180
rect 6480 4080 6560 4140
rect 6480 4040 6500 4080
rect 6540 4040 6560 4080
rect 6480 3980 6560 4040
rect 6480 3940 6500 3980
rect 6540 3940 6560 3980
rect 6480 3920 6560 3940
rect 6640 4280 6820 4300
rect 6640 4240 6660 4280
rect 6700 4240 6760 4280
rect 6800 4240 6820 4280
rect 6640 4180 6820 4240
rect 6640 4140 6660 4180
rect 6700 4140 6760 4180
rect 6800 4140 6820 4180
rect 6640 4080 6820 4140
rect 6640 4040 6660 4080
rect 6700 4040 6760 4080
rect 6800 4040 6820 4080
rect 6640 3980 6820 4040
rect 6640 3940 6660 3980
rect 6700 3940 6760 3980
rect 6800 3940 6820 3980
rect 6640 3920 6820 3940
rect 6870 4280 6950 4300
rect 6870 4240 6890 4280
rect 6930 4240 6950 4280
rect 6870 4180 6950 4240
rect 6870 4140 6890 4180
rect 6930 4140 6950 4180
rect 6870 4080 6950 4140
rect 6870 4040 6890 4080
rect 6930 4040 6950 4080
rect 6870 3980 6950 4040
rect 6870 3940 6890 3980
rect 6930 3940 6950 3980
rect 8050 4290 8070 4330
rect 8110 4290 8170 4330
rect 8210 4290 8230 4330
rect 8050 4230 8230 4290
rect 8050 4190 8070 4230
rect 8110 4190 8170 4230
rect 8210 4190 8230 4230
rect 8050 4130 8230 4190
rect 8050 4090 8070 4130
rect 8110 4090 8170 4130
rect 8210 4090 8230 4130
rect 8050 4030 8230 4090
rect 8050 3990 8070 4030
rect 8110 3990 8170 4030
rect 8210 3990 8230 4030
rect 8050 3970 8230 3990
rect 8370 4330 8450 4520
rect 8370 4290 8390 4330
rect 8430 4290 8450 4330
rect 8370 4230 8450 4290
rect 8370 4190 8390 4230
rect 8430 4190 8450 4230
rect 8370 4130 8450 4190
rect 8370 4090 8390 4130
rect 8430 4090 8450 4130
rect 8370 4030 8450 4090
rect 8370 3990 8390 4030
rect 8430 3990 8450 4030
rect 8370 3970 8450 3990
rect 8590 4330 8670 4350
rect 8590 4290 8610 4330
rect 8650 4290 8670 4330
rect 8590 4230 8670 4290
rect 8590 4190 8610 4230
rect 8650 4190 8670 4230
rect 8590 4130 8670 4190
rect 8590 4090 8610 4130
rect 8650 4090 8670 4130
rect 8590 4030 8670 4090
rect 8590 3990 8610 4030
rect 8650 3990 8670 4030
rect 6870 3920 6950 3940
rect 8590 3930 8670 3990
rect 8810 4330 8890 4520
rect 8810 4290 8830 4330
rect 8870 4290 8890 4330
rect 8810 4230 8890 4290
rect 8810 4190 8830 4230
rect 8870 4190 8890 4230
rect 8810 4130 8890 4190
rect 8810 4090 8830 4130
rect 8870 4090 8890 4130
rect 8810 4030 8890 4090
rect 8810 3990 8830 4030
rect 8870 3990 8890 4030
rect 8810 3970 8890 3990
rect 9030 4330 9110 4350
rect 9030 4290 9050 4330
rect 9090 4290 9110 4330
rect 9030 4230 9110 4290
rect 9030 4190 9050 4230
rect 9090 4190 9110 4230
rect 9030 4130 9110 4190
rect 9030 4090 9050 4130
rect 9090 4090 9110 4130
rect 9030 4030 9110 4090
rect 9030 3990 9050 4030
rect 9090 3990 9110 4030
rect 9030 3930 9110 3990
rect 9250 4330 9330 4520
rect 9570 4350 9650 4520
rect 9250 4290 9270 4330
rect 9310 4290 9330 4330
rect 9250 4230 9330 4290
rect 9250 4190 9270 4230
rect 9310 4190 9330 4230
rect 9250 4130 9330 4190
rect 9250 4090 9270 4130
rect 9310 4090 9330 4130
rect 9250 4030 9330 4090
rect 9250 3990 9270 4030
rect 9310 3990 9330 4030
rect 9250 3970 9330 3990
rect 9470 4330 9750 4350
rect 9470 4290 9490 4330
rect 9530 4290 9590 4330
rect 9630 4290 9690 4330
rect 9730 4290 9750 4330
rect 9470 4230 9750 4290
rect 9470 4190 9490 4230
rect 9530 4190 9590 4230
rect 9630 4190 9690 4230
rect 9730 4190 9750 4230
rect 9470 4130 9750 4190
rect 9470 4090 9490 4130
rect 9530 4090 9590 4130
rect 9630 4090 9690 4130
rect 9730 4090 9750 4130
rect 9470 4030 9750 4090
rect 9470 3990 9490 4030
rect 9530 3990 9590 4030
rect 9630 3990 9690 4030
rect 9730 3990 9750 4030
rect 9470 3970 9750 3990
rect 9890 4330 9970 4520
rect 9890 4290 9910 4330
rect 9950 4290 9970 4330
rect 9890 4230 9970 4290
rect 9890 4190 9910 4230
rect 9950 4190 9970 4230
rect 9890 4130 9970 4190
rect 9890 4090 9910 4130
rect 9950 4090 9970 4130
rect 9890 4030 9970 4090
rect 9890 3990 9910 4030
rect 9950 3990 9970 4030
rect 9890 3970 9970 3990
rect 10110 4330 10190 4350
rect 10110 4290 10130 4330
rect 10170 4290 10190 4330
rect 10110 4230 10190 4290
rect 10110 4190 10130 4230
rect 10170 4190 10190 4230
rect 10110 4130 10190 4190
rect 10110 4090 10130 4130
rect 10170 4090 10190 4130
rect 10110 4030 10190 4090
rect 10110 3990 10130 4030
rect 10170 3990 10190 4030
rect 1900 3760 2000 3780
rect 1900 3700 1920 3760
rect 1980 3750 2000 3760
rect 2160 3750 2200 3920
rect 2900 3750 2940 3920
rect 3060 3750 3100 3920
rect 3800 3750 3840 3920
rect 4060 3750 4100 3920
rect 4140 3860 4220 3880
rect 4140 3820 4160 3860
rect 4200 3820 4220 3860
rect 4140 3800 4220 3820
rect 4320 3750 4360 3920
rect 4540 3750 4580 3920
rect 4870 3750 4910 3920
rect 5300 3750 5340 3920
rect 5690 3750 5730 3920
rect 6080 3750 6120 3920
rect 6760 3750 6800 3920
rect 8460 3880 8540 3900
rect 8460 3840 8480 3880
rect 8520 3840 8540 3880
rect 8460 3820 8540 3840
rect 8590 3850 9110 3930
rect 9570 3910 9650 3970
rect 9570 3870 9590 3910
rect 9630 3870 9650 3910
rect 10110 3930 10190 3990
rect 10330 4330 10410 4520
rect 10330 4290 10350 4330
rect 10390 4290 10410 4330
rect 10330 4230 10410 4290
rect 10330 4190 10350 4230
rect 10390 4190 10410 4230
rect 10330 4130 10410 4190
rect 10330 4090 10350 4130
rect 10390 4090 10410 4130
rect 10330 4030 10410 4090
rect 10330 3990 10350 4030
rect 10390 3990 10410 4030
rect 10330 3970 10410 3990
rect 10550 4330 10630 4350
rect 10550 4290 10570 4330
rect 10610 4290 10630 4330
rect 10550 4230 10630 4290
rect 10550 4190 10570 4230
rect 10610 4190 10630 4230
rect 10550 4130 10630 4190
rect 10550 4090 10570 4130
rect 10610 4090 10630 4130
rect 10550 4030 10630 4090
rect 10550 3990 10570 4030
rect 10610 3990 10630 4030
rect 10550 3930 10630 3990
rect 10770 4330 10850 4520
rect 10770 4290 10790 4330
rect 10830 4290 10850 4330
rect 10770 4230 10850 4290
rect 10770 4190 10790 4230
rect 10830 4190 10850 4230
rect 10770 4130 10850 4190
rect 10770 4090 10790 4130
rect 10830 4090 10850 4130
rect 10770 4030 10850 4090
rect 10770 3990 10790 4030
rect 10830 3990 10850 4030
rect 10770 3970 10850 3990
rect 10990 4450 11070 4520
rect 10990 4410 11010 4450
rect 11050 4410 11070 4450
rect 10990 4350 11070 4410
rect 10990 4330 11170 4350
rect 10990 4290 11010 4330
rect 11050 4290 11110 4330
rect 11150 4290 11170 4330
rect 10990 4230 11170 4290
rect 10990 4190 11010 4230
rect 11050 4190 11110 4230
rect 11150 4190 11170 4230
rect 10990 4130 11170 4190
rect 10990 4090 11010 4130
rect 11050 4090 11110 4130
rect 11150 4090 11170 4130
rect 10990 4030 11170 4090
rect 10990 3990 11010 4030
rect 11050 3990 11110 4030
rect 11150 3990 11170 4030
rect 10990 3970 11170 3990
rect 9570 3850 9650 3870
rect 9980 3880 10060 3900
rect 8590 3790 8670 3850
rect 7200 3760 7300 3790
rect 7200 3750 7230 3760
rect 1980 3710 2080 3750
rect 2120 3710 2180 3750
rect 2220 3710 2280 3750
rect 2320 3710 2380 3750
rect 2420 3710 2480 3750
rect 2520 3710 2580 3750
rect 2620 3710 2680 3750
rect 2720 3710 2780 3750
rect 2820 3710 2880 3750
rect 2920 3710 2980 3750
rect 3020 3710 3080 3750
rect 3120 3710 3180 3750
rect 3220 3710 3280 3750
rect 3320 3710 3380 3750
rect 3420 3710 3480 3750
rect 3520 3710 3580 3750
rect 3620 3710 3680 3750
rect 3720 3710 3780 3750
rect 3820 3710 3880 3750
rect 3920 3710 3980 3750
rect 4020 3710 4080 3750
rect 4120 3710 4180 3750
rect 4220 3710 4280 3750
rect 4320 3710 4380 3750
rect 4420 3710 4480 3750
rect 4520 3710 4580 3750
rect 4620 3710 4680 3750
rect 4720 3710 4780 3750
rect 4820 3710 4880 3750
rect 4920 3710 4980 3750
rect 5020 3710 5080 3750
rect 5120 3710 5180 3750
rect 5220 3710 5280 3750
rect 5320 3710 5380 3750
rect 5420 3710 5480 3750
rect 5520 3710 5580 3750
rect 5620 3710 5680 3750
rect 5720 3710 5780 3750
rect 5820 3710 5880 3750
rect 5920 3710 5980 3750
rect 6020 3710 6080 3750
rect 6120 3710 6180 3750
rect 6220 3710 6280 3750
rect 6320 3710 6380 3750
rect 6420 3710 6480 3750
rect 6520 3710 6580 3750
rect 6620 3710 6680 3750
rect 6720 3710 6780 3750
rect 6820 3710 6880 3750
rect 6920 3710 6980 3750
rect 7020 3710 7080 3750
rect 7120 3720 7230 3750
rect 7270 3720 7300 3760
rect 8590 3750 8610 3790
rect 8650 3750 8670 3790
rect 8590 3730 8670 3750
rect 7120 3710 7300 3720
rect 1980 3700 2000 3710
rect 1900 3680 2000 3700
rect 2160 3540 2200 3710
rect 2590 3640 2670 3660
rect 2590 3600 2610 3640
rect 2650 3600 2670 3640
rect 2590 3580 2670 3600
rect 2590 3540 2630 3580
rect 2900 3540 2940 3710
rect 3060 3540 3100 3710
rect 3800 3540 3840 3710
rect 4200 3540 4240 3710
rect 4530 3540 4570 3710
rect 4860 3540 4900 3710
rect 5300 3540 5340 3710
rect 5710 3640 5790 3660
rect 5710 3600 5730 3640
rect 5770 3600 5790 3640
rect 5710 3580 5790 3600
rect 6080 3540 6120 3710
rect 7200 3690 7300 3710
rect 9030 3700 9110 3850
rect 9980 3840 10000 3880
rect 10040 3840 10060 3880
rect 10110 3850 10630 3930
rect 11350 3910 11460 3930
rect 11350 3900 11370 3910
rect 9980 3820 10060 3840
rect 10550 3710 10630 3850
rect 10680 3880 11370 3900
rect 10680 3840 10700 3880
rect 10740 3840 11370 3880
rect 11440 3840 11460 3910
rect 10680 3820 11460 3840
rect 11180 3710 11260 3730
rect 6360 3630 6720 3670
rect 6360 3540 6400 3630
rect 6640 3610 6720 3630
rect 9030 3620 9550 3700
rect 6640 3570 6660 3610
rect 6700 3570 6720 3610
rect 6640 3550 6720 3570
rect 8390 3610 8470 3620
rect 8390 3560 8410 3610
rect 8450 3560 8470 3610
rect 2070 3520 2210 3540
rect 2070 3480 2080 3520
rect 2120 3480 2160 3520
rect 2200 3480 2210 3520
rect 2070 3420 2210 3480
rect 2070 3380 2080 3420
rect 2120 3380 2160 3420
rect 2200 3380 2210 3420
rect 2070 3320 2210 3380
rect 2070 3280 2080 3320
rect 2120 3280 2160 3320
rect 2200 3280 2210 3320
rect 2070 3220 2210 3280
rect 2070 3180 2080 3220
rect 2120 3180 2160 3220
rect 2200 3180 2210 3220
rect 2070 3160 2210 3180
rect 2260 3520 2320 3540
rect 2260 3480 2270 3520
rect 2310 3480 2320 3520
rect 2260 3420 2320 3480
rect 2260 3380 2270 3420
rect 2310 3380 2320 3420
rect 2260 3320 2320 3380
rect 2260 3280 2270 3320
rect 2310 3280 2320 3320
rect 2260 3220 2320 3280
rect 2260 3180 2270 3220
rect 2310 3180 2320 3220
rect 2260 3160 2320 3180
rect 2370 3520 2550 3540
rect 2370 3480 2380 3520
rect 2420 3490 2490 3520
rect 2420 3480 2430 3490
rect 2370 3420 2430 3480
rect 2470 3480 2490 3490
rect 2530 3480 2550 3520
rect 2470 3460 2550 3480
rect 2590 3520 2730 3540
rect 2590 3500 2680 3520
rect 2370 3380 2380 3420
rect 2420 3380 2430 3420
rect 2370 3320 2430 3380
rect 2370 3280 2380 3320
rect 2420 3280 2430 3320
rect 2370 3220 2430 3280
rect 2370 3180 2380 3220
rect 2420 3180 2430 3220
rect 2370 3160 2430 3180
rect 2380 3120 2420 3160
rect 2260 3080 2420 3120
rect 2020 3030 2100 3050
rect 2020 2990 2040 3030
rect 2080 2990 2100 3030
rect 2020 2970 2100 2990
rect 2260 2920 2300 3080
rect 2590 3040 2630 3500
rect 2670 3480 2680 3500
rect 2720 3480 2730 3520
rect 2670 3420 2730 3480
rect 2670 3380 2680 3420
rect 2720 3380 2730 3420
rect 2670 3320 2730 3380
rect 2670 3280 2680 3320
rect 2720 3280 2730 3320
rect 2670 3220 2730 3280
rect 2670 3180 2680 3220
rect 2720 3180 2730 3220
rect 2670 3160 2730 3180
rect 2780 3520 2840 3540
rect 2780 3480 2790 3520
rect 2830 3480 2840 3520
rect 2780 3420 2840 3480
rect 2780 3380 2790 3420
rect 2830 3380 2840 3420
rect 2780 3320 2840 3380
rect 2780 3280 2790 3320
rect 2830 3280 2840 3320
rect 2780 3220 2840 3280
rect 2780 3180 2790 3220
rect 2830 3180 2840 3220
rect 2780 3160 2840 3180
rect 2890 3520 3110 3540
rect 2890 3480 2900 3520
rect 2940 3480 2980 3520
rect 3020 3480 3060 3520
rect 3100 3480 3110 3520
rect 2890 3420 3110 3480
rect 2890 3380 2900 3420
rect 2940 3380 2980 3420
rect 3020 3380 3060 3420
rect 3100 3380 3110 3420
rect 2890 3320 3110 3380
rect 2890 3280 2900 3320
rect 2940 3280 2980 3320
rect 3020 3280 3060 3320
rect 3100 3280 3110 3320
rect 2890 3220 3110 3280
rect 2890 3180 2900 3220
rect 2940 3180 2980 3220
rect 3020 3180 3060 3220
rect 3100 3180 3110 3220
rect 2890 3160 3110 3180
rect 3160 3520 3220 3540
rect 3160 3480 3170 3520
rect 3210 3480 3220 3520
rect 3160 3420 3220 3480
rect 3160 3380 3170 3420
rect 3210 3380 3220 3420
rect 3160 3320 3220 3380
rect 3160 3280 3170 3320
rect 3210 3280 3220 3320
rect 3160 3220 3220 3280
rect 3160 3180 3170 3220
rect 3210 3180 3220 3220
rect 3160 3160 3220 3180
rect 3270 3520 3450 3540
rect 3270 3480 3280 3520
rect 3320 3490 3390 3520
rect 3320 3480 3330 3490
rect 3270 3420 3330 3480
rect 3370 3480 3390 3490
rect 3430 3480 3450 3520
rect 3370 3460 3450 3480
rect 3490 3520 3630 3540
rect 3490 3500 3580 3520
rect 3270 3380 3280 3420
rect 3320 3380 3330 3420
rect 3270 3320 3330 3380
rect 3270 3280 3280 3320
rect 3320 3280 3330 3320
rect 3270 3220 3330 3280
rect 3270 3180 3280 3220
rect 3320 3180 3330 3220
rect 3270 3160 3330 3180
rect 2680 3120 2720 3160
rect 3280 3120 3320 3160
rect 2680 3080 2830 3120
rect 2350 3020 2630 3040
rect 2350 2980 2370 3020
rect 2410 3000 2630 3020
rect 2410 2980 2430 3000
rect 2350 2960 2430 2980
rect 2790 2920 2830 3080
rect 2870 3100 3320 3120
rect 2870 3060 2890 3100
rect 2930 3080 3320 3100
rect 2930 3060 2950 3080
rect 2870 3040 2950 3060
rect 3160 2920 3200 3080
rect 3490 3040 3530 3500
rect 3570 3480 3580 3500
rect 3620 3480 3630 3520
rect 3570 3420 3630 3480
rect 3570 3380 3580 3420
rect 3620 3380 3630 3420
rect 3570 3320 3630 3380
rect 3570 3280 3580 3320
rect 3620 3280 3630 3320
rect 3570 3220 3630 3280
rect 3570 3180 3580 3220
rect 3620 3180 3630 3220
rect 3570 3160 3630 3180
rect 3680 3520 3740 3540
rect 3680 3480 3690 3520
rect 3730 3480 3740 3520
rect 3680 3420 3740 3480
rect 3680 3380 3690 3420
rect 3730 3380 3740 3420
rect 3680 3320 3740 3380
rect 3680 3280 3690 3320
rect 3730 3280 3740 3320
rect 3680 3220 3740 3280
rect 3680 3180 3690 3220
rect 3730 3180 3740 3220
rect 3680 3160 3740 3180
rect 3790 3520 3930 3540
rect 3790 3480 3800 3520
rect 3840 3480 3880 3520
rect 3920 3480 3930 3520
rect 3790 3420 3930 3480
rect 3790 3380 3800 3420
rect 3840 3380 3880 3420
rect 3920 3380 3930 3420
rect 3790 3320 3930 3380
rect 3790 3280 3800 3320
rect 3840 3280 3880 3320
rect 3920 3280 3930 3320
rect 3790 3220 3930 3280
rect 3790 3180 3800 3220
rect 3840 3180 3880 3220
rect 3920 3180 3930 3220
rect 3790 3160 3930 3180
rect 4080 3520 4140 3540
rect 4080 3480 4090 3520
rect 4130 3480 4140 3520
rect 4080 3420 4140 3480
rect 4080 3380 4090 3420
rect 4130 3380 4140 3420
rect 4080 3320 4140 3380
rect 4080 3280 4090 3320
rect 4130 3280 4140 3320
rect 4080 3220 4140 3280
rect 4080 3180 4090 3220
rect 4130 3180 4140 3220
rect 4080 3160 4140 3180
rect 4190 3520 4330 3540
rect 4190 3480 4200 3520
rect 4240 3480 4280 3520
rect 4320 3480 4330 3520
rect 4190 3420 4330 3480
rect 4190 3380 4200 3420
rect 4240 3380 4280 3420
rect 4320 3380 4330 3420
rect 4190 3320 4330 3380
rect 4190 3280 4200 3320
rect 4240 3280 4280 3320
rect 4320 3280 4330 3320
rect 4190 3220 4330 3280
rect 4190 3180 4200 3220
rect 4240 3180 4280 3220
rect 4320 3180 4330 3220
rect 4190 3160 4330 3180
rect 4410 3520 4470 3540
rect 4410 3480 4420 3520
rect 4460 3480 4470 3520
rect 4410 3420 4470 3480
rect 4410 3380 4420 3420
rect 4460 3380 4470 3420
rect 4410 3320 4470 3380
rect 4410 3280 4420 3320
rect 4460 3280 4470 3320
rect 4410 3220 4470 3280
rect 4410 3180 4420 3220
rect 4460 3180 4470 3220
rect 4410 3160 4470 3180
rect 4520 3520 4660 3540
rect 4520 3480 4530 3520
rect 4570 3480 4610 3520
rect 4650 3480 4660 3520
rect 4520 3420 4660 3480
rect 4520 3380 4530 3420
rect 4570 3380 4610 3420
rect 4650 3380 4660 3420
rect 4520 3320 4660 3380
rect 4520 3280 4530 3320
rect 4570 3280 4610 3320
rect 4650 3280 4660 3320
rect 4520 3220 4660 3280
rect 4520 3180 4530 3220
rect 4570 3180 4610 3220
rect 4650 3180 4660 3220
rect 4520 3160 4660 3180
rect 4740 3520 4800 3540
rect 4740 3480 4750 3520
rect 4790 3480 4800 3520
rect 4740 3420 4800 3480
rect 4740 3380 4750 3420
rect 4790 3380 4800 3420
rect 4740 3320 4800 3380
rect 4740 3280 4750 3320
rect 4790 3280 4800 3320
rect 4740 3220 4800 3280
rect 4740 3180 4750 3220
rect 4790 3180 4800 3220
rect 4740 3160 4800 3180
rect 4850 3520 4990 3540
rect 4850 3480 4860 3520
rect 4900 3480 4940 3520
rect 4980 3480 4990 3520
rect 4850 3420 4990 3480
rect 4850 3380 4860 3420
rect 4900 3380 4940 3420
rect 4980 3380 4990 3420
rect 4850 3320 4990 3380
rect 4850 3280 4860 3320
rect 4900 3280 4940 3320
rect 4980 3280 4990 3320
rect 4850 3220 4990 3280
rect 4850 3180 4860 3220
rect 4900 3180 4940 3220
rect 4980 3180 4990 3220
rect 4850 3160 4990 3180
rect 5180 3520 5360 3540
rect 5180 3480 5200 3520
rect 5240 3480 5300 3520
rect 5340 3480 5360 3520
rect 5180 3420 5360 3480
rect 5180 3380 5200 3420
rect 5240 3380 5300 3420
rect 5340 3380 5360 3420
rect 5180 3320 5360 3380
rect 5180 3280 5200 3320
rect 5240 3280 5300 3320
rect 5340 3280 5360 3320
rect 5180 3220 5360 3280
rect 5180 3180 5200 3220
rect 5240 3180 5300 3220
rect 5340 3180 5360 3220
rect 5180 3160 5360 3180
rect 5410 3520 5490 3540
rect 5410 3480 5430 3520
rect 5470 3480 5490 3520
rect 5410 3420 5490 3480
rect 5410 3380 5430 3420
rect 5470 3380 5490 3420
rect 5410 3320 5490 3380
rect 5410 3280 5430 3320
rect 5470 3280 5490 3320
rect 5410 3220 5490 3280
rect 5410 3180 5430 3220
rect 5470 3180 5490 3220
rect 5410 3160 5490 3180
rect 5670 3520 5750 3540
rect 5670 3480 5690 3520
rect 5730 3480 5750 3520
rect 5670 3420 5750 3480
rect 5670 3380 5690 3420
rect 5730 3380 5750 3420
rect 5670 3320 5750 3380
rect 5670 3280 5690 3320
rect 5730 3280 5750 3320
rect 5670 3220 5750 3280
rect 5670 3180 5690 3220
rect 5730 3180 5750 3220
rect 5670 3160 5750 3180
rect 5800 3520 5880 3540
rect 5800 3480 5820 3520
rect 5860 3480 5880 3520
rect 5800 3420 5880 3480
rect 5800 3380 5820 3420
rect 5860 3380 5880 3420
rect 5800 3320 5880 3380
rect 5800 3280 5820 3320
rect 5860 3280 5880 3320
rect 5800 3220 5880 3280
rect 5800 3180 5820 3220
rect 5860 3180 5880 3220
rect 5800 3160 5880 3180
rect 5960 3520 6140 3540
rect 5960 3480 5980 3520
rect 6020 3480 6080 3520
rect 6120 3480 6140 3520
rect 5960 3420 6140 3480
rect 5960 3380 5980 3420
rect 6020 3380 6080 3420
rect 6120 3380 6140 3420
rect 5960 3320 6140 3380
rect 5960 3280 5980 3320
rect 6020 3280 6080 3320
rect 6120 3280 6140 3320
rect 5960 3220 6140 3280
rect 5960 3180 5980 3220
rect 6020 3180 6080 3220
rect 6120 3180 6140 3220
rect 5960 3160 6140 3180
rect 6190 3520 6270 3540
rect 6190 3480 6210 3520
rect 6250 3480 6270 3520
rect 6190 3420 6270 3480
rect 6190 3380 6210 3420
rect 6250 3380 6270 3420
rect 6190 3320 6270 3380
rect 6190 3280 6210 3320
rect 6250 3280 6270 3320
rect 6190 3220 6270 3280
rect 6190 3180 6210 3220
rect 6250 3180 6270 3220
rect 6190 3160 6270 3180
rect 6350 3520 6430 3540
rect 6350 3480 6370 3520
rect 6410 3480 6430 3520
rect 6350 3420 6430 3480
rect 6350 3380 6370 3420
rect 6410 3380 6430 3420
rect 6350 3320 6430 3380
rect 6350 3280 6370 3320
rect 6410 3280 6430 3320
rect 6350 3220 6430 3280
rect 6350 3180 6370 3220
rect 6410 3180 6430 3220
rect 6350 3160 6430 3180
rect 6480 3520 6560 3540
rect 6480 3480 6500 3520
rect 6540 3480 6560 3520
rect 6480 3420 6560 3480
rect 6480 3380 6500 3420
rect 6540 3380 6560 3420
rect 6480 3320 6560 3380
rect 6480 3280 6500 3320
rect 6540 3280 6560 3320
rect 6480 3220 6560 3280
rect 6480 3180 6500 3220
rect 6540 3180 6560 3220
rect 6480 3160 6560 3180
rect 7850 3350 8030 3370
rect 7850 3310 7870 3350
rect 7910 3310 7970 3350
rect 8010 3310 8030 3350
rect 7850 3250 8030 3310
rect 7850 3210 7870 3250
rect 7910 3210 7970 3250
rect 8010 3210 8030 3250
rect 3580 3120 3620 3160
rect 3580 3080 3730 3120
rect 4080 3090 4120 3160
rect 4410 3090 4450 3160
rect 4740 3090 4780 3160
rect 5430 3120 5470 3160
rect 5690 3120 5730 3160
rect 3250 3020 3530 3040
rect 3250 2980 3270 3020
rect 3310 3000 3530 3020
rect 3310 2980 3330 3000
rect 3250 2960 3330 2980
rect 3690 2920 3730 3080
rect 3860 3070 3940 3090
rect 3860 3030 3880 3070
rect 3920 3030 3940 3070
rect 3860 3010 3940 3030
rect 4020 3070 4120 3090
rect 4020 3030 4040 3070
rect 4080 3030 4120 3070
rect 4020 3010 4120 3030
rect 4350 3070 4450 3090
rect 4350 3030 4370 3070
rect 4410 3030 4450 3070
rect 4350 3010 4450 3030
rect 4680 3070 4780 3090
rect 4680 3030 4700 3070
rect 4740 3030 4780 3070
rect 4680 3010 4780 3030
rect 4940 3070 5020 3090
rect 5430 3080 5730 3120
rect 4940 3030 4960 3070
rect 5000 3030 5020 3070
rect 4940 3010 5020 3030
rect 5140 3060 5220 3080
rect 5140 3020 5160 3060
rect 5200 3020 5220 3060
rect 4080 2920 4120 3010
rect 4410 2920 4450 3010
rect 4740 2920 4780 3010
rect 5140 3000 5220 3020
rect 5430 2920 5470 3080
rect 5690 2920 5730 3080
rect 5820 3110 5860 3160
rect 5820 3090 5920 3110
rect 5820 3050 5860 3090
rect 5900 3050 5920 3090
rect 5820 3030 5920 3050
rect 5820 2920 5860 3030
rect 6230 3020 6270 3160
rect 6230 3010 6310 3020
rect 6230 2970 6250 3010
rect 6290 2970 6310 3010
rect 6230 2950 6310 2970
rect 6230 2920 6270 2950
rect 6370 2920 6410 3160
rect 6500 3040 6540 3160
rect 7850 3150 8030 3210
rect 7850 3110 7870 3150
rect 7910 3110 7970 3150
rect 8010 3110 8030 3150
rect 6890 3070 6970 3090
rect 6890 3040 6910 3070
rect 6500 3030 6910 3040
rect 6950 3030 6970 3070
rect 6500 3010 6970 3030
rect 7850 3050 8030 3110
rect 7850 3010 7870 3050
rect 7910 3010 7970 3050
rect 8010 3010 8030 3050
rect 6500 3000 6930 3010
rect 6500 2920 6540 3000
rect 6890 2920 6930 3000
rect 7850 2990 8030 3010
rect 7950 2930 8030 2990
rect 2070 2900 2210 2920
rect 2070 2860 2080 2900
rect 2120 2860 2160 2900
rect 2200 2860 2210 2900
rect 2070 2800 2210 2860
rect 2070 2760 2080 2800
rect 2120 2760 2160 2800
rect 2200 2760 2210 2800
rect 2070 2740 2210 2760
rect 2260 2900 2320 2920
rect 2260 2860 2270 2900
rect 2310 2860 2320 2900
rect 2260 2800 2320 2860
rect 2260 2760 2270 2800
rect 2310 2760 2320 2800
rect 2260 2740 2320 2760
rect 2370 2900 2430 2920
rect 2370 2860 2380 2900
rect 2420 2860 2430 2900
rect 2370 2800 2430 2860
rect 2370 2760 2380 2800
rect 2420 2760 2430 2800
rect 2370 2740 2430 2760
rect 2670 2900 2730 2920
rect 2670 2860 2680 2900
rect 2720 2860 2730 2900
rect 2670 2800 2730 2860
rect 2670 2760 2680 2800
rect 2720 2760 2730 2800
rect 2670 2740 2730 2760
rect 2780 2900 2840 2920
rect 2780 2860 2790 2900
rect 2830 2860 2840 2900
rect 2780 2800 2840 2860
rect 2780 2760 2790 2800
rect 2830 2760 2840 2800
rect 2780 2740 2840 2760
rect 2890 2900 3110 2920
rect 2890 2860 2900 2900
rect 2940 2860 2980 2900
rect 3020 2860 3060 2900
rect 3100 2860 3110 2900
rect 2890 2800 3110 2860
rect 2890 2760 2900 2800
rect 2940 2760 2980 2800
rect 3020 2760 3060 2800
rect 3100 2760 3110 2800
rect 2890 2740 3110 2760
rect 3160 2900 3220 2920
rect 3160 2860 3170 2900
rect 3210 2860 3220 2900
rect 3160 2800 3220 2860
rect 3160 2760 3170 2800
rect 3210 2760 3220 2800
rect 3160 2740 3220 2760
rect 3270 2900 3330 2920
rect 3270 2860 3280 2900
rect 3320 2860 3330 2900
rect 3270 2800 3330 2860
rect 3270 2760 3280 2800
rect 3320 2760 3330 2800
rect 3270 2740 3330 2760
rect 3570 2900 3630 2920
rect 3570 2860 3580 2900
rect 3620 2860 3630 2900
rect 3570 2800 3630 2860
rect 3570 2760 3580 2800
rect 3620 2760 3630 2800
rect 3570 2740 3630 2760
rect 3680 2900 3740 2920
rect 3680 2860 3690 2900
rect 3730 2860 3740 2900
rect 3680 2800 3740 2860
rect 3680 2760 3690 2800
rect 3730 2760 3740 2800
rect 3680 2740 3740 2760
rect 3790 2900 3930 2920
rect 3790 2860 3800 2900
rect 3840 2860 3880 2900
rect 3920 2860 3930 2900
rect 3790 2800 3930 2860
rect 3790 2760 3800 2800
rect 3840 2760 3880 2800
rect 3920 2760 3930 2800
rect 3790 2740 3930 2760
rect 4080 2900 4140 2920
rect 4080 2860 4090 2900
rect 4130 2860 4140 2900
rect 4080 2800 4140 2860
rect 4080 2760 4090 2800
rect 4130 2760 4140 2800
rect 4080 2740 4140 2760
rect 4190 2900 4330 2920
rect 4190 2860 4200 2900
rect 4240 2860 4280 2900
rect 4320 2860 4330 2900
rect 4190 2800 4330 2860
rect 4190 2760 4200 2800
rect 4240 2760 4280 2800
rect 4320 2760 4330 2800
rect 4190 2740 4330 2760
rect 4410 2900 4470 2920
rect 4410 2860 4420 2900
rect 4460 2860 4470 2900
rect 4410 2800 4470 2860
rect 4410 2760 4420 2800
rect 4460 2760 4470 2800
rect 4410 2740 4470 2760
rect 4520 2900 4660 2920
rect 4520 2860 4530 2900
rect 4570 2860 4610 2900
rect 4650 2860 4660 2900
rect 4520 2800 4660 2860
rect 4520 2760 4530 2800
rect 4570 2760 4610 2800
rect 4650 2760 4660 2800
rect 4520 2740 4660 2760
rect 4740 2900 4800 2920
rect 4740 2860 4750 2900
rect 4790 2860 4800 2900
rect 4740 2800 4800 2860
rect 4740 2760 4750 2800
rect 4790 2760 4800 2800
rect 4740 2740 4800 2760
rect 4850 2900 4990 2920
rect 4850 2860 4860 2900
rect 4900 2860 4940 2900
rect 4980 2860 4990 2900
rect 4850 2800 4990 2860
rect 4850 2760 4860 2800
rect 4900 2760 4940 2800
rect 4980 2760 4990 2800
rect 4850 2740 4990 2760
rect 5180 2900 5360 2920
rect 5180 2860 5200 2900
rect 5240 2860 5300 2900
rect 5340 2860 5360 2900
rect 5180 2800 5360 2860
rect 5180 2760 5200 2800
rect 5240 2760 5300 2800
rect 5340 2760 5360 2800
rect 5180 2740 5360 2760
rect 5410 2900 5490 2920
rect 5410 2860 5430 2900
rect 5470 2860 5490 2900
rect 5410 2800 5490 2860
rect 5410 2760 5430 2800
rect 5470 2760 5490 2800
rect 5410 2740 5490 2760
rect 5670 2900 5750 2920
rect 5670 2860 5690 2900
rect 5730 2860 5750 2900
rect 5670 2800 5750 2860
rect 5670 2760 5690 2800
rect 5730 2760 5750 2800
rect 5670 2740 5750 2760
rect 5800 2900 5880 2920
rect 5800 2860 5820 2900
rect 5860 2860 5880 2900
rect 5800 2800 5880 2860
rect 5800 2760 5820 2800
rect 5860 2760 5880 2800
rect 5800 2740 5880 2760
rect 5960 2900 6140 2920
rect 5960 2860 5980 2900
rect 6020 2860 6080 2900
rect 6120 2860 6140 2900
rect 5960 2800 6140 2860
rect 5960 2760 5980 2800
rect 6020 2760 6080 2800
rect 6120 2760 6140 2800
rect 5960 2740 6140 2760
rect 6190 2900 6270 2920
rect 6190 2860 6210 2900
rect 6250 2860 6270 2900
rect 6190 2800 6270 2860
rect 6190 2760 6210 2800
rect 6250 2760 6270 2800
rect 6190 2740 6270 2760
rect 6350 2900 6430 2920
rect 6350 2860 6370 2900
rect 6410 2860 6430 2900
rect 6350 2800 6430 2860
rect 6350 2760 6370 2800
rect 6410 2760 6430 2800
rect 6350 2740 6430 2760
rect 6480 2900 6560 2920
rect 6480 2860 6500 2900
rect 6540 2860 6560 2900
rect 6480 2800 6560 2860
rect 6480 2760 6500 2800
rect 6540 2760 6560 2800
rect 6480 2740 6560 2760
rect 6640 2900 6820 2920
rect 6640 2860 6660 2900
rect 6700 2860 6760 2900
rect 6800 2860 6820 2900
rect 6640 2800 6820 2860
rect 6640 2760 6660 2800
rect 6700 2760 6760 2800
rect 6800 2760 6820 2800
rect 6640 2740 6820 2760
rect 6870 2900 6950 2920
rect 6870 2860 6890 2900
rect 6930 2860 6950 2900
rect 6870 2800 6950 2860
rect 7950 2890 7970 2930
rect 8010 2890 8030 2930
rect 7950 2840 8030 2890
rect 8170 3350 8250 3370
rect 8170 3310 8190 3350
rect 8230 3310 8250 3350
rect 8170 3250 8250 3310
rect 8170 3210 8190 3250
rect 8230 3210 8250 3250
rect 8170 3150 8250 3210
rect 8170 3110 8190 3150
rect 8230 3110 8250 3150
rect 8170 3050 8250 3110
rect 8170 3010 8190 3050
rect 8230 3010 8250 3050
rect 8170 2840 8250 3010
rect 8390 3350 8470 3560
rect 8930 3470 9010 3490
rect 8930 3430 8950 3470
rect 8990 3430 9010 3470
rect 8930 3370 9010 3430
rect 8390 3310 8410 3350
rect 8450 3310 8470 3350
rect 8390 3250 8470 3310
rect 8390 3210 8410 3250
rect 8450 3210 8470 3250
rect 8390 3150 8470 3210
rect 8390 3110 8410 3150
rect 8450 3110 8470 3150
rect 8390 3050 8470 3110
rect 8390 3010 8410 3050
rect 8450 3010 8470 3050
rect 8390 2990 8470 3010
rect 8610 3350 8690 3370
rect 8610 3310 8630 3350
rect 8670 3310 8690 3350
rect 8610 3250 8690 3310
rect 8610 3210 8630 3250
rect 8670 3210 8690 3250
rect 8610 3150 8690 3210
rect 8610 3110 8630 3150
rect 8670 3110 8690 3150
rect 8610 3050 8690 3110
rect 8610 3010 8630 3050
rect 8670 3010 8690 3050
rect 8610 2840 8690 3010
rect 8830 3350 9110 3370
rect 8830 3310 8850 3350
rect 8890 3310 8950 3350
rect 8990 3310 9050 3350
rect 9090 3310 9110 3350
rect 8830 3250 9110 3310
rect 8830 3210 8850 3250
rect 8890 3210 8950 3250
rect 8990 3210 9050 3250
rect 9090 3210 9110 3250
rect 8830 3150 9110 3210
rect 8830 3110 8850 3150
rect 8890 3110 8950 3150
rect 8990 3110 9050 3150
rect 9090 3110 9110 3150
rect 8830 3050 9110 3110
rect 8830 3010 8850 3050
rect 8890 3010 8950 3050
rect 8990 3010 9050 3050
rect 9090 3010 9110 3050
rect 8830 2990 9110 3010
rect 9250 3350 9330 3370
rect 9250 3310 9270 3350
rect 9310 3310 9330 3350
rect 9250 3250 9330 3310
rect 9250 3210 9270 3250
rect 9310 3210 9330 3250
rect 9250 3150 9330 3210
rect 9250 3110 9270 3150
rect 9310 3110 9330 3150
rect 9250 3050 9330 3110
rect 9250 3010 9270 3050
rect 9310 3010 9330 3050
rect 8930 2840 9010 2990
rect 9250 2840 9330 3010
rect 9470 3350 9550 3620
rect 10550 3670 11200 3710
rect 11240 3670 11260 3710
rect 10550 3630 11260 3670
rect 10420 3500 10500 3520
rect 10010 3470 10090 3490
rect 10010 3430 10030 3470
rect 10070 3430 10090 3470
rect 10420 3460 10440 3500
rect 10480 3460 10500 3500
rect 10420 3440 10500 3460
rect 10010 3370 10090 3430
rect 9470 3310 9490 3350
rect 9530 3310 9550 3350
rect 9470 3250 9550 3310
rect 9470 3210 9490 3250
rect 9530 3210 9550 3250
rect 9470 3150 9550 3210
rect 9470 3110 9490 3150
rect 9530 3110 9550 3150
rect 9470 3050 9550 3110
rect 9470 3010 9490 3050
rect 9530 3010 9550 3050
rect 9470 2990 9550 3010
rect 9690 3350 9770 3370
rect 9690 3310 9710 3350
rect 9750 3310 9770 3350
rect 9690 3250 9770 3310
rect 9690 3210 9710 3250
rect 9750 3210 9770 3250
rect 9690 3150 9770 3210
rect 9690 3110 9710 3150
rect 9750 3110 9770 3150
rect 9690 3050 9770 3110
rect 9690 3010 9710 3050
rect 9750 3010 9770 3050
rect 9690 2840 9770 3010
rect 9910 3350 10190 3370
rect 9910 3310 9930 3350
rect 9970 3310 10030 3350
rect 10070 3310 10130 3350
rect 10170 3310 10190 3350
rect 9910 3250 10190 3310
rect 9910 3210 9930 3250
rect 9970 3210 10030 3250
rect 10070 3210 10130 3250
rect 10170 3210 10190 3250
rect 9910 3150 10190 3210
rect 9910 3110 9930 3150
rect 9970 3110 10030 3150
rect 10070 3110 10130 3150
rect 10170 3110 10190 3150
rect 9910 3050 10190 3110
rect 9910 3010 9930 3050
rect 9970 3010 10030 3050
rect 10070 3010 10130 3050
rect 10170 3010 10190 3050
rect 9910 2990 10190 3010
rect 10330 3350 10410 3370
rect 10330 3310 10350 3350
rect 10390 3310 10410 3350
rect 10330 3250 10410 3310
rect 10330 3210 10350 3250
rect 10390 3210 10410 3250
rect 10330 3150 10410 3210
rect 10330 3110 10350 3150
rect 10390 3110 10410 3150
rect 10330 3050 10410 3110
rect 10330 3010 10350 3050
rect 10390 3010 10410 3050
rect 10010 2840 10090 2990
rect 10330 2840 10410 3010
rect 10550 3350 10630 3630
rect 10680 3500 11460 3520
rect 10680 3460 10700 3500
rect 10740 3460 11370 3500
rect 10680 3440 11370 3460
rect 11350 3430 11370 3440
rect 11440 3430 11460 3500
rect 11350 3410 11460 3430
rect 10550 3310 10570 3350
rect 10610 3310 10630 3350
rect 10550 3250 10630 3310
rect 10550 3210 10570 3250
rect 10610 3210 10630 3250
rect 10550 3150 10630 3210
rect 10550 3110 10570 3150
rect 10610 3110 10630 3150
rect 10550 3050 10630 3110
rect 10550 3010 10570 3050
rect 10610 3010 10630 3050
rect 10550 2990 10630 3010
rect 10770 3350 10850 3370
rect 10770 3310 10790 3350
rect 10830 3310 10850 3350
rect 10770 3250 10850 3310
rect 10770 3210 10790 3250
rect 10830 3210 10850 3250
rect 10770 3150 10850 3210
rect 10770 3110 10790 3150
rect 10830 3110 10850 3150
rect 10770 3050 10850 3110
rect 10770 3010 10790 3050
rect 10830 3010 10850 3050
rect 10770 2840 10850 3010
rect 10990 3350 11170 3370
rect 10990 3310 11010 3350
rect 11050 3310 11110 3350
rect 11150 3310 11170 3350
rect 10990 3250 11170 3310
rect 10990 3210 11010 3250
rect 11050 3210 11110 3250
rect 11150 3210 11170 3250
rect 10990 3150 11170 3210
rect 10990 3110 11010 3150
rect 11050 3110 11110 3150
rect 11150 3110 11170 3150
rect 10990 3050 11170 3110
rect 10990 3010 11010 3050
rect 11050 3010 11110 3050
rect 11150 3010 11170 3050
rect 10990 2990 11170 3010
rect 10990 2930 11070 2990
rect 10990 2890 11010 2930
rect 11050 2890 11070 2930
rect 10990 2840 11070 2890
rect 7850 2800 7910 2840
rect 7950 2800 8010 2840
rect 8050 2800 8110 2840
rect 8150 2800 8210 2840
rect 8250 2800 8310 2840
rect 8350 2800 8410 2840
rect 8450 2800 8510 2840
rect 8550 2800 8610 2840
rect 8650 2800 8710 2840
rect 8750 2800 8810 2840
rect 8850 2800 8910 2840
rect 8950 2800 9010 2840
rect 9050 2800 9110 2840
rect 9150 2800 9210 2840
rect 9250 2800 9310 2840
rect 9350 2800 9410 2840
rect 9450 2800 9510 2840
rect 9550 2800 9610 2840
rect 9650 2800 9710 2840
rect 9750 2800 9810 2840
rect 9850 2800 9910 2840
rect 9950 2800 10010 2840
rect 10050 2800 10110 2840
rect 10150 2800 10210 2840
rect 10250 2800 10310 2840
rect 10350 2800 10410 2840
rect 10450 2800 10510 2840
rect 10550 2800 10610 2840
rect 10650 2800 10710 2840
rect 10750 2800 10810 2840
rect 10850 2800 10910 2840
rect 10950 2800 11010 2840
rect 11050 2800 11070 2840
rect 6870 2760 6890 2800
rect 6930 2760 6950 2800
rect 6870 2740 6950 2760
rect 1720 2580 1820 2610
rect 1720 2540 1750 2580
rect 1790 2570 1820 2580
rect 2160 2570 2200 2740
rect 2380 2570 2420 2740
rect 2680 2570 2720 2740
rect 2910 2570 2950 2740
rect 3060 2570 3100 2740
rect 3280 2570 3320 2740
rect 3580 2570 3620 2740
rect 3800 2570 3840 2740
rect 4200 2570 4240 2740
rect 4530 2570 4570 2740
rect 4860 2570 4900 2740
rect 5300 2570 5340 2740
rect 5790 2680 5870 2700
rect 5790 2640 5810 2680
rect 5850 2640 5870 2680
rect 5790 2620 5870 2640
rect 6080 2570 6120 2740
rect 6430 2680 6510 2700
rect 6430 2640 6450 2680
rect 6490 2640 6510 2680
rect 6430 2620 6510 2640
rect 6760 2570 6800 2740
rect 17090 2730 17200 2750
rect 11700 2710 11810 2730
rect 11700 2640 11720 2710
rect 11790 2640 11810 2710
rect 17090 2660 17110 2730
rect 17180 2680 17200 2730
rect 17590 2730 17700 2750
rect 17590 2680 17610 2730
rect 17180 2660 17610 2680
rect 17680 2660 17700 2730
rect 17090 2650 17700 2660
rect 17090 2640 17380 2650
rect 11700 2620 11810 2640
rect 17350 2610 17380 2640
rect 17420 2640 17700 2650
rect 17420 2610 17450 2640
rect 17350 2580 17450 2610
rect 1790 2540 1880 2570
rect 1720 2530 1880 2540
rect 1920 2530 1980 2570
rect 2020 2530 2080 2570
rect 2120 2530 2180 2570
rect 2220 2530 2280 2570
rect 2320 2530 2380 2570
rect 2420 2530 2480 2570
rect 2520 2530 2580 2570
rect 2620 2530 2680 2570
rect 2720 2530 2780 2570
rect 2820 2530 2880 2570
rect 2920 2530 2980 2570
rect 3020 2530 3080 2570
rect 3120 2530 3180 2570
rect 3220 2530 3280 2570
rect 3320 2530 3380 2570
rect 3420 2530 3480 2570
rect 3520 2530 3580 2570
rect 3620 2530 3680 2570
rect 3720 2530 3780 2570
rect 3820 2530 3880 2570
rect 3920 2530 3980 2570
rect 4020 2530 4080 2570
rect 4120 2530 4180 2570
rect 4220 2530 4280 2570
rect 4320 2530 4380 2570
rect 4420 2530 4480 2570
rect 4520 2530 4580 2570
rect 4620 2530 4680 2570
rect 4720 2530 4780 2570
rect 4820 2530 4880 2570
rect 4920 2530 4980 2570
rect 5020 2530 5080 2570
rect 5120 2530 5180 2570
rect 5220 2530 5280 2570
rect 5320 2530 5380 2570
rect 5420 2530 5480 2570
rect 5520 2530 5580 2570
rect 5620 2530 5680 2570
rect 5720 2530 5780 2570
rect 5820 2530 5880 2570
rect 5920 2530 5980 2570
rect 6020 2530 6080 2570
rect 6120 2530 6180 2570
rect 6220 2530 6280 2570
rect 6320 2530 6380 2570
rect 6420 2530 6480 2570
rect 6520 2530 6580 2570
rect 6620 2530 6680 2570
rect 6720 2530 6780 2570
rect 6820 2530 6880 2570
rect 6920 2530 7040 2570
rect 1720 2510 1820 2530
rect 14410 2520 14510 2540
rect 14410 2460 14430 2520
rect 14490 2460 14510 2520
rect 14410 2440 14510 2460
rect 12170 2160 12270 2180
rect 17380 2160 17420 2580
rect 23100 2500 23180 2510
rect 23100 2450 23110 2500
rect 23160 2450 23180 2500
rect 23100 2440 23180 2450
rect 25532 2500 25612 2510
rect 25532 2450 25552 2500
rect 25602 2450 25612 2500
rect 25532 2440 25612 2450
rect 7140 2120 7200 2160
rect 7240 2120 7300 2160
rect 7340 2120 7400 2160
rect 7440 2120 7500 2160
rect 7540 2120 7600 2160
rect 7640 2120 7700 2160
rect 7740 2120 7800 2160
rect 7840 2120 7900 2160
rect 7940 2120 8000 2160
rect 8040 2120 8100 2160
rect 8140 2120 8200 2160
rect 8240 2120 8300 2160
rect 8340 2120 8400 2160
rect 8440 2120 8500 2160
rect 8540 2120 8600 2160
rect 8640 2120 8700 2160
rect 8740 2120 8800 2160
rect 8840 2120 8900 2160
rect 8940 2120 9000 2160
rect 9040 2120 9100 2160
rect 9140 2120 9200 2160
rect 9240 2120 9300 2160
rect 9340 2120 9400 2160
rect 9440 2120 9500 2160
rect 9540 2120 9600 2160
rect 9640 2120 9700 2160
rect 9740 2120 9800 2160
rect 9840 2120 9900 2160
rect 9940 2120 10000 2160
rect 10040 2120 10100 2160
rect 10140 2120 10200 2160
rect 10240 2120 10300 2160
rect 10340 2120 10400 2160
rect 10440 2120 10500 2160
rect 10540 2120 10600 2160
rect 10640 2120 10700 2160
rect 10740 2120 10800 2160
rect 10840 2120 10900 2160
rect 10940 2120 11000 2160
rect 11040 2120 11100 2160
rect 11140 2120 11200 2160
rect 11240 2120 11300 2160
rect 11340 2120 11400 2160
rect 11440 2120 11500 2160
rect 11540 2120 11600 2160
rect 11640 2120 11700 2160
rect 11740 2120 11800 2160
rect 11840 2120 11900 2160
rect 11940 2120 12000 2160
rect 12040 2120 12100 2160
rect 12140 2120 12190 2160
rect 12170 2100 12190 2120
rect 12250 2120 12300 2160
rect 12340 2120 12400 2160
rect 12440 2120 12500 2160
rect 12540 2120 12600 2160
rect 12640 2120 12700 2160
rect 12740 2120 12800 2160
rect 12840 2120 12900 2160
rect 12940 2120 13000 2160
rect 13040 2120 13100 2160
rect 13140 2120 13200 2160
rect 13240 2120 13300 2160
rect 13340 2120 13400 2160
rect 13440 2120 13500 2160
rect 13540 2120 13600 2160
rect 13640 2120 13700 2160
rect 13740 2120 13800 2160
rect 13840 2120 13900 2160
rect 13940 2120 14000 2160
rect 14040 2120 14100 2160
rect 14140 2120 14200 2160
rect 14240 2120 14300 2160
rect 14340 2120 14400 2160
rect 14440 2120 14500 2160
rect 14540 2120 14600 2160
rect 14640 2120 14700 2160
rect 14740 2120 14800 2160
rect 14840 2120 14900 2160
rect 14940 2120 15000 2160
rect 15040 2120 15100 2160
rect 15140 2120 15200 2160
rect 15240 2120 15300 2160
rect 15340 2120 15400 2160
rect 15440 2120 15500 2160
rect 15540 2120 15600 2160
rect 15640 2120 15700 2160
rect 15740 2120 15800 2160
rect 15840 2120 15900 2160
rect 15940 2120 16000 2160
rect 16040 2120 16100 2160
rect 16140 2120 16200 2160
rect 16240 2120 16300 2160
rect 16340 2120 16400 2160
rect 16440 2120 16500 2160
rect 16540 2120 16600 2160
rect 16640 2120 16700 2160
rect 16740 2120 16800 2160
rect 16840 2120 16900 2160
rect 16940 2120 17000 2160
rect 17040 2120 17100 2160
rect 17140 2120 17200 2160
rect 17240 2120 17300 2160
rect 17340 2120 17420 2160
rect 12250 2100 12270 2120
rect 12170 2080 12270 2100
rect 12520 1990 12580 2120
rect 13120 1990 13180 2120
rect 13800 1990 13860 2120
rect 12410 1970 12470 1990
rect 12410 1930 12420 1970
rect 12460 1930 12470 1970
rect 12410 1870 12470 1930
rect 12410 1830 12420 1870
rect 12460 1830 12470 1870
rect 12170 1660 12270 1680
rect 12170 1640 12190 1660
rect 1720 1600 1770 1640
rect 1810 1600 1870 1640
rect 1910 1600 1970 1640
rect 2010 1600 2070 1640
rect 2110 1600 2170 1640
rect 2210 1600 2270 1640
rect 2310 1600 2370 1640
rect 2410 1600 2470 1640
rect 2510 1600 2570 1640
rect 2610 1600 2670 1640
rect 2710 1600 2770 1640
rect 2810 1600 2870 1640
rect 2910 1600 2970 1640
rect 3010 1600 3070 1640
rect 3110 1600 3170 1640
rect 3210 1600 3270 1640
rect 3310 1600 3370 1640
rect 3410 1600 3470 1640
rect 3510 1600 3570 1640
rect 3610 1600 3670 1640
rect 3710 1600 3770 1640
rect 3810 1600 3870 1640
rect 3910 1600 3970 1640
rect 4010 1600 4070 1640
rect 4110 1600 4170 1640
rect 4210 1600 4270 1640
rect 4310 1600 4370 1640
rect 4410 1600 4470 1640
rect 4510 1600 4570 1640
rect 4610 1600 4670 1640
rect 4710 1600 4770 1640
rect 4810 1600 4870 1640
rect 4910 1600 4970 1640
rect 5010 1600 5070 1640
rect 5110 1600 5170 1640
rect 5210 1600 5270 1640
rect 5310 1600 5370 1640
rect 5410 1600 5470 1640
rect 5510 1600 5570 1640
rect 5610 1600 5670 1640
rect 5710 1600 5770 1640
rect 5810 1600 5870 1640
rect 5910 1600 5970 1640
rect 6010 1600 6070 1640
rect 6110 1600 6170 1640
rect 6210 1600 6270 1640
rect 6310 1600 6370 1640
rect 6410 1600 6470 1640
rect 6510 1600 6570 1640
rect 6610 1600 6670 1640
rect 6710 1600 6770 1640
rect 6810 1600 6870 1640
rect 6910 1600 6970 1640
rect 7010 1600 7070 1640
rect 7110 1600 7170 1640
rect 7210 1600 7270 1640
rect 7310 1600 7370 1640
rect 7410 1600 7470 1640
rect 7510 1600 7570 1640
rect 7610 1600 7670 1640
rect 7710 1600 7770 1640
rect 7810 1600 7870 1640
rect 7910 1600 7970 1640
rect 8010 1600 8070 1640
rect 8110 1600 8170 1640
rect 8210 1600 8270 1640
rect 8310 1600 8370 1640
rect 8410 1600 8470 1640
rect 8510 1600 8570 1640
rect 8610 1600 8670 1640
rect 8710 1600 8770 1640
rect 8810 1600 8870 1640
rect 8910 1600 8970 1640
rect 9010 1600 9070 1640
rect 9110 1600 9170 1640
rect 9210 1600 9270 1640
rect 9310 1600 9370 1640
rect 9410 1600 9470 1640
rect 9510 1600 9570 1640
rect 9610 1600 9670 1640
rect 9710 1600 9770 1640
rect 9810 1600 9870 1640
rect 9910 1600 9970 1640
rect 10010 1600 10070 1640
rect 10110 1600 10170 1640
rect 10210 1600 10270 1640
rect 10310 1600 10370 1640
rect 10410 1600 10470 1640
rect 10510 1600 10570 1640
rect 10610 1600 10670 1640
rect 10710 1600 10770 1640
rect 10810 1600 10870 1640
rect 10910 1600 10970 1640
rect 11010 1600 11070 1640
rect 11110 1600 11170 1640
rect 11210 1600 11270 1640
rect 11310 1600 11370 1640
rect 11410 1600 11470 1640
rect 11510 1600 11570 1640
rect 11610 1600 11670 1640
rect 11710 1600 11770 1640
rect 11810 1600 11870 1640
rect 11910 1600 11970 1640
rect 12010 1600 12070 1640
rect 12110 1600 12190 1640
rect 12250 1600 12270 1660
rect 1780 1530 1860 1550
rect 1780 1490 1800 1530
rect 1840 1490 1860 1530
rect 1780 1470 1860 1490
rect 1800 1430 1840 1470
rect 1960 1430 2000 1600
rect 2180 1430 2220 1600
rect 2650 1430 2690 1600
rect 2730 1510 2810 1530
rect 2730 1470 2750 1510
rect 2790 1470 2810 1510
rect 2860 1520 2940 1540
rect 2860 1480 2880 1520
rect 2920 1480 2940 1520
rect 2860 1470 2940 1480
rect 2730 1450 2810 1470
rect 2880 1430 2920 1470
rect 2990 1430 3030 1600
rect 3210 1430 3250 1600
rect 3650 1430 3690 1600
rect 3800 1520 3880 1540
rect 3800 1480 3820 1520
rect 3860 1480 3880 1520
rect 3800 1470 3880 1480
rect 4330 1430 4370 1600
rect 4550 1430 4590 1600
rect 5020 1430 5060 1600
rect 5360 1520 5440 1540
rect 5360 1480 5380 1520
rect 5420 1480 5440 1520
rect 5360 1470 5440 1480
rect 5480 1430 5520 1600
rect 5830 1430 5870 1600
rect 6080 1430 6120 1600
rect 6300 1430 6340 1600
rect 6630 1430 6670 1600
rect 7290 1430 7330 1600
rect 7510 1430 7550 1600
rect 7974 1530 8040 1550
rect 7974 1490 7984 1530
rect 8024 1490 8040 1530
rect 7974 1470 8040 1490
rect 8080 1430 8120 1600
rect 8340 1520 8380 1600
rect 8590 1520 8630 1600
rect 8810 1520 8850 1600
rect 9360 1520 9400 1600
rect 9640 1520 9680 1600
rect 9890 1520 9930 1600
rect 10110 1520 10150 1600
rect 10660 1520 10700 1600
rect 10940 1520 10980 1600
rect 11190 1520 11230 1600
rect 11410 1520 11450 1600
rect 11960 1520 12000 1600
rect 12170 1580 12270 1600
rect 12410 1640 12470 1830
rect 12410 1600 12420 1640
rect 12460 1600 12470 1640
rect 8330 1500 8390 1520
rect 8470 1500 8530 1520
rect 8330 1460 8340 1500
rect 8380 1460 8390 1500
rect 8330 1440 8390 1460
rect 8430 1460 8480 1500
rect 8520 1460 8530 1500
rect 8430 1440 8530 1460
rect 8580 1500 8640 1520
rect 8580 1460 8590 1500
rect 8630 1460 8640 1500
rect 8580 1440 8640 1460
rect 8690 1500 8750 1520
rect 8690 1460 8700 1500
rect 8740 1460 8750 1500
rect 8690 1440 8750 1460
rect 8800 1500 8860 1520
rect 8800 1460 8810 1500
rect 8850 1460 8860 1500
rect 8800 1440 8860 1460
rect 8910 1500 8970 1520
rect 8910 1460 8920 1500
rect 8960 1460 8970 1500
rect 9130 1500 9190 1520
rect 9130 1480 9140 1500
rect 8910 1440 8970 1460
rect 9010 1460 9140 1480
rect 9180 1460 9190 1500
rect 9010 1440 9190 1460
rect 9240 1500 9300 1520
rect 9240 1460 9250 1500
rect 9290 1460 9300 1500
rect 9240 1440 9300 1460
rect 9350 1500 9410 1520
rect 9350 1460 9360 1500
rect 9400 1460 9410 1500
rect 9350 1440 9410 1460
rect 9460 1500 9520 1520
rect 9460 1460 9470 1500
rect 9510 1460 9520 1500
rect 9460 1440 9520 1460
rect 9630 1500 9690 1520
rect 9770 1500 9830 1520
rect 9630 1460 9640 1500
rect 9680 1460 9690 1500
rect 9630 1440 9690 1460
rect 9730 1460 9780 1500
rect 9820 1460 9830 1500
rect 9730 1440 9830 1460
rect 9880 1500 9940 1520
rect 9880 1460 9890 1500
rect 9930 1460 9940 1500
rect 9880 1440 9940 1460
rect 9990 1500 10050 1520
rect 9990 1460 10000 1500
rect 10040 1460 10050 1500
rect 9990 1440 10050 1460
rect 10100 1500 10160 1520
rect 10100 1460 10110 1500
rect 10150 1460 10160 1500
rect 10100 1440 10160 1460
rect 10210 1500 10270 1520
rect 10210 1460 10220 1500
rect 10260 1460 10270 1500
rect 10430 1500 10490 1520
rect 10430 1480 10440 1500
rect 10210 1440 10270 1460
rect 10310 1460 10440 1480
rect 10480 1460 10490 1500
rect 10310 1440 10490 1460
rect 10540 1500 10600 1520
rect 10540 1460 10550 1500
rect 10590 1460 10600 1500
rect 10540 1440 10600 1460
rect 10650 1500 10710 1520
rect 10650 1460 10660 1500
rect 10700 1460 10710 1500
rect 10650 1440 10710 1460
rect 10760 1500 10820 1520
rect 10760 1460 10770 1500
rect 10810 1460 10820 1500
rect 10760 1440 10820 1460
rect 10930 1500 10990 1520
rect 11070 1500 11130 1520
rect 10930 1460 10940 1500
rect 10980 1460 10990 1500
rect 10930 1440 10990 1460
rect 11030 1460 11080 1500
rect 11120 1460 11130 1500
rect 11030 1440 11130 1460
rect 11180 1500 11240 1520
rect 11180 1460 11190 1500
rect 11230 1460 11240 1500
rect 11180 1440 11240 1460
rect 11290 1500 11350 1520
rect 11290 1460 11300 1500
rect 11340 1460 11350 1500
rect 11290 1440 11350 1460
rect 11400 1500 11460 1520
rect 11400 1460 11410 1500
rect 11450 1460 11460 1500
rect 11400 1440 11460 1460
rect 11510 1500 11570 1520
rect 11510 1460 11520 1500
rect 11560 1460 11570 1500
rect 11730 1500 11790 1520
rect 11730 1480 11740 1500
rect 11510 1440 11570 1460
rect 11610 1460 11740 1480
rect 11780 1460 11790 1500
rect 11610 1440 11790 1460
rect 11840 1500 11900 1520
rect 11840 1460 11850 1500
rect 11890 1460 11900 1500
rect 11840 1440 11900 1460
rect 11950 1500 12010 1520
rect 11950 1460 11960 1500
rect 12000 1460 12010 1500
rect 11950 1440 12010 1460
rect 12060 1500 12120 1520
rect 12060 1460 12070 1500
rect 12110 1460 12120 1500
rect 12060 1440 12120 1460
rect 1800 1410 1900 1430
rect 1800 1370 1850 1410
rect 1890 1370 1900 1410
rect 1800 1350 1900 1370
rect 1950 1410 2010 1430
rect 1950 1370 1960 1410
rect 2000 1370 2010 1410
rect 1950 1350 2010 1370
rect 2060 1410 2120 1430
rect 2060 1370 2070 1410
rect 2110 1370 2120 1410
rect 2060 1350 2120 1370
rect 2170 1410 2230 1430
rect 2170 1370 2180 1410
rect 2220 1370 2230 1410
rect 2170 1350 2230 1370
rect 2280 1410 2340 1430
rect 2420 1410 2480 1430
rect 2280 1370 2290 1410
rect 2330 1370 2340 1410
rect 2280 1350 2340 1370
rect 2380 1370 2430 1410
rect 2470 1370 2480 1410
rect 2380 1350 2480 1370
rect 2530 1410 2590 1430
rect 2530 1370 2540 1410
rect 2580 1370 2590 1410
rect 2530 1350 2590 1370
rect 2640 1410 2700 1430
rect 2640 1370 2650 1410
rect 2690 1370 2700 1410
rect 2640 1350 2700 1370
rect 2870 1410 2930 1430
rect 2870 1370 2880 1410
rect 2920 1370 2930 1410
rect 2870 1350 2930 1370
rect 2980 1410 3040 1430
rect 2980 1370 2990 1410
rect 3030 1370 3040 1410
rect 2980 1350 3040 1370
rect 3090 1410 3150 1430
rect 3090 1370 3100 1410
rect 3140 1370 3150 1410
rect 3090 1350 3150 1370
rect 3200 1410 3260 1430
rect 3200 1370 3210 1410
rect 3250 1370 3260 1410
rect 3200 1350 3260 1370
rect 3310 1410 3370 1430
rect 3310 1370 3320 1410
rect 3360 1370 3370 1410
rect 3310 1350 3370 1370
rect 3530 1410 3590 1430
rect 3530 1370 3540 1410
rect 3580 1370 3590 1410
rect 3530 1350 3590 1370
rect 3640 1410 3700 1430
rect 3640 1370 3650 1410
rect 3690 1370 3700 1410
rect 3640 1350 3700 1370
rect 3750 1410 3810 1430
rect 3750 1370 3760 1410
rect 3800 1370 3810 1410
rect 3750 1350 3810 1370
rect 3860 1410 3920 1430
rect 3860 1370 3870 1410
rect 3910 1370 3920 1410
rect 3860 1350 3920 1370
rect 3970 1410 4030 1430
rect 4210 1410 4270 1430
rect 3970 1370 3980 1410
rect 4020 1370 4070 1410
rect 3970 1350 4070 1370
rect 1610 1260 1690 1280
rect 1610 1220 1630 1260
rect 1670 1240 1690 1260
rect 1800 1240 1840 1350
rect 2070 1310 2110 1350
rect 2290 1310 2330 1350
rect 1670 1220 1840 1240
rect 1890 1290 2330 1310
rect 1890 1250 1910 1290
rect 1950 1270 2330 1290
rect 1950 1250 1970 1270
rect 1890 1230 1970 1250
rect 1610 1200 1840 1220
rect 1800 1110 1840 1200
rect 1760 1090 1840 1110
rect 2000 1090 2060 1110
rect 1760 1050 1780 1090
rect 1820 1050 2010 1090
rect 2050 1050 2060 1090
rect 1760 1030 1840 1050
rect 2000 1030 2060 1050
rect 2110 1090 2250 1110
rect 2110 1050 2120 1090
rect 2160 1050 2200 1090
rect 2240 1050 2250 1090
rect 2290 1090 2330 1270
rect 2380 1190 2420 1350
rect 2870 1310 2910 1350
rect 3090 1310 3130 1350
rect 3310 1310 3350 1350
rect 3540 1310 3580 1350
rect 3760 1310 3800 1350
rect 2470 1290 2550 1310
rect 2810 1290 2910 1310
rect 2470 1250 2490 1290
rect 2530 1250 2830 1290
rect 2870 1250 2910 1290
rect 2470 1230 2550 1250
rect 2810 1230 2910 1250
rect 3050 1270 3350 1310
rect 3050 1230 3090 1270
rect 2380 1150 2690 1190
rect 2650 1110 2690 1150
rect 2420 1090 2480 1110
rect 2290 1050 2430 1090
rect 2470 1050 2480 1090
rect 2110 1030 2250 1050
rect 2420 1030 2480 1050
rect 2530 1090 2590 1110
rect 2530 1050 2540 1090
rect 2580 1050 2590 1090
rect 2530 1030 2590 1050
rect 2640 1090 2700 1110
rect 2640 1050 2650 1090
rect 2690 1050 2700 1090
rect 2870 1090 2910 1230
rect 3010 1210 3090 1230
rect 3010 1170 3030 1210
rect 3070 1170 3090 1210
rect 3010 1150 3090 1170
rect 3310 1110 3350 1270
rect 3390 1290 3470 1310
rect 3390 1250 3410 1290
rect 3450 1250 3470 1290
rect 3540 1270 3800 1310
rect 3910 1290 3990 1310
rect 3390 1240 3470 1250
rect 3910 1250 3930 1290
rect 3970 1250 3990 1290
rect 3910 1240 3990 1250
rect 4030 1190 4070 1350
rect 3410 1170 4070 1190
rect 3410 1130 3430 1170
rect 3470 1150 4070 1170
rect 4170 1370 4220 1410
rect 4260 1370 4270 1410
rect 4170 1350 4270 1370
rect 4320 1410 4380 1430
rect 4320 1370 4330 1410
rect 4370 1370 4380 1410
rect 4320 1350 4380 1370
rect 4430 1410 4490 1430
rect 4430 1370 4440 1410
rect 4480 1370 4490 1410
rect 4430 1350 4490 1370
rect 4540 1410 4600 1430
rect 4540 1370 4550 1410
rect 4590 1370 4600 1410
rect 4540 1350 4600 1370
rect 4650 1410 4710 1430
rect 4790 1410 4850 1430
rect 4650 1370 4660 1410
rect 4700 1370 4710 1410
rect 4650 1350 4710 1370
rect 4750 1370 4800 1410
rect 4840 1370 4850 1410
rect 4750 1350 4850 1370
rect 4900 1410 4960 1430
rect 4900 1370 4910 1410
rect 4950 1370 4960 1410
rect 4900 1350 4960 1370
rect 5010 1410 5150 1430
rect 5350 1410 5410 1430
rect 5010 1370 5020 1410
rect 5060 1370 5100 1410
rect 5140 1370 5150 1410
rect 5010 1350 5150 1370
rect 5190 1370 5360 1410
rect 5400 1370 5410 1410
rect 3470 1130 3490 1150
rect 3410 1110 3490 1130
rect 3540 1110 3580 1150
rect 3870 1110 3910 1150
rect 4170 1110 4210 1350
rect 4440 1310 4480 1350
rect 4660 1310 4700 1350
rect 4260 1290 4700 1310
rect 4260 1250 4280 1290
rect 4320 1270 4700 1290
rect 4320 1250 4340 1270
rect 4260 1240 4340 1250
rect 3090 1090 3150 1110
rect 2870 1050 3100 1090
rect 3140 1050 3150 1090
rect 2640 1030 2700 1050
rect 3090 1030 3150 1050
rect 3200 1090 3260 1110
rect 3200 1050 3210 1090
rect 3250 1050 3260 1090
rect 3200 1030 3260 1050
rect 3310 1090 3370 1110
rect 3310 1050 3320 1090
rect 3360 1050 3370 1090
rect 3310 1030 3370 1050
rect 3530 1090 3590 1110
rect 3530 1050 3540 1090
rect 3580 1050 3590 1090
rect 3530 1030 3590 1050
rect 3640 1090 3700 1110
rect 3640 1050 3650 1090
rect 3690 1050 3700 1090
rect 3640 1030 3700 1050
rect 3750 1090 3820 1110
rect 3750 1050 3760 1090
rect 3800 1050 3820 1090
rect 3750 1030 3820 1050
rect 3860 1090 3920 1110
rect 3860 1050 3870 1090
rect 3910 1050 3920 1090
rect 3860 1030 3920 1050
rect 4130 1090 4210 1110
rect 4370 1090 4430 1110
rect 4130 1050 4150 1090
rect 4190 1050 4380 1090
rect 4420 1050 4430 1090
rect 4130 1030 4210 1050
rect 4370 1030 4430 1050
rect 4480 1090 4620 1110
rect 4480 1050 4490 1090
rect 4530 1050 4570 1090
rect 4610 1050 4620 1090
rect 4660 1090 4700 1270
rect 4750 1190 4790 1350
rect 4840 1290 4920 1310
rect 5050 1290 5130 1310
rect 4840 1250 4860 1290
rect 4900 1250 5070 1290
rect 5110 1250 5130 1290
rect 4840 1230 4920 1250
rect 5050 1240 5130 1250
rect 5190 1190 5230 1370
rect 5350 1350 5410 1370
rect 5460 1410 5520 1430
rect 5460 1370 5470 1410
rect 5510 1370 5520 1410
rect 5460 1350 5520 1370
rect 5710 1410 5770 1430
rect 5710 1370 5720 1410
rect 5760 1370 5770 1410
rect 5710 1350 5770 1370
rect 5820 1410 5880 1430
rect 5820 1370 5830 1410
rect 5870 1370 5880 1410
rect 5820 1350 5880 1370
rect 5960 1410 6020 1430
rect 5960 1370 5970 1410
rect 6010 1370 6020 1410
rect 5960 1350 6020 1370
rect 6070 1410 6130 1430
rect 6070 1370 6080 1410
rect 6120 1370 6130 1410
rect 6070 1350 6130 1370
rect 6180 1410 6240 1430
rect 6180 1370 6190 1410
rect 6230 1370 6240 1410
rect 6180 1350 6240 1370
rect 6290 1410 6350 1430
rect 6290 1370 6300 1410
rect 6340 1370 6350 1410
rect 6290 1350 6350 1370
rect 6400 1410 6460 1430
rect 6400 1370 6410 1410
rect 6450 1370 6460 1410
rect 6400 1350 6460 1370
rect 6540 1410 6680 1430
rect 6540 1370 6550 1410
rect 6590 1370 6630 1410
rect 6670 1370 6680 1410
rect 6540 1350 6680 1370
rect 6730 1410 6790 1430
rect 6730 1370 6740 1410
rect 6780 1370 6790 1410
rect 6730 1350 6790 1370
rect 6840 1410 6900 1430
rect 6840 1370 6850 1410
rect 6890 1370 6900 1410
rect 6840 1350 6900 1370
rect 6950 1410 7010 1430
rect 7170 1410 7230 1430
rect 6950 1370 6960 1410
rect 7000 1370 7050 1410
rect 6950 1350 7050 1370
rect 5290 1290 5370 1310
rect 5720 1300 5760 1350
rect 5290 1250 5310 1290
rect 5350 1270 5370 1290
rect 5630 1280 5760 1300
rect 5630 1270 5650 1280
rect 5350 1250 5650 1270
rect 5290 1240 5650 1250
rect 5690 1240 5760 1280
rect 5960 1260 6000 1350
rect 6180 1310 6220 1350
rect 6400 1310 6440 1350
rect 5290 1230 5760 1240
rect 5630 1220 5760 1230
rect 4750 1150 5060 1190
rect 5020 1110 5060 1150
rect 5110 1170 5510 1190
rect 5110 1130 5130 1170
rect 5170 1150 5510 1170
rect 5170 1130 5190 1150
rect 5110 1110 5190 1130
rect 5250 1110 5290 1150
rect 5470 1110 5510 1150
rect 5720 1110 5760 1220
rect 5900 1240 6000 1260
rect 5900 1200 5920 1240
rect 5960 1200 6000 1240
rect 6140 1270 6440 1310
rect 6140 1230 6180 1270
rect 5900 1180 6000 1200
rect 4790 1090 4850 1110
rect 4660 1050 4800 1090
rect 4840 1050 4850 1090
rect 4480 1030 4620 1050
rect 4790 1030 4850 1050
rect 4900 1090 4960 1110
rect 4900 1050 4910 1090
rect 4950 1050 4960 1090
rect 4900 1030 4960 1050
rect 5010 1090 5070 1110
rect 5010 1050 5020 1090
rect 5060 1050 5070 1090
rect 5010 1030 5070 1050
rect 5240 1090 5300 1110
rect 5240 1050 5250 1090
rect 5290 1050 5300 1090
rect 5240 1030 5300 1050
rect 5350 1090 5410 1110
rect 5350 1050 5360 1090
rect 5400 1050 5410 1090
rect 5350 1030 5410 1050
rect 5460 1090 5520 1110
rect 5460 1050 5470 1090
rect 5510 1050 5520 1090
rect 5460 1030 5520 1050
rect 5600 1090 5660 1110
rect 5600 1050 5610 1090
rect 5650 1050 5660 1090
rect 5600 1030 5660 1050
rect 5710 1090 5770 1110
rect 5710 1050 5720 1090
rect 5760 1050 5770 1090
rect 5710 1030 5770 1050
rect 5820 1090 5880 1110
rect 5820 1050 5830 1090
rect 5870 1050 5880 1090
rect 5960 1090 6000 1180
rect 6100 1210 6180 1230
rect 6100 1170 6120 1210
rect 6160 1170 6180 1210
rect 6100 1150 6180 1170
rect 6400 1110 6440 1270
rect 6530 1290 6610 1310
rect 6890 1290 6970 1310
rect 6530 1250 6550 1290
rect 6590 1250 6910 1290
rect 6950 1250 6970 1290
rect 6530 1240 6610 1250
rect 6890 1240 6970 1250
rect 6500 1170 6890 1190
rect 6500 1130 6520 1170
rect 6560 1150 6890 1170
rect 6560 1130 6580 1150
rect 6500 1110 6580 1130
rect 6630 1110 6670 1150
rect 6850 1110 6890 1150
rect 6180 1090 6240 1110
rect 5960 1050 6190 1090
rect 6230 1050 6240 1090
rect 5820 1030 5880 1050
rect 6180 1030 6240 1050
rect 6290 1090 6350 1110
rect 6290 1050 6300 1090
rect 6340 1050 6350 1090
rect 6290 1030 6350 1050
rect 6400 1090 6460 1110
rect 6400 1050 6410 1090
rect 6450 1050 6460 1090
rect 6400 1030 6460 1050
rect 6620 1090 6680 1110
rect 6620 1050 6630 1090
rect 6670 1050 6680 1090
rect 6620 1030 6680 1050
rect 6730 1090 6790 1110
rect 6730 1050 6740 1090
rect 6780 1050 6790 1090
rect 6730 1030 6790 1050
rect 6840 1090 6900 1110
rect 7010 1090 7050 1350
rect 7130 1370 7180 1410
rect 7220 1370 7230 1410
rect 7130 1350 7230 1370
rect 7280 1410 7340 1430
rect 7280 1370 7290 1410
rect 7330 1370 7340 1410
rect 7280 1350 7340 1370
rect 7390 1410 7450 1430
rect 7390 1370 7400 1410
rect 7440 1370 7450 1410
rect 7390 1350 7450 1370
rect 7500 1410 7560 1430
rect 7500 1370 7510 1410
rect 7550 1370 7560 1410
rect 7500 1350 7560 1370
rect 7610 1410 7670 1430
rect 7610 1370 7620 1410
rect 7660 1370 7670 1410
rect 7830 1410 7890 1430
rect 7830 1390 7840 1410
rect 7610 1350 7670 1370
rect 7710 1370 7840 1390
rect 7880 1370 7890 1410
rect 7710 1350 7890 1370
rect 7940 1410 8000 1430
rect 7940 1370 7950 1410
rect 7990 1370 8000 1410
rect 7940 1350 8000 1370
rect 8050 1410 8120 1430
rect 8050 1370 8060 1410
rect 8100 1370 8120 1410
rect 8050 1350 8120 1370
rect 8160 1410 8220 1430
rect 8160 1370 8170 1410
rect 8210 1370 8220 1410
rect 8160 1350 8220 1370
rect 7130 1110 7170 1350
rect 7400 1310 7440 1350
rect 7620 1310 7660 1350
rect 7220 1290 7660 1310
rect 7220 1250 7240 1290
rect 7280 1270 7660 1290
rect 7280 1250 7300 1270
rect 7220 1240 7300 1250
rect 7550 1110 7590 1270
rect 7710 1230 7750 1350
rect 8170 1310 8210 1350
rect 7800 1290 8210 1310
rect 7800 1250 7820 1290
rect 7860 1270 8210 1290
rect 7860 1250 7880 1270
rect 7800 1230 7880 1250
rect 7630 1210 7750 1230
rect 7630 1170 7650 1210
rect 7690 1190 7750 1210
rect 7690 1170 7850 1190
rect 7630 1150 7850 1170
rect 7810 1110 7850 1150
rect 7950 1110 7990 1270
rect 8170 1110 8210 1270
rect 8270 1270 8350 1290
rect 8270 1230 8290 1270
rect 8330 1250 8350 1270
rect 8430 1250 8470 1440
rect 8700 1400 8740 1440
rect 8920 1400 8960 1440
rect 8520 1380 8960 1400
rect 8520 1340 8540 1380
rect 8580 1360 8960 1380
rect 8580 1340 8600 1360
rect 8520 1320 8600 1340
rect 8330 1230 8470 1250
rect 8270 1210 8470 1230
rect 6840 1050 6850 1090
rect 6890 1050 7050 1090
rect 7090 1090 7170 1110
rect 7240 1090 7300 1110
rect 7090 1050 7110 1090
rect 7150 1050 7250 1090
rect 7290 1050 7300 1090
rect 6840 1030 6900 1050
rect 7090 1030 7170 1050
rect 7240 1030 7300 1050
rect 7350 1090 7490 1110
rect 7350 1050 7360 1090
rect 7400 1050 7440 1090
rect 7480 1050 7490 1090
rect 7350 1030 7490 1050
rect 7550 1090 7640 1110
rect 7550 1050 7590 1090
rect 7630 1050 7640 1090
rect 7550 1030 7640 1050
rect 7690 1090 7750 1110
rect 7690 1050 7700 1090
rect 7740 1050 7750 1090
rect 7690 1030 7750 1050
rect 7800 1090 7860 1110
rect 7800 1050 7810 1090
rect 7850 1050 7860 1090
rect 7800 1030 7860 1050
rect 7940 1090 8000 1110
rect 7940 1050 7950 1090
rect 7990 1050 8000 1090
rect 7940 1030 8000 1050
rect 8050 1090 8110 1110
rect 8050 1050 8060 1090
rect 8100 1050 8110 1090
rect 8050 1030 8110 1050
rect 8160 1090 8220 1110
rect 8160 1050 8170 1090
rect 8210 1050 8220 1090
rect 8430 1090 8470 1210
rect 8850 1110 8890 1360
rect 9010 1230 9050 1440
rect 9470 1400 9510 1440
rect 9100 1380 9510 1400
rect 9100 1340 9120 1380
rect 9160 1360 9510 1380
rect 9160 1340 9180 1360
rect 9100 1320 9180 1340
rect 8930 1210 9050 1230
rect 8930 1170 8950 1210
rect 8990 1190 9050 1210
rect 8990 1170 9150 1190
rect 8930 1150 9150 1170
rect 9110 1110 9150 1150
rect 9250 1110 9290 1360
rect 9470 1110 9510 1360
rect 9570 1270 9650 1290
rect 9570 1230 9590 1270
rect 9630 1250 9650 1270
rect 9730 1250 9770 1440
rect 10000 1400 10040 1440
rect 10220 1400 10260 1440
rect 9820 1380 10260 1400
rect 9820 1340 9840 1380
rect 9880 1360 10260 1380
rect 9880 1340 9900 1360
rect 9820 1320 9900 1340
rect 9630 1230 9770 1250
rect 9570 1210 9770 1230
rect 8540 1090 8600 1110
rect 8430 1050 8550 1090
rect 8590 1050 8600 1090
rect 8160 1030 8220 1050
rect 8540 1030 8600 1050
rect 8650 1090 8790 1110
rect 8650 1050 8660 1090
rect 8700 1050 8740 1090
rect 8780 1050 8790 1090
rect 8650 1030 8790 1050
rect 8850 1090 8940 1110
rect 8850 1050 8890 1090
rect 8930 1050 8940 1090
rect 8850 1030 8940 1050
rect 8990 1090 9050 1110
rect 8990 1050 9000 1090
rect 9040 1050 9050 1090
rect 8990 1030 9050 1050
rect 9100 1090 9160 1110
rect 9100 1050 9110 1090
rect 9150 1050 9160 1090
rect 9100 1030 9160 1050
rect 9240 1090 9300 1110
rect 9240 1050 9250 1090
rect 9290 1050 9300 1090
rect 9240 1030 9300 1050
rect 9350 1090 9410 1110
rect 9350 1050 9360 1090
rect 9400 1050 9410 1090
rect 9350 1030 9410 1050
rect 9460 1090 9520 1110
rect 9460 1050 9470 1090
rect 9510 1050 9520 1090
rect 9730 1090 9770 1210
rect 10150 1110 10190 1360
rect 10310 1230 10350 1440
rect 10770 1400 10810 1440
rect 10400 1380 10810 1400
rect 10400 1340 10420 1380
rect 10460 1360 10810 1380
rect 10460 1340 10480 1360
rect 10400 1320 10480 1340
rect 10230 1210 10350 1230
rect 10230 1170 10250 1210
rect 10290 1190 10350 1210
rect 10290 1170 10450 1190
rect 10230 1150 10450 1170
rect 10410 1110 10450 1150
rect 10550 1110 10590 1360
rect 10770 1110 10810 1360
rect 10870 1270 10950 1290
rect 10870 1230 10890 1270
rect 10930 1250 10950 1270
rect 11030 1250 11070 1440
rect 11300 1400 11340 1440
rect 11520 1400 11560 1440
rect 11120 1380 11560 1400
rect 11120 1340 11140 1380
rect 11180 1360 11560 1380
rect 11180 1340 11200 1360
rect 11120 1320 11200 1340
rect 10930 1230 11070 1250
rect 10870 1210 11070 1230
rect 9840 1090 9900 1110
rect 9730 1050 9850 1090
rect 9890 1050 9900 1090
rect 9460 1030 9520 1050
rect 9840 1030 9900 1050
rect 9950 1090 10090 1110
rect 9950 1050 9960 1090
rect 10000 1050 10040 1090
rect 10080 1050 10090 1090
rect 9950 1030 10090 1050
rect 10150 1090 10240 1110
rect 10150 1050 10190 1090
rect 10230 1050 10240 1090
rect 10150 1030 10240 1050
rect 10290 1090 10350 1110
rect 10290 1050 10300 1090
rect 10340 1050 10350 1090
rect 10290 1030 10350 1050
rect 10400 1090 10460 1110
rect 10400 1050 10410 1090
rect 10450 1050 10460 1090
rect 10400 1030 10460 1050
rect 10540 1090 10600 1110
rect 10540 1050 10550 1090
rect 10590 1050 10600 1090
rect 10540 1030 10600 1050
rect 10650 1090 10710 1110
rect 10650 1050 10660 1090
rect 10700 1050 10710 1090
rect 10650 1030 10710 1050
rect 10760 1090 10820 1110
rect 10760 1050 10770 1090
rect 10810 1050 10820 1090
rect 11030 1090 11070 1210
rect 11450 1110 11490 1360
rect 11610 1230 11650 1440
rect 12070 1400 12110 1440
rect 11700 1380 12110 1400
rect 11700 1340 11720 1380
rect 11760 1360 12110 1380
rect 11760 1340 11780 1360
rect 11700 1320 11780 1340
rect 11530 1210 11650 1230
rect 11530 1170 11550 1210
rect 11590 1190 11650 1210
rect 11590 1170 11750 1190
rect 11530 1150 11750 1170
rect 11710 1110 11750 1150
rect 11850 1110 11890 1360
rect 12070 1110 12110 1360
rect 12410 1400 12470 1600
rect 12520 1970 12660 1990
rect 12520 1930 12530 1970
rect 12570 1930 12610 1970
rect 12650 1930 12660 1970
rect 12520 1870 12660 1930
rect 12520 1830 12530 1870
rect 12570 1830 12610 1870
rect 12650 1830 12660 1870
rect 12520 1810 12660 1830
rect 13010 1970 13070 1990
rect 13010 1930 13020 1970
rect 13060 1930 13070 1970
rect 13010 1870 13070 1930
rect 13010 1830 13020 1870
rect 13060 1830 13070 1870
rect 12520 1660 12580 1810
rect 12520 1640 12660 1660
rect 12520 1600 12530 1640
rect 12570 1600 12610 1640
rect 12650 1600 12660 1640
rect 12520 1580 12660 1600
rect 13010 1640 13070 1830
rect 13010 1600 13020 1640
rect 13060 1600 13070 1640
rect 12630 1520 12710 1540
rect 12630 1480 12650 1520
rect 12690 1480 12710 1520
rect 12630 1460 12710 1480
rect 12410 1360 12420 1400
rect 12460 1360 12470 1400
rect 12410 1340 12470 1360
rect 12520 1400 12580 1420
rect 12520 1360 12530 1400
rect 12570 1360 12580 1400
rect 12520 1310 12580 1360
rect 13010 1400 13070 1600
rect 13120 1970 13260 1990
rect 13120 1930 13130 1970
rect 13170 1930 13210 1970
rect 13250 1930 13260 1970
rect 13120 1870 13260 1930
rect 13120 1830 13130 1870
rect 13170 1830 13210 1870
rect 13250 1830 13260 1870
rect 13120 1810 13260 1830
rect 13610 1970 13670 1990
rect 13610 1930 13620 1970
rect 13660 1930 13670 1970
rect 13610 1870 13670 1930
rect 13610 1830 13620 1870
rect 13660 1830 13670 1870
rect 13120 1660 13180 1810
rect 13120 1640 13260 1660
rect 13120 1600 13130 1640
rect 13170 1600 13210 1640
rect 13250 1600 13260 1640
rect 13120 1580 13260 1600
rect 13610 1640 13670 1830
rect 13610 1600 13620 1640
rect 13660 1600 13670 1640
rect 13230 1520 13310 1540
rect 13230 1480 13250 1520
rect 13290 1480 13310 1520
rect 13230 1460 13310 1480
rect 13010 1360 13020 1400
rect 13060 1360 13070 1400
rect 13010 1340 13070 1360
rect 13120 1400 13180 1420
rect 13120 1360 13130 1400
rect 13170 1360 13180 1400
rect 13120 1310 13180 1360
rect 13610 1400 13670 1600
rect 13720 1970 13940 1990
rect 13720 1930 13730 1970
rect 13770 1930 13810 1970
rect 13850 1930 13890 1970
rect 13930 1930 13940 1970
rect 13720 1870 13940 1930
rect 13720 1830 13730 1870
rect 13770 1830 13810 1870
rect 13850 1830 13890 1870
rect 13930 1830 13940 1870
rect 13720 1810 13940 1830
rect 13990 1970 14050 1990
rect 13990 1930 14000 1970
rect 14040 1930 14050 1970
rect 13990 1870 14050 1930
rect 13990 1830 14000 1870
rect 14040 1850 14050 1870
rect 14040 1830 14260 1850
rect 13990 1810 14260 1830
rect 13720 1660 13780 1810
rect 13720 1640 13860 1660
rect 13720 1600 13730 1640
rect 13770 1600 13810 1640
rect 13850 1600 13860 1640
rect 13720 1580 13860 1600
rect 13830 1520 13910 1540
rect 13830 1480 13850 1520
rect 13890 1480 13910 1520
rect 13830 1460 13910 1480
rect 13610 1360 13620 1400
rect 13660 1360 13670 1400
rect 13610 1340 13670 1360
rect 13720 1400 13780 1420
rect 13720 1360 13730 1400
rect 13770 1360 13780 1400
rect 13720 1310 13780 1360
rect 12290 1290 12370 1310
rect 12290 1250 12310 1290
rect 12350 1250 12370 1290
rect 12290 1230 12370 1250
rect 12520 1290 12970 1310
rect 12520 1250 12910 1290
rect 12950 1250 12970 1290
rect 12520 1230 12970 1250
rect 13120 1290 13570 1310
rect 13120 1250 13510 1290
rect 13550 1250 13570 1290
rect 13120 1230 13570 1250
rect 13720 1290 14140 1310
rect 13720 1250 14080 1290
rect 14120 1250 14140 1290
rect 13720 1230 14140 1250
rect 12410 1190 12470 1210
rect 12410 1150 12420 1190
rect 12460 1150 12470 1190
rect 11140 1090 11200 1110
rect 11030 1050 11150 1090
rect 11190 1050 11200 1090
rect 10760 1030 10820 1050
rect 11140 1030 11200 1050
rect 11250 1090 11390 1110
rect 11250 1050 11260 1090
rect 11300 1050 11340 1090
rect 11380 1050 11390 1090
rect 11250 1030 11390 1050
rect 11450 1090 11540 1110
rect 11450 1050 11490 1090
rect 11530 1050 11540 1090
rect 11450 1030 11540 1050
rect 11590 1090 11650 1110
rect 11590 1050 11600 1090
rect 11640 1050 11650 1090
rect 11590 1030 11650 1050
rect 11700 1090 11760 1110
rect 11700 1050 11710 1090
rect 11750 1050 11760 1090
rect 11700 1030 11760 1050
rect 11840 1090 11900 1110
rect 11840 1050 11850 1090
rect 11890 1050 11900 1090
rect 11840 1030 11900 1050
rect 11950 1090 12010 1110
rect 11950 1050 11960 1090
rect 12000 1050 12010 1090
rect 11950 1030 12010 1050
rect 12060 1090 12120 1110
rect 12060 1050 12070 1090
rect 12110 1050 12120 1090
rect 12060 1030 12120 1050
rect 12410 1090 12470 1150
rect 12410 1050 12420 1090
rect 12460 1050 12470 1090
rect 1620 880 1720 900
rect 1620 820 1640 880
rect 1700 860 1720 880
rect 2120 860 2160 1030
rect 2420 970 2500 990
rect 2420 930 2440 970
rect 2480 930 2500 970
rect 2420 910 2500 930
rect 2540 860 2580 1030
rect 2650 990 2690 1030
rect 2620 970 2690 990
rect 2620 930 2630 970
rect 2670 930 2690 970
rect 2730 990 2810 1010
rect 2730 950 2750 990
rect 2790 950 2810 990
rect 2730 930 2810 950
rect 2620 910 2690 930
rect 3210 860 3250 1030
rect 3540 970 3620 990
rect 3540 930 3560 970
rect 3600 930 3620 970
rect 3540 910 3620 930
rect 3680 970 3740 990
rect 3680 930 3690 970
rect 3730 930 3740 970
rect 3680 910 3740 930
rect 3780 860 3820 1030
rect 4490 860 4530 1030
rect 4800 970 4880 990
rect 4800 930 4820 970
rect 4860 930 4880 970
rect 4800 910 4880 930
rect 4920 860 4960 1030
rect 5020 990 5060 1030
rect 5020 970 5100 990
rect 5020 930 5040 970
rect 5080 930 5100 970
rect 5020 910 5100 930
rect 5360 860 5400 1030
rect 5610 860 5650 1030
rect 5830 860 5870 1030
rect 6190 980 6230 1030
rect 6150 960 6230 980
rect 6150 920 6170 960
rect 6210 920 6230 960
rect 6150 910 6230 920
rect 6300 860 6340 1030
rect 6560 960 6640 980
rect 6560 920 6580 960
rect 6620 920 6640 960
rect 6560 910 6640 920
rect 6740 860 6780 1030
rect 7360 860 7400 1030
rect 7700 860 7740 1030
rect 8060 860 8100 1030
rect 8550 990 8590 1030
rect 8510 970 8590 990
rect 8510 930 8530 970
rect 8570 930 8590 970
rect 8510 910 8590 930
rect 8660 860 8700 1030
rect 9000 860 9040 1030
rect 9090 970 9170 990
rect 9090 930 9110 970
rect 9150 930 9170 970
rect 9090 910 9170 930
rect 9360 860 9400 1030
rect 9850 990 9890 1030
rect 9810 970 9890 990
rect 9810 930 9830 970
rect 9870 930 9890 970
rect 9810 910 9890 930
rect 9960 860 10000 1030
rect 10300 860 10340 1030
rect 10390 970 10470 990
rect 10390 930 10410 970
rect 10450 930 10470 970
rect 10390 910 10470 930
rect 10660 860 10700 1030
rect 11150 990 11190 1030
rect 11110 970 11190 990
rect 11110 930 11130 970
rect 11170 930 11190 970
rect 11110 910 11190 930
rect 11260 860 11300 1030
rect 11600 860 11640 1030
rect 11690 970 11770 990
rect 11690 930 11710 970
rect 11750 930 11770 970
rect 11690 910 11770 930
rect 11960 860 12000 1030
rect 12170 860 12270 880
rect 1700 820 1770 860
rect 1810 820 1870 860
rect 1910 820 1970 860
rect 2010 820 2070 860
rect 2110 820 2170 860
rect 2210 820 2270 860
rect 2310 820 2370 860
rect 2410 820 2470 860
rect 2510 820 2570 860
rect 2610 820 2670 860
rect 2710 820 2770 860
rect 2810 820 2870 860
rect 2910 820 2970 860
rect 3010 820 3070 860
rect 3110 820 3170 860
rect 3210 820 3270 860
rect 3310 820 3370 860
rect 3410 820 3470 860
rect 3510 820 3570 860
rect 3610 820 3670 860
rect 3710 820 3770 860
rect 3810 820 3870 860
rect 3910 820 3970 860
rect 4010 820 4070 860
rect 4110 820 4170 860
rect 4210 820 4270 860
rect 4310 820 4370 860
rect 4410 820 4470 860
rect 4510 820 4570 860
rect 4610 820 4670 860
rect 4710 820 4770 860
rect 4810 820 4870 860
rect 4910 820 4970 860
rect 5010 820 5070 860
rect 5110 820 5170 860
rect 5210 820 5270 860
rect 5310 820 5370 860
rect 5410 820 5470 860
rect 5510 820 5570 860
rect 5610 820 5670 860
rect 5710 820 5770 860
rect 5810 820 5870 860
rect 5910 820 5970 860
rect 6010 820 6070 860
rect 6110 820 6170 860
rect 6210 820 6270 860
rect 6310 820 6370 860
rect 6410 820 6470 860
rect 6510 820 6570 860
rect 6610 820 6670 860
rect 6710 820 6770 860
rect 6810 820 6870 860
rect 6910 820 6970 860
rect 7010 820 7070 860
rect 7110 820 7170 860
rect 7210 820 7270 860
rect 7310 820 7370 860
rect 7410 820 7470 860
rect 7510 820 7570 860
rect 7610 820 7670 860
rect 7710 820 7770 860
rect 7810 820 7870 860
rect 7910 820 7970 860
rect 8010 820 8070 860
rect 8110 820 8170 860
rect 8210 820 8270 860
rect 8310 820 8370 860
rect 8410 820 8470 860
rect 8510 820 8570 860
rect 8610 820 8670 860
rect 8710 820 8770 860
rect 8810 820 8870 860
rect 8910 820 8970 860
rect 9010 820 9070 860
rect 9110 820 9170 860
rect 9210 820 9270 860
rect 9310 820 9370 860
rect 9410 820 9470 860
rect 9510 820 9570 860
rect 9610 820 9670 860
rect 9710 820 9770 860
rect 9810 820 9870 860
rect 9910 820 9970 860
rect 10010 820 10070 860
rect 10110 820 10170 860
rect 10210 820 10270 860
rect 10310 820 10370 860
rect 10410 820 10470 860
rect 10510 820 10570 860
rect 10610 820 10670 860
rect 10710 820 10770 860
rect 10810 820 10870 860
rect 10910 820 10970 860
rect 11010 820 11070 860
rect 11110 820 11170 860
rect 11210 820 11270 860
rect 11310 820 11370 860
rect 11410 820 11470 860
rect 11510 820 11570 860
rect 11610 820 11670 860
rect 11710 820 11770 860
rect 11810 820 11870 860
rect 11910 820 11970 860
rect 12010 820 12070 860
rect 12110 820 12190 860
rect 1620 800 1720 820
rect 12170 800 12190 820
rect 12250 800 12270 860
rect 12170 780 12270 800
rect 12410 850 12470 1050
rect 12520 1190 12580 1230
rect 12520 1150 12530 1190
rect 12570 1150 12580 1190
rect 12520 1090 12580 1150
rect 12520 1050 12530 1090
rect 12570 1050 12580 1090
rect 12520 1030 12580 1050
rect 13010 1190 13070 1210
rect 13010 1150 13020 1190
rect 13060 1150 13070 1190
rect 13010 1090 13070 1150
rect 13010 1050 13020 1090
rect 13060 1050 13070 1090
rect 12700 970 12780 990
rect 12700 930 12720 970
rect 12760 930 12780 970
rect 12700 910 12780 930
rect 12410 810 12420 850
rect 12460 810 12470 850
rect 12410 750 12470 810
rect 12410 710 12420 750
rect 12460 710 12470 750
rect 12410 500 12470 710
rect 12520 850 12670 870
rect 12520 810 12530 850
rect 12570 810 12610 850
rect 12650 810 12670 850
rect 12520 750 12670 810
rect 13010 850 13070 1050
rect 13120 1190 13180 1230
rect 13120 1150 13130 1190
rect 13170 1150 13180 1190
rect 13120 1090 13180 1150
rect 13120 1050 13130 1090
rect 13170 1050 13180 1090
rect 13120 1030 13180 1050
rect 13610 1190 13670 1210
rect 13610 1150 13620 1190
rect 13660 1150 13670 1190
rect 13610 1090 13670 1150
rect 13610 1050 13620 1090
rect 13660 1050 13670 1090
rect 13300 970 13380 990
rect 13300 930 13320 970
rect 13360 930 13380 970
rect 13300 910 13380 930
rect 13010 810 13020 850
rect 13060 810 13070 850
rect 13010 750 13070 810
rect 12520 710 12530 750
rect 12570 710 12610 750
rect 12650 710 12850 750
rect 12520 690 12850 710
rect 12410 460 12420 500
rect 12460 460 12470 500
rect 12410 400 12470 460
rect 12410 360 12420 400
rect 12460 360 12470 400
rect 12410 300 12470 360
rect 12410 260 12420 300
rect 12460 260 12470 300
rect 12410 200 12470 260
rect 12410 160 12420 200
rect 12460 160 12470 200
rect 12410 140 12470 160
rect 12790 520 12850 690
rect 13010 710 13020 750
rect 13060 710 13070 750
rect 12790 500 12930 520
rect 12790 460 12800 500
rect 12840 460 12880 500
rect 12920 460 12930 500
rect 12790 400 12930 460
rect 12790 360 12800 400
rect 12840 360 12880 400
rect 12920 360 12930 400
rect 12790 300 12930 360
rect 12790 260 12800 300
rect 12840 260 12880 300
rect 12920 260 12930 300
rect 12790 200 12930 260
rect 12790 160 12800 200
rect 12840 160 12880 200
rect 12920 160 12930 200
rect 12790 140 12930 160
rect 13010 500 13070 710
rect 13120 850 13270 870
rect 13120 810 13130 850
rect 13170 810 13210 850
rect 13250 810 13270 850
rect 13120 750 13270 810
rect 13610 850 13670 1050
rect 13720 1190 13780 1230
rect 13720 1150 13730 1190
rect 13770 1150 13780 1190
rect 13720 1090 13780 1150
rect 13720 1050 13730 1090
rect 13770 1050 13780 1090
rect 13720 1030 13780 1050
rect 13900 970 13980 990
rect 13900 930 13920 970
rect 13960 930 13980 970
rect 13900 910 13980 930
rect 13610 810 13620 850
rect 13660 810 13670 850
rect 13610 750 13670 810
rect 13120 710 13130 750
rect 13170 710 13210 750
rect 13250 710 13450 750
rect 13120 690 13450 710
rect 13010 460 13020 500
rect 13060 460 13070 500
rect 13010 400 13070 460
rect 13010 360 13020 400
rect 13060 360 13070 400
rect 13010 300 13070 360
rect 13010 260 13020 300
rect 13060 260 13070 300
rect 13010 200 13070 260
rect 13010 160 13020 200
rect 13060 160 13070 200
rect 13010 140 13070 160
rect 13390 520 13450 690
rect 13610 710 13620 750
rect 13660 710 13670 750
rect 13390 500 13530 520
rect 13390 460 13400 500
rect 13440 460 13480 500
rect 13520 460 13530 500
rect 13390 400 13530 460
rect 13390 360 13400 400
rect 13440 360 13480 400
rect 13520 360 13530 400
rect 13390 300 13530 360
rect 13390 260 13400 300
rect 13440 260 13480 300
rect 13520 260 13530 300
rect 13390 200 13530 260
rect 13390 160 13400 200
rect 13440 160 13480 200
rect 13520 160 13530 200
rect 13390 140 13530 160
rect 13610 500 13670 710
rect 13720 850 13870 870
rect 13720 810 13730 850
rect 13770 810 13810 850
rect 13850 810 13870 850
rect 13720 750 13870 810
rect 13720 710 13730 750
rect 13770 710 13810 750
rect 13850 710 14130 750
rect 13720 690 14130 710
rect 14070 520 14130 690
rect 14220 640 14260 1810
rect 14300 1810 14380 1830
rect 14300 1770 14320 1810
rect 14360 1770 14380 1810
rect 14300 1750 14380 1770
rect 14220 620 14590 640
rect 14220 580 14230 620
rect 14270 580 14350 620
rect 14390 580 14470 620
rect 14510 580 14590 620
rect 14220 560 14590 580
rect 13610 460 13620 500
rect 13660 460 13670 500
rect 13610 400 13670 460
rect 13610 360 13620 400
rect 13660 360 13670 400
rect 13610 300 13670 360
rect 13610 260 13620 300
rect 13660 260 13670 300
rect 13610 200 13670 260
rect 13610 160 13620 200
rect 13660 160 13670 200
rect 13610 140 13670 160
rect 13990 500 14210 520
rect 13990 460 14000 500
rect 14040 460 14080 500
rect 14120 460 14160 500
rect 14200 460 14210 500
rect 13990 400 14210 460
rect 13990 360 14000 400
rect 14040 360 14080 400
rect 14120 360 14160 400
rect 14200 360 14210 400
rect 13990 300 14210 360
rect 13990 260 14000 300
rect 14040 260 14080 300
rect 14120 260 14160 300
rect 14200 260 14210 300
rect 13990 200 14210 260
rect 13990 160 14000 200
rect 14040 160 14080 200
rect 14120 160 14160 200
rect 14200 160 14210 200
rect 13990 140 14210 160
rect 14530 500 14590 560
rect 14530 460 14540 500
rect 14580 460 14590 500
rect 14530 400 14590 460
rect 14530 360 14540 400
rect 14580 360 14590 400
rect 14530 300 14590 360
rect 14530 260 14540 300
rect 14580 260 14590 300
rect 14530 200 14590 260
rect 14530 160 14540 200
rect 14580 160 14590 200
rect 14530 140 14590 160
rect 12170 80 12270 100
rect 12170 20 12190 80
rect 12250 60 12270 80
rect 12790 60 12850 140
rect 13390 60 13450 140
rect 14070 60 14130 140
rect 12250 20 12300 60
rect 12340 20 12400 60
rect 12440 20 12500 60
rect 12540 20 12600 60
rect 12640 20 12700 60
rect 12740 20 12800 60
rect 12840 20 12900 60
rect 12940 20 13000 60
rect 13040 20 13100 60
rect 13140 20 13200 60
rect 13240 20 13300 60
rect 13340 20 13400 60
rect 13440 20 13500 60
rect 13540 20 13600 60
rect 13640 20 13700 60
rect 13740 20 13800 60
rect 13840 20 13900 60
rect 13940 20 14000 60
rect 14040 20 14100 60
rect 14140 20 14200 60
rect 14240 20 14300 60
rect 14340 20 14400 60
rect 14440 20 14500 60
rect 14540 20 14640 60
rect 12170 0 12270 20
<< viali >>
rect 3250 15040 3290 15080
rect 3250 14960 3290 15000
rect 3250 14880 3290 14920
rect 920 14498 970 14548
rect 490 14348 540 14398
rect 130 14138 180 14188
rect 1650 14402 1656 14424
rect 1656 14402 1684 14424
rect 1650 14390 1684 14402
rect 1750 14390 1784 14424
rect 1850 14390 1884 14424
rect 1950 14402 1982 14424
rect 1982 14402 1984 14424
rect 2050 14402 2072 14424
rect 2072 14402 2084 14424
rect 2150 14402 2162 14424
rect 2162 14402 2184 14424
rect 1950 14390 1984 14402
rect 2050 14390 2084 14402
rect 2150 14390 2184 14402
rect 1650 14312 1656 14324
rect 1656 14312 1684 14324
rect 1650 14290 1684 14312
rect 1750 14290 1784 14324
rect 1850 14290 1884 14324
rect 1950 14312 1982 14324
rect 1982 14312 1984 14324
rect 2050 14312 2072 14324
rect 2072 14312 2084 14324
rect 2150 14312 2162 14324
rect 2162 14312 2184 14324
rect 1950 14290 1984 14312
rect 2050 14290 2084 14312
rect 2150 14290 2184 14312
rect 1650 14222 1656 14224
rect 1656 14222 1684 14224
rect 1650 14190 1684 14222
rect 1750 14190 1784 14224
rect 1850 14190 1884 14224
rect 1950 14222 1982 14224
rect 1982 14222 1984 14224
rect 2050 14222 2072 14224
rect 2072 14222 2084 14224
rect 2150 14222 2162 14224
rect 2162 14222 2184 14224
rect 1950 14190 1984 14222
rect 2050 14190 2084 14222
rect 2150 14190 2184 14222
rect 1650 14090 1684 14124
rect 1750 14090 1784 14124
rect 1850 14090 1884 14124
rect 1950 14090 1984 14124
rect 2050 14090 2084 14124
rect 2150 14090 2184 14124
rect 1650 13990 1684 14024
rect 1750 13990 1784 14024
rect 1850 13990 1884 14024
rect 1950 13990 1984 14024
rect 2050 13990 2084 14024
rect 2150 13990 2184 14024
rect 1650 13896 1684 13924
rect 1650 13890 1656 13896
rect 1656 13890 1684 13896
rect 1750 13890 1784 13924
rect 1850 13890 1884 13924
rect 1950 13896 1984 13924
rect 2050 13896 2084 13924
rect 2150 13896 2184 13924
rect 1950 13890 1982 13896
rect 1982 13890 1984 13896
rect 2050 13890 2072 13896
rect 2072 13890 2084 13896
rect 2150 13890 2162 13896
rect 2162 13890 2184 13896
rect 3010 14402 3016 14424
rect 3016 14402 3044 14424
rect 3010 14390 3044 14402
rect 3110 14390 3144 14424
rect 3210 14390 3244 14424
rect 3310 14402 3342 14424
rect 3342 14402 3344 14424
rect 3410 14402 3432 14424
rect 3432 14402 3444 14424
rect 3510 14402 3522 14424
rect 3522 14402 3544 14424
rect 3310 14390 3344 14402
rect 3410 14390 3444 14402
rect 3510 14390 3544 14402
rect 3010 14312 3016 14324
rect 3016 14312 3044 14324
rect 3010 14290 3044 14312
rect 3110 14290 3144 14324
rect 3210 14290 3244 14324
rect 3310 14312 3342 14324
rect 3342 14312 3344 14324
rect 3410 14312 3432 14324
rect 3432 14312 3444 14324
rect 3510 14312 3522 14324
rect 3522 14312 3544 14324
rect 3310 14290 3344 14312
rect 3410 14290 3444 14312
rect 3510 14290 3544 14312
rect 3010 14222 3016 14224
rect 3016 14222 3044 14224
rect 3010 14190 3044 14222
rect 3110 14190 3144 14224
rect 3210 14190 3244 14224
rect 3310 14222 3342 14224
rect 3342 14222 3344 14224
rect 3410 14222 3432 14224
rect 3432 14222 3444 14224
rect 3510 14222 3522 14224
rect 3522 14222 3544 14224
rect 3310 14190 3344 14222
rect 3410 14190 3444 14222
rect 3510 14190 3544 14222
rect 3010 14090 3044 14124
rect 3110 14090 3144 14124
rect 3210 14090 3244 14124
rect 3310 14090 3344 14124
rect 3410 14090 3444 14124
rect 3510 14090 3544 14124
rect 3010 13990 3044 14024
rect 3110 13990 3144 14024
rect 3210 13990 3244 14024
rect 3310 13990 3344 14024
rect 3410 13990 3444 14024
rect 3510 13990 3544 14024
rect 3010 13896 3044 13924
rect 3010 13890 3016 13896
rect 3016 13890 3044 13896
rect 3110 13890 3144 13924
rect 3210 13890 3244 13924
rect 3310 13896 3344 13924
rect 3410 13896 3444 13924
rect 3510 13896 3544 13924
rect 3310 13890 3342 13896
rect 3342 13890 3344 13896
rect 3410 13890 3432 13896
rect 3432 13890 3444 13896
rect 3510 13890 3522 13896
rect 3522 13890 3544 13896
rect 4370 14402 4376 14424
rect 4376 14402 4404 14424
rect 4370 14390 4404 14402
rect 4470 14390 4504 14424
rect 4570 14390 4604 14424
rect 4670 14402 4702 14424
rect 4702 14402 4704 14424
rect 4770 14402 4792 14424
rect 4792 14402 4804 14424
rect 4870 14402 4882 14424
rect 4882 14402 4904 14424
rect 4670 14390 4704 14402
rect 4770 14390 4804 14402
rect 4870 14390 4904 14402
rect 4370 14312 4376 14324
rect 4376 14312 4404 14324
rect 4370 14290 4404 14312
rect 4470 14290 4504 14324
rect 4570 14290 4604 14324
rect 4670 14312 4702 14324
rect 4702 14312 4704 14324
rect 4770 14312 4792 14324
rect 4792 14312 4804 14324
rect 4870 14312 4882 14324
rect 4882 14312 4904 14324
rect 4670 14290 4704 14312
rect 4770 14290 4804 14312
rect 4870 14290 4904 14312
rect 4370 14222 4376 14224
rect 4376 14222 4404 14224
rect 4370 14190 4404 14222
rect 4470 14190 4504 14224
rect 4570 14190 4604 14224
rect 4670 14222 4702 14224
rect 4702 14222 4704 14224
rect 4770 14222 4792 14224
rect 4792 14222 4804 14224
rect 4870 14222 4882 14224
rect 4882 14222 4904 14224
rect 4670 14190 4704 14222
rect 4770 14190 4804 14222
rect 4870 14190 4904 14222
rect 4370 14090 4404 14124
rect 4470 14090 4504 14124
rect 4570 14090 4604 14124
rect 4670 14090 4704 14124
rect 4770 14090 4804 14124
rect 4870 14090 4904 14124
rect 4370 13990 4404 14024
rect 4470 13990 4504 14024
rect 4570 13990 4604 14024
rect 4670 13990 4704 14024
rect 4770 13990 4804 14024
rect 4870 13990 4904 14024
rect 4370 13896 4404 13924
rect 4370 13890 4376 13896
rect 4376 13890 4404 13896
rect 4470 13890 4504 13924
rect 4570 13890 4604 13924
rect 4670 13896 4704 13924
rect 4770 13896 4804 13924
rect 4870 13896 4904 13924
rect 4670 13890 4702 13896
rect 4702 13890 4704 13896
rect 4770 13890 4792 13896
rect 4792 13890 4804 13896
rect 4870 13890 4882 13896
rect 4882 13890 4904 13896
rect 5450 14498 5500 14548
rect 5810 14348 5860 14398
rect 6470 14348 6520 14398
rect 130 12790 180 12840
rect 250 12740 300 12790
rect 680 12360 730 12410
rect 1650 13042 1656 13064
rect 1656 13042 1684 13064
rect 1650 13030 1684 13042
rect 1750 13030 1784 13064
rect 1850 13030 1884 13064
rect 1950 13042 1982 13064
rect 1982 13042 1984 13064
rect 2050 13042 2072 13064
rect 2072 13042 2084 13064
rect 2150 13042 2162 13064
rect 2162 13042 2184 13064
rect 1950 13030 1984 13042
rect 2050 13030 2084 13042
rect 2150 13030 2184 13042
rect 1650 12952 1656 12964
rect 1656 12952 1684 12964
rect 1650 12930 1684 12952
rect 1750 12930 1784 12964
rect 1850 12930 1884 12964
rect 1950 12952 1982 12964
rect 1982 12952 1984 12964
rect 2050 12952 2072 12964
rect 2072 12952 2084 12964
rect 2150 12952 2162 12964
rect 2162 12952 2184 12964
rect 1950 12930 1984 12952
rect 2050 12930 2084 12952
rect 2150 12930 2184 12952
rect 1650 12862 1656 12864
rect 1656 12862 1684 12864
rect 1650 12830 1684 12862
rect 1750 12830 1784 12864
rect 1850 12830 1884 12864
rect 1950 12862 1982 12864
rect 1982 12862 1984 12864
rect 2050 12862 2072 12864
rect 2072 12862 2084 12864
rect 2150 12862 2162 12864
rect 2162 12862 2184 12864
rect 1950 12830 1984 12862
rect 2050 12830 2084 12862
rect 2150 12830 2184 12862
rect 1650 12730 1684 12764
rect 1750 12730 1784 12764
rect 1850 12730 1884 12764
rect 1950 12730 1984 12764
rect 2050 12730 2084 12764
rect 2150 12730 2184 12764
rect 1650 12630 1684 12664
rect 1750 12630 1784 12664
rect 1850 12630 1884 12664
rect 1950 12630 1984 12664
rect 2050 12630 2084 12664
rect 2150 12630 2184 12664
rect 1650 12536 1684 12564
rect 1650 12530 1656 12536
rect 1656 12530 1684 12536
rect 1750 12530 1784 12564
rect 1850 12530 1884 12564
rect 1950 12536 1984 12564
rect 2050 12536 2084 12564
rect 2150 12536 2184 12564
rect 1950 12530 1982 12536
rect 1982 12530 1984 12536
rect 2050 12530 2072 12536
rect 2072 12530 2084 12536
rect 2150 12530 2162 12536
rect 2162 12530 2184 12536
rect 3010 13042 3016 13064
rect 3016 13042 3044 13064
rect 3010 13030 3044 13042
rect 3110 13030 3144 13064
rect 3210 13030 3244 13064
rect 3310 13042 3342 13064
rect 3342 13042 3344 13064
rect 3410 13042 3432 13064
rect 3432 13042 3444 13064
rect 3510 13042 3522 13064
rect 3522 13042 3544 13064
rect 3310 13030 3344 13042
rect 3410 13030 3444 13042
rect 3510 13030 3544 13042
rect 3010 12952 3016 12964
rect 3016 12952 3044 12964
rect 3010 12930 3044 12952
rect 3110 12930 3144 12964
rect 3210 12930 3244 12964
rect 3310 12952 3342 12964
rect 3342 12952 3344 12964
rect 3410 12952 3432 12964
rect 3432 12952 3444 12964
rect 3510 12952 3522 12964
rect 3522 12952 3544 12964
rect 3310 12930 3344 12952
rect 3410 12930 3444 12952
rect 3510 12930 3544 12952
rect 3010 12862 3016 12864
rect 3016 12862 3044 12864
rect 3010 12830 3044 12862
rect 3110 12830 3144 12864
rect 3210 12830 3244 12864
rect 3310 12862 3342 12864
rect 3342 12862 3344 12864
rect 3410 12862 3432 12864
rect 3432 12862 3444 12864
rect 3510 12862 3522 12864
rect 3522 12862 3544 12864
rect 3310 12830 3344 12862
rect 3410 12830 3444 12862
rect 3510 12830 3544 12862
rect 3010 12730 3044 12764
rect 3110 12730 3144 12764
rect 3210 12730 3244 12764
rect 3310 12730 3344 12764
rect 3410 12730 3444 12764
rect 3510 12730 3544 12764
rect 3010 12630 3044 12664
rect 3110 12630 3144 12664
rect 3210 12630 3244 12664
rect 3310 12630 3344 12664
rect 3410 12630 3444 12664
rect 3510 12630 3544 12664
rect 3010 12536 3044 12564
rect 3010 12530 3016 12536
rect 3016 12530 3044 12536
rect 3110 12530 3144 12564
rect 3210 12530 3244 12564
rect 3310 12536 3344 12564
rect 3410 12536 3444 12564
rect 3510 12536 3544 12564
rect 3310 12530 3342 12536
rect 3342 12530 3344 12536
rect 3410 12530 3432 12536
rect 3432 12530 3444 12536
rect 3510 12530 3522 12536
rect 3522 12530 3544 12536
rect 4370 13042 4376 13064
rect 4376 13042 4404 13064
rect 4370 13030 4404 13042
rect 4470 13030 4504 13064
rect 4570 13030 4604 13064
rect 4670 13042 4702 13064
rect 4702 13042 4704 13064
rect 4770 13042 4792 13064
rect 4792 13042 4804 13064
rect 4870 13042 4882 13064
rect 4882 13042 4904 13064
rect 4670 13030 4704 13042
rect 4770 13030 4804 13042
rect 4870 13030 4904 13042
rect 4370 12952 4376 12964
rect 4376 12952 4404 12964
rect 4370 12930 4404 12952
rect 4470 12930 4504 12964
rect 4570 12930 4604 12964
rect 4670 12952 4702 12964
rect 4702 12952 4704 12964
rect 4770 12952 4792 12964
rect 4792 12952 4804 12964
rect 4870 12952 4882 12964
rect 4882 12952 4904 12964
rect 4670 12930 4704 12952
rect 4770 12930 4804 12952
rect 4870 12930 4904 12952
rect 4370 12862 4376 12864
rect 4376 12862 4404 12864
rect 4370 12830 4404 12862
rect 4470 12830 4504 12864
rect 4570 12830 4604 12864
rect 4670 12862 4702 12864
rect 4702 12862 4704 12864
rect 4770 12862 4792 12864
rect 4792 12862 4804 12864
rect 4870 12862 4882 12864
rect 4882 12862 4904 12864
rect 4670 12830 4704 12862
rect 4770 12830 4804 12862
rect 4870 12830 4904 12862
rect 4370 12730 4404 12764
rect 4470 12730 4504 12764
rect 4570 12730 4604 12764
rect 4670 12730 4704 12764
rect 4770 12730 4804 12764
rect 4870 12730 4904 12764
rect 4370 12630 4404 12664
rect 4470 12630 4504 12664
rect 4570 12630 4604 12664
rect 4670 12630 4704 12664
rect 4770 12630 4804 12664
rect 4870 12630 4904 12664
rect 4370 12536 4404 12564
rect 4370 12530 4376 12536
rect 4376 12530 4404 12536
rect 4470 12530 4504 12564
rect 4570 12530 4604 12564
rect 4670 12536 4704 12564
rect 4770 12536 4804 12564
rect 4870 12536 4904 12564
rect 4670 12530 4702 12536
rect 4702 12530 4704 12536
rect 4770 12530 4792 12536
rect 4792 12530 4804 12536
rect 4870 12530 4882 12536
rect 4882 12530 4904 12536
rect 5810 13210 5860 13260
rect 6470 13002 6520 13052
rect 5690 12360 5740 12410
rect 1650 11682 1656 11704
rect 1656 11682 1684 11704
rect 1650 11670 1684 11682
rect 1750 11670 1784 11704
rect 1850 11670 1884 11704
rect 1950 11682 1982 11704
rect 1982 11682 1984 11704
rect 2050 11682 2072 11704
rect 2072 11682 2084 11704
rect 2150 11682 2162 11704
rect 2162 11682 2184 11704
rect 1950 11670 1984 11682
rect 2050 11670 2084 11682
rect 2150 11670 2184 11682
rect 1650 11592 1656 11604
rect 1656 11592 1684 11604
rect 1650 11570 1684 11592
rect 1750 11570 1784 11604
rect 1850 11570 1884 11604
rect 1950 11592 1982 11604
rect 1982 11592 1984 11604
rect 2050 11592 2072 11604
rect 2072 11592 2084 11604
rect 2150 11592 2162 11604
rect 2162 11592 2184 11604
rect 1950 11570 1984 11592
rect 2050 11570 2084 11592
rect 2150 11570 2184 11592
rect 1650 11502 1656 11504
rect 1656 11502 1684 11504
rect 1650 11470 1684 11502
rect 1750 11470 1784 11504
rect 1850 11470 1884 11504
rect 1950 11502 1982 11504
rect 1982 11502 1984 11504
rect 2050 11502 2072 11504
rect 2072 11502 2084 11504
rect 2150 11502 2162 11504
rect 2162 11502 2184 11504
rect 1950 11470 1984 11502
rect 2050 11470 2084 11502
rect 2150 11470 2184 11502
rect 1650 11370 1684 11404
rect 1750 11370 1784 11404
rect 1850 11370 1884 11404
rect 1950 11370 1984 11404
rect 2050 11370 2084 11404
rect 2150 11370 2184 11404
rect 1650 11270 1684 11304
rect 1750 11270 1784 11304
rect 1850 11270 1884 11304
rect 1950 11270 1984 11304
rect 2050 11270 2084 11304
rect 2150 11270 2184 11304
rect 1650 11176 1684 11204
rect 1650 11170 1656 11176
rect 1656 11170 1684 11176
rect 1750 11170 1784 11204
rect 1850 11170 1884 11204
rect 1950 11176 1984 11204
rect 2050 11176 2084 11204
rect 2150 11176 2184 11204
rect 1950 11170 1982 11176
rect 1982 11170 1984 11176
rect 2050 11170 2072 11176
rect 2072 11170 2084 11176
rect 2150 11170 2162 11176
rect 2162 11170 2184 11176
rect 3010 11682 3016 11704
rect 3016 11682 3044 11704
rect 3010 11670 3044 11682
rect 3110 11670 3144 11704
rect 3210 11670 3244 11704
rect 3310 11682 3342 11704
rect 3342 11682 3344 11704
rect 3410 11682 3432 11704
rect 3432 11682 3444 11704
rect 3510 11682 3522 11704
rect 3522 11682 3544 11704
rect 3310 11670 3344 11682
rect 3410 11670 3444 11682
rect 3510 11670 3544 11682
rect 3010 11592 3016 11604
rect 3016 11592 3044 11604
rect 3010 11570 3044 11592
rect 3110 11570 3144 11604
rect 3210 11570 3244 11604
rect 3310 11592 3342 11604
rect 3342 11592 3344 11604
rect 3410 11592 3432 11604
rect 3432 11592 3444 11604
rect 3510 11592 3522 11604
rect 3522 11592 3544 11604
rect 3310 11570 3344 11592
rect 3410 11570 3444 11592
rect 3510 11570 3544 11592
rect 3010 11502 3016 11504
rect 3016 11502 3044 11504
rect 3010 11470 3044 11502
rect 3110 11470 3144 11504
rect 3210 11470 3244 11504
rect 3310 11502 3342 11504
rect 3342 11502 3344 11504
rect 3410 11502 3432 11504
rect 3432 11502 3444 11504
rect 3510 11502 3522 11504
rect 3522 11502 3544 11504
rect 3310 11470 3344 11502
rect 3410 11470 3444 11502
rect 3510 11470 3544 11502
rect 3010 11370 3044 11404
rect 3110 11370 3144 11404
rect 3210 11370 3244 11404
rect 3310 11370 3344 11404
rect 3410 11370 3444 11404
rect 3510 11370 3544 11404
rect 3010 11270 3044 11304
rect 3110 11270 3144 11304
rect 3210 11270 3244 11304
rect 3310 11270 3344 11304
rect 3410 11270 3444 11304
rect 3510 11270 3544 11304
rect 3010 11176 3044 11204
rect 3010 11170 3016 11176
rect 3016 11170 3044 11176
rect 3110 11170 3144 11204
rect 3210 11170 3244 11204
rect 3310 11176 3344 11204
rect 3410 11176 3444 11204
rect 3510 11176 3544 11204
rect 3310 11170 3342 11176
rect 3342 11170 3344 11176
rect 3410 11170 3432 11176
rect 3432 11170 3444 11176
rect 3510 11170 3522 11176
rect 3522 11170 3544 11176
rect 4370 11682 4376 11704
rect 4376 11682 4404 11704
rect 4370 11670 4404 11682
rect 4470 11670 4504 11704
rect 4570 11670 4604 11704
rect 4670 11682 4702 11704
rect 4702 11682 4704 11704
rect 4770 11682 4792 11704
rect 4792 11682 4804 11704
rect 4870 11682 4882 11704
rect 4882 11682 4904 11704
rect 4670 11670 4704 11682
rect 4770 11670 4804 11682
rect 4870 11670 4904 11682
rect 4370 11592 4376 11604
rect 4376 11592 4404 11604
rect 4370 11570 4404 11592
rect 4470 11570 4504 11604
rect 4570 11570 4604 11604
rect 4670 11592 4702 11604
rect 4702 11592 4704 11604
rect 4770 11592 4792 11604
rect 4792 11592 4804 11604
rect 4870 11592 4882 11604
rect 4882 11592 4904 11604
rect 4670 11570 4704 11592
rect 4770 11570 4804 11592
rect 4870 11570 4904 11592
rect 4370 11502 4376 11504
rect 4376 11502 4404 11504
rect 4370 11470 4404 11502
rect 4470 11470 4504 11504
rect 4570 11470 4604 11504
rect 4670 11502 4702 11504
rect 4702 11502 4704 11504
rect 4770 11502 4792 11504
rect 4792 11502 4804 11504
rect 4870 11502 4882 11504
rect 4882 11502 4904 11504
rect 4670 11470 4704 11502
rect 4770 11470 4804 11502
rect 4870 11470 4904 11502
rect 4370 11370 4404 11404
rect 4470 11370 4504 11404
rect 4570 11370 4604 11404
rect 4670 11370 4704 11404
rect 4770 11370 4804 11404
rect 4870 11370 4904 11404
rect 4370 11270 4404 11304
rect 4470 11270 4504 11304
rect 4570 11270 4604 11304
rect 4670 11270 4704 11304
rect 4770 11270 4804 11304
rect 4870 11270 4904 11304
rect 4370 11176 4404 11204
rect 4370 11170 4376 11176
rect 4376 11170 4404 11176
rect 4470 11170 4504 11204
rect 4570 11170 4604 11204
rect 4670 11176 4704 11204
rect 4770 11176 4804 11204
rect 4870 11176 4904 11204
rect 4670 11170 4702 11176
rect 4702 11170 4704 11176
rect 4770 11170 4792 11176
rect 4792 11170 4804 11176
rect 4870 11170 4882 11176
rect 4882 11170 4904 11176
rect 2552 10560 2602 10610
rect 3950 10560 4000 10610
rect 1090 10170 1130 10210
rect 5480 10210 5520 10250
rect 5480 10130 5520 10170
rect 1170 10000 1210 10040
rect 1330 10000 1370 10040
rect 1490 10000 1530 10040
rect 1650 10000 1690 10040
rect 1810 10000 1850 10040
rect 1970 10000 2010 10040
rect 2130 10000 2170 10040
rect 2290 10000 2330 10040
rect 2450 10000 2490 10040
rect 2610 10000 2650 10040
rect 2770 10000 2810 10040
rect 2930 10000 2970 10040
rect 3090 10000 3130 10040
rect 3250 10000 3290 10040
rect 3410 10000 3450 10040
rect 3570 10000 3610 10040
rect 3730 10000 3770 10040
rect 3890 10000 3930 10040
rect 4050 10000 4090 10040
rect 4210 10000 4250 10040
rect 4370 10000 4410 10040
rect 4530 10000 4570 10040
rect 4690 10000 4730 10040
rect 4850 10000 4890 10040
rect 5010 10000 5050 10040
rect 5170 10000 5210 10040
rect 1910 9730 1950 9770
rect 4590 9730 4630 9770
rect 11770 9750 11830 9810
rect 750 9130 790 9170
rect 930 9090 970 9130
rect 1170 9090 1210 9130
rect 1410 9090 1450 9130
rect 1650 9090 1690 9130
rect 2290 9090 2330 9130
rect 2530 9090 2570 9130
rect 2770 9090 2810 9130
rect 3070 9120 3110 9160
rect 5750 9610 5790 9650
rect 5750 9510 5790 9550
rect 5750 9410 5790 9450
rect 5750 9310 5790 9350
rect 5750 9210 5790 9250
rect 3430 9120 3470 9160
rect 3730 9090 3770 9130
rect 3970 9090 4010 9130
rect 4210 9090 4250 9130
rect 4850 9090 4890 9130
rect 5090 9090 5130 9130
rect 5330 9090 5370 9130
rect 5570 9090 5610 9130
rect 1433 8718 1467 8752
rect 1793 8718 1827 8752
rect 1913 8718 1947 8752
rect 2273 8718 2307 8752
rect 2393 8718 2427 8752
rect 2810 8690 2850 8730
rect 1370 8600 1410 8640
rect 1490 8600 1530 8640
rect 1610 8600 1650 8640
rect 1730 8600 1770 8640
rect 1850 8600 1890 8640
rect 1970 8600 2010 8640
rect 2090 8600 2130 8640
rect 2210 8600 2250 8640
rect 2330 8600 2370 8640
rect 2450 8600 2490 8640
rect 2570 8600 2610 8640
rect 2810 8610 2850 8650
rect 1534 8488 1568 8522
rect 1692 8488 1726 8522
rect 2016 8488 2050 8522
rect 2170 8488 2204 8522
rect 2494 8488 2528 8522
rect 2810 8530 2850 8570
rect 3690 8690 3730 8730
rect 4113 8718 4147 8752
rect 4233 8718 4267 8752
rect 4593 8718 4627 8752
rect 4713 8718 4747 8752
rect 5073 8718 5107 8752
rect 3690 8610 3730 8650
rect 3930 8600 3970 8640
rect 4050 8600 4090 8640
rect 4170 8600 4210 8640
rect 4290 8600 4330 8640
rect 4410 8600 4450 8640
rect 4530 8600 4570 8640
rect 4650 8600 4690 8640
rect 4770 8600 4810 8640
rect 4890 8600 4930 8640
rect 5010 8600 5050 8640
rect 5130 8600 5170 8640
rect 3690 8530 3730 8570
rect 4012 8488 4046 8522
rect 4336 8488 4370 8522
rect 4490 8488 4524 8522
rect 4814 8488 4848 8522
rect 4972 8488 5006 8522
rect 710 7890 750 7930
rect 890 7880 930 7920
rect 1370 7880 1410 7920
rect 1610 7880 1650 7920
rect 2090 7880 2130 7920
rect 2330 7880 2370 7920
rect 2750 7880 2790 7920
rect 3750 7880 3790 7920
rect 4170 7880 4210 7920
rect 4410 7880 4450 7920
rect 4890 7880 4930 7920
rect 5130 7880 5170 7920
rect 5610 7880 5650 7920
rect 5790 7890 5830 7930
rect 530 7760 570 7800
rect 530 7660 570 7700
rect 650 7760 690 7800
rect 650 7660 690 7700
rect 770 7760 810 7800
rect 770 7660 810 7700
rect 890 7760 930 7800
rect 890 7660 930 7700
rect 1010 7760 1050 7800
rect 1010 7660 1050 7700
rect 1130 7760 1170 7800
rect 1130 7660 1170 7700
rect 1250 7760 1290 7800
rect 1250 7660 1290 7700
rect 1370 7760 1410 7800
rect 1370 7660 1410 7700
rect 1490 7760 1530 7800
rect 1490 7660 1530 7700
rect 1610 7760 1650 7800
rect 1610 7660 1650 7700
rect 1730 7760 1770 7800
rect 1730 7660 1770 7700
rect 1850 7760 1890 7800
rect 1850 7660 1890 7700
rect 1970 7760 2010 7800
rect 1970 7660 2010 7700
rect 2090 7760 2130 7800
rect 2090 7660 2130 7700
rect 2210 7760 2250 7800
rect 2210 7660 2250 7700
rect 2330 7760 2370 7800
rect 2330 7660 2370 7700
rect 2450 7760 2490 7800
rect 2450 7660 2490 7700
rect 2570 7760 2610 7800
rect 2570 7660 2610 7700
rect 2690 7760 2730 7800
rect 2690 7660 2730 7700
rect 2810 7760 2850 7800
rect 2810 7660 2850 7700
rect 2930 7760 2970 7800
rect 2930 7660 2970 7700
rect 3570 7760 3610 7800
rect 3570 7660 3610 7700
rect 3690 7760 3730 7800
rect 3690 7660 3730 7700
rect 3810 7760 3850 7800
rect 3810 7660 3850 7700
rect 3930 7760 3970 7800
rect 3930 7660 3970 7700
rect 4050 7760 4090 7800
rect 4050 7660 4090 7700
rect 4170 7760 4210 7800
rect 4170 7660 4210 7700
rect 4290 7760 4330 7800
rect 4290 7660 4330 7700
rect 4410 7760 4450 7800
rect 4410 7660 4450 7700
rect 4530 7760 4570 7800
rect 4530 7660 4570 7700
rect 4650 7760 4690 7800
rect 4650 7660 4690 7700
rect 4770 7760 4810 7800
rect 4770 7660 4810 7700
rect 4890 7760 4930 7800
rect 4890 7660 4930 7700
rect 5010 7760 5050 7800
rect 5010 7660 5050 7700
rect 5130 7760 5170 7800
rect 5130 7660 5170 7700
rect 5250 7760 5290 7800
rect 5250 7660 5290 7700
rect 5370 7760 5410 7800
rect 5370 7660 5410 7700
rect 5490 7760 5530 7800
rect 5490 7660 5530 7700
rect 5610 7760 5650 7800
rect 5610 7660 5650 7700
rect 5730 7760 5770 7800
rect 5730 7660 5770 7700
rect 5850 7760 5890 7800
rect 5850 7660 5890 7700
rect 5970 7760 6010 7800
rect 5970 7660 6010 7700
rect 530 7540 570 7580
rect 2930 7540 2970 7580
rect 3570 7540 3610 7580
rect 5970 7540 6010 7580
rect 1900 6720 1940 6760
rect 2080 6720 2120 6760
rect 2260 6720 2300 6760
rect 2440 6720 2480 6760
rect 2620 6720 2660 6760
rect 2800 6720 2840 6760
rect 2980 6720 3020 6760
rect 3160 6720 3200 6760
rect 3340 6720 3380 6760
rect 3520 6720 3560 6760
rect 3700 6720 3740 6760
rect 3880 6720 3920 6760
rect 4060 6720 4100 6760
rect 4240 6720 4280 6760
rect 4420 6720 4460 6760
rect 4600 6720 4640 6760
rect 1630 6600 1670 6640
rect 1630 6500 1670 6540
rect 1630 6400 1670 6440
rect 1630 6300 1670 6340
rect 1630 6200 1670 6240
rect 1630 6100 1670 6140
rect 1810 6600 1850 6640
rect 1810 6500 1850 6540
rect 1810 6400 1850 6440
rect 1810 6300 1850 6340
rect 1810 6200 1850 6240
rect 1810 6100 1850 6140
rect 1990 6600 2030 6640
rect 1990 6500 2030 6540
rect 1990 6400 2030 6440
rect 1990 6300 2030 6340
rect 1990 6200 2030 6240
rect 1990 6100 2030 6140
rect 2170 6600 2210 6640
rect 2170 6500 2210 6540
rect 2170 6400 2210 6440
rect 2170 6300 2210 6340
rect 2170 6200 2210 6240
rect 2170 6100 2210 6140
rect 2350 6600 2390 6640
rect 2350 6500 2390 6540
rect 2350 6400 2390 6440
rect 2350 6300 2390 6340
rect 2350 6200 2390 6240
rect 2350 6100 2390 6140
rect 2530 6600 2570 6640
rect 2530 6500 2570 6540
rect 2530 6400 2570 6440
rect 2530 6300 2570 6340
rect 2530 6200 2570 6240
rect 2530 6100 2570 6140
rect 2710 6600 2750 6640
rect 2710 6500 2750 6540
rect 2710 6400 2750 6440
rect 2710 6300 2750 6340
rect 2710 6200 2750 6240
rect 2710 6100 2750 6140
rect 2890 6600 2930 6640
rect 2890 6500 2930 6540
rect 2890 6400 2930 6440
rect 2890 6300 2930 6340
rect 2890 6200 2930 6240
rect 2890 6100 2930 6140
rect 3070 6600 3110 6640
rect 3070 6500 3110 6540
rect 3070 6400 3110 6440
rect 3070 6300 3110 6340
rect 3070 6200 3110 6240
rect 3070 6100 3110 6140
rect 3250 6600 3290 6640
rect 3250 6500 3290 6540
rect 3250 6400 3290 6440
rect 3250 6300 3290 6340
rect 3250 6200 3290 6240
rect 3250 6100 3290 6140
rect 3430 6600 3470 6640
rect 3430 6500 3470 6540
rect 3430 6400 3470 6440
rect 3430 6300 3470 6340
rect 3430 6200 3470 6240
rect 3430 6100 3470 6140
rect 3610 6600 3650 6640
rect 3610 6500 3650 6540
rect 3610 6400 3650 6440
rect 3610 6300 3650 6340
rect 3610 6200 3650 6240
rect 3610 6100 3650 6140
rect 3790 6600 3830 6640
rect 3790 6500 3830 6540
rect 3790 6400 3830 6440
rect 3790 6300 3830 6340
rect 3790 6200 3830 6240
rect 3790 6100 3830 6140
rect 3970 6600 4010 6640
rect 3970 6500 4010 6540
rect 3970 6400 4010 6440
rect 3970 6300 4010 6340
rect 3970 6200 4010 6240
rect 3970 6100 4010 6140
rect 4150 6600 4190 6640
rect 4150 6500 4190 6540
rect 4150 6400 4190 6440
rect 4150 6300 4190 6340
rect 4150 6200 4190 6240
rect 4150 6100 4190 6140
rect 4330 6600 4370 6640
rect 4330 6500 4370 6540
rect 4330 6400 4370 6440
rect 4330 6300 4370 6340
rect 4330 6200 4370 6240
rect 4330 6100 4370 6140
rect 4510 6600 4550 6640
rect 4510 6500 4550 6540
rect 4510 6400 4550 6440
rect 4510 6300 4550 6340
rect 4510 6200 4550 6240
rect 4510 6100 4550 6140
rect 4690 6600 4730 6640
rect 4690 6500 4730 6540
rect 4690 6400 4730 6440
rect 4690 6300 4730 6340
rect 4690 6200 4730 6240
rect 4690 6100 4730 6140
rect 4870 6600 4910 6640
rect 4870 6500 4910 6540
rect 5600 6520 5640 6560
rect 5720 6520 5760 6560
rect 5840 6520 5880 6560
rect 4870 6400 4910 6440
rect 4870 6300 4910 6340
rect 5500 6400 5540 6440
rect 5500 6300 5540 6340
rect 5610 6400 5650 6440
rect 5610 6300 5650 6340
rect 5720 6400 5760 6440
rect 5720 6300 5760 6340
rect 5830 6400 5870 6440
rect 5830 6300 5870 6340
rect 5940 6400 5980 6440
rect 5940 6300 5980 6340
rect 4870 6200 4910 6240
rect 5500 6180 5540 6220
rect 5720 6180 5760 6220
rect 5940 6180 5980 6220
rect 8430 8530 8470 8580
rect 8430 8390 8470 8440
rect 8830 8530 8870 8580
rect 8830 8390 8870 8440
rect 9230 8530 9270 8580
rect 9230 8390 9270 8440
rect 9630 8530 9670 8580
rect 9630 8390 9670 8440
rect 10030 8530 10070 8580
rect 10030 8390 10070 8440
rect 8230 8270 8270 8310
rect 9810 8230 9850 8270
rect 10230 8270 10270 8310
rect 7990 8120 8030 8160
rect 8090 8120 8130 8160
rect 8190 8120 8230 8160
rect 8290 8120 8330 8160
rect 8390 8120 8430 8160
rect 8490 8120 8530 8160
rect 8590 8120 8630 8160
rect 8690 8120 8730 8160
rect 8790 8120 8830 8160
rect 8890 8120 8930 8160
rect 8990 8120 9030 8160
rect 9090 8120 9130 8160
rect 9190 8120 9230 8160
rect 9290 8120 9330 8160
rect 9390 8120 9430 8160
rect 9490 8120 9530 8160
rect 9590 8120 9630 8160
rect 9690 8120 9730 8160
rect 9790 8120 9830 8160
rect 9890 8120 9930 8160
rect 9990 8120 10030 8160
rect 10090 8120 10130 8160
rect 10190 8120 10230 8160
rect 10290 8120 10330 8160
rect 10390 8120 10430 8160
rect 10490 8120 10530 8160
rect 10590 8120 10630 8160
rect 10690 8120 10730 8160
rect 10790 8120 10830 8160
rect 10890 8120 10930 8160
rect 9810 8010 9850 8050
rect 8450 7400 8490 7440
rect 9590 7730 9630 7770
rect 9350 7560 9390 7600
rect 8890 7400 8930 7440
rect 10030 7710 10070 7750
rect 11770 7810 11840 7880
rect 10730 7610 10770 7650
rect 11940 7560 11980 7600
rect 8770 7020 8810 7060
rect 11770 7310 11840 7380
rect 7990 6910 8030 6950
rect 8090 6910 8130 6950
rect 8190 6910 8230 6950
rect 8290 6910 8330 6950
rect 8390 6910 8430 6950
rect 8490 6910 8530 6950
rect 8590 6910 8630 6950
rect 8690 6910 8730 6950
rect 8790 6910 8830 6950
rect 8890 6910 8930 6950
rect 8990 6910 9030 6950
rect 9090 6910 9130 6950
rect 9190 6910 9230 6950
rect 9290 6910 9330 6950
rect 9390 6910 9430 6950
rect 9490 6910 9530 6950
rect 9590 6910 9630 6950
rect 9690 6910 9730 6950
rect 9790 6910 9830 6950
rect 9890 6910 9930 6950
rect 9990 6910 10030 6950
rect 10090 6910 10130 6950
rect 10190 6910 10230 6950
rect 10290 6910 10330 6950
rect 10390 6910 10430 6950
rect 10490 6910 10530 6950
rect 10590 6910 10630 6950
rect 10690 6910 10730 6950
rect 10790 6910 10830 6950
rect 10890 6910 10930 6950
rect 8350 6750 8390 6790
rect 8770 6800 8810 6840
rect 8550 6630 8590 6670
rect 8550 6530 8590 6570
rect 8550 6430 8590 6470
rect 8550 6330 8590 6370
rect 8550 6230 8590 6270
rect 8950 6630 8990 6670
rect 8950 6530 8990 6570
rect 8950 6430 8990 6470
rect 8950 6330 8990 6370
rect 8950 6230 8990 6270
rect 9350 6630 9390 6670
rect 9350 6530 9390 6570
rect 9350 6430 9390 6470
rect 9350 6330 9390 6370
rect 9350 6230 9390 6270
rect 9750 6630 9790 6670
rect 9750 6530 9790 6570
rect 9750 6430 9790 6470
rect 9750 6330 9790 6370
rect 9750 6230 9790 6270
rect 10150 6630 10190 6670
rect 10150 6530 10190 6570
rect 10150 6430 10190 6470
rect 10150 6330 10190 6370
rect 10150 6230 10190 6270
rect 4870 6100 4910 6140
rect 1630 5980 1670 6020
rect 1990 5980 2030 6020
rect 2350 5980 2390 6020
rect 2710 5980 2750 6020
rect 3070 5980 3110 6020
rect 3430 5980 3470 6020
rect 3790 5980 3830 6020
rect 4150 5980 4190 6020
rect 4510 5980 4550 6020
rect 4870 5980 4910 6020
rect 1808 5718 1842 5752
rect 1918 5718 1952 5752
rect 2028 5718 2062 5752
rect 2138 5718 2172 5752
rect 2248 5718 2282 5752
rect 2358 5718 2392 5752
rect 2468 5718 2502 5752
rect 2578 5718 2612 5752
rect 2688 5718 2722 5752
rect 2798 5718 2832 5752
rect 3708 5718 3742 5752
rect 3818 5718 3852 5752
rect 3928 5718 3962 5752
rect 4038 5718 4072 5752
rect 4148 5718 4182 5752
rect 4258 5718 4292 5752
rect 4368 5718 4402 5752
rect 4478 5718 4512 5752
rect 4588 5718 4622 5752
rect 4698 5718 4732 5752
rect 1560 5600 1600 5640
rect 1640 5600 1680 5640
rect 1560 5500 1600 5540
rect 1640 5500 1680 5540
rect 1750 5600 1790 5640
rect 1750 5500 1790 5540
rect 1860 5600 1900 5640
rect 1860 5500 1900 5540
rect 1970 5600 2010 5640
rect 1970 5500 2010 5540
rect 2080 5600 2120 5640
rect 2080 5500 2120 5540
rect 2190 5600 2230 5640
rect 2190 5500 2230 5540
rect 2300 5600 2340 5640
rect 2300 5500 2340 5540
rect 2410 5600 2450 5640
rect 2410 5500 2450 5540
rect 2520 5600 2560 5640
rect 2520 5500 2560 5540
rect 2630 5600 2670 5640
rect 2630 5500 2670 5540
rect 2740 5600 2780 5640
rect 2740 5500 2780 5540
rect 2850 5600 2890 5640
rect 2850 5500 2890 5540
rect 2960 5600 3000 5640
rect 3040 5600 3080 5640
rect 2960 5500 3000 5540
rect 3040 5500 3080 5540
rect 3460 5600 3500 5640
rect 3540 5600 3580 5640
rect 3460 5500 3500 5540
rect 3540 5500 3580 5540
rect 3650 5600 3690 5640
rect 3650 5500 3690 5540
rect 3760 5600 3800 5640
rect 3760 5500 3800 5540
rect 3870 5600 3910 5640
rect 3870 5500 3910 5540
rect 3980 5600 4020 5640
rect 3980 5500 4020 5540
rect 4090 5600 4130 5640
rect 4090 5500 4130 5540
rect 4200 5600 4240 5640
rect 4200 5500 4240 5540
rect 4310 5600 4350 5640
rect 4310 5500 4350 5540
rect 4420 5600 4460 5640
rect 4420 5500 4460 5540
rect 4530 5600 4570 5640
rect 4530 5500 4570 5540
rect 4640 5600 4680 5640
rect 4640 5500 4680 5540
rect 4750 5600 4790 5640
rect 4750 5500 4790 5540
rect 4860 5600 4900 5640
rect 4940 5600 4980 5640
rect 4860 5500 4900 5540
rect 4940 5500 4980 5540
rect 1640 5380 1680 5420
rect 2960 5380 3000 5420
rect 3540 5380 3580 5420
rect 4860 5380 4900 5420
rect 11770 5380 11830 5440
rect 11610 5020 11680 5090
rect 1750 4880 1790 4920
rect 1880 4890 1920 4930
rect 1980 4890 2020 4930
rect 2080 4890 2120 4930
rect 2180 4890 2220 4930
rect 2280 4890 2320 4930
rect 2380 4890 2420 4930
rect 2480 4890 2520 4930
rect 2580 4890 2620 4930
rect 2680 4890 2720 4930
rect 2780 4890 2820 4930
rect 2880 4890 2920 4930
rect 2980 4890 3020 4930
rect 3080 4890 3120 4930
rect 3180 4890 3220 4930
rect 3280 4890 3320 4930
rect 3380 4890 3420 4930
rect 3480 4890 3520 4930
rect 3580 4890 3620 4930
rect 3680 4890 3720 4930
rect 3780 4890 3820 4930
rect 3880 4890 3920 4930
rect 3980 4890 4020 4930
rect 4080 4890 4120 4930
rect 4180 4890 4220 4930
rect 4280 4890 4320 4930
rect 4380 4890 4420 4930
rect 4480 4890 4520 4930
rect 4580 4890 4620 4930
rect 4680 4890 4720 4930
rect 4780 4890 4820 4930
rect 4880 4890 4920 4930
rect 4980 4890 5020 4930
rect 5080 4890 5120 4930
rect 5180 4890 5220 4930
rect 5280 4890 5320 4930
rect 5380 4890 5420 4930
rect 5480 4890 5520 4930
rect 5580 4890 5620 4930
rect 5680 4890 5720 4930
rect 5780 4890 5820 4930
rect 5880 4890 5920 4930
rect 5980 4890 6020 4930
rect 6080 4890 6120 4930
rect 6180 4890 6220 4930
rect 6280 4890 6320 4930
rect 6380 4890 6420 4930
rect 6480 4890 6520 4930
rect 6580 4890 6620 4930
rect 6680 4890 6720 4930
rect 6780 4890 6820 4930
rect 6880 4890 6920 4930
rect 2570 4780 2610 4820
rect 1950 4430 1990 4470
rect 4290 4780 4330 4820
rect 6360 4780 6400 4820
rect 3860 4430 3900 4470
rect 5030 4390 5070 4430
rect 5160 4420 5200 4460
rect 7900 4520 7940 4560
rect 8000 4520 8040 4560
rect 8100 4520 8140 4560
rect 8200 4520 8240 4560
rect 8300 4520 8340 4560
rect 8400 4520 8440 4560
rect 8500 4520 8540 4560
rect 8600 4520 8640 4560
rect 8700 4520 8740 4560
rect 8800 4520 8840 4560
rect 8900 4520 8940 4560
rect 9000 4520 9040 4560
rect 9100 4520 9140 4560
rect 9200 4520 9240 4560
rect 9300 4520 9340 4560
rect 9400 4520 9440 4560
rect 9500 4520 9540 4560
rect 9600 4520 9640 4560
rect 9700 4520 9740 4560
rect 9800 4520 9840 4560
rect 9900 4520 9940 4560
rect 10000 4520 10040 4560
rect 10100 4520 10140 4560
rect 10200 4520 10240 4560
rect 10300 4520 10340 4560
rect 10400 4520 10440 4560
rect 10500 4520 10540 4560
rect 10600 4520 10640 4560
rect 10700 4520 10740 4560
rect 10800 4520 10840 4560
rect 10900 4520 10940 4560
rect 11000 4520 11040 4560
rect 6660 4360 6700 4400
rect 6900 4360 6940 4400
rect 1920 3700 1980 3760
rect 4160 3820 4200 3860
rect 8480 3840 8520 3880
rect 2080 3710 2120 3750
rect 2180 3710 2220 3750
rect 2280 3710 2320 3750
rect 2380 3710 2420 3750
rect 2480 3710 2520 3750
rect 2580 3710 2620 3750
rect 2680 3710 2720 3750
rect 2780 3710 2820 3750
rect 2880 3710 2920 3750
rect 2980 3710 3020 3750
rect 3080 3710 3120 3750
rect 3180 3710 3220 3750
rect 3280 3710 3320 3750
rect 3380 3710 3420 3750
rect 3480 3710 3520 3750
rect 3580 3710 3620 3750
rect 3680 3710 3720 3750
rect 3780 3710 3820 3750
rect 3880 3710 3920 3750
rect 3980 3710 4020 3750
rect 4080 3710 4120 3750
rect 4180 3710 4220 3750
rect 4280 3710 4320 3750
rect 4380 3710 4420 3750
rect 4480 3710 4520 3750
rect 4580 3710 4620 3750
rect 4680 3710 4720 3750
rect 4780 3710 4820 3750
rect 4880 3710 4920 3750
rect 4980 3710 5020 3750
rect 5080 3710 5120 3750
rect 5180 3710 5220 3750
rect 5280 3710 5320 3750
rect 5380 3710 5420 3750
rect 5480 3710 5520 3750
rect 5580 3710 5620 3750
rect 5680 3710 5720 3750
rect 5780 3710 5820 3750
rect 5880 3710 5920 3750
rect 5980 3710 6020 3750
rect 6080 3710 6120 3750
rect 6180 3710 6220 3750
rect 6280 3710 6320 3750
rect 6380 3710 6420 3750
rect 6480 3710 6520 3750
rect 6580 3710 6620 3750
rect 6680 3710 6720 3750
rect 6780 3710 6820 3750
rect 6880 3710 6920 3750
rect 6980 3710 7020 3750
rect 7080 3710 7120 3750
rect 7230 3720 7270 3760
rect 8610 3750 8650 3790
rect 2610 3600 2650 3640
rect 5730 3600 5770 3640
rect 10000 3840 10040 3880
rect 11370 3840 11440 3910
rect 6660 3570 6700 3610
rect 8410 3600 8450 3610
rect 8410 3570 8450 3600
rect 2040 2990 2080 3030
rect 3880 3030 3920 3070
rect 4960 3030 5000 3070
rect 5160 3020 5200 3060
rect 6910 3030 6950 3070
rect 11200 3670 11240 3710
rect 10440 3460 10480 3500
rect 11370 3430 11440 3500
rect 7910 2800 7950 2840
rect 8010 2800 8050 2840
rect 8110 2800 8150 2840
rect 8210 2800 8250 2840
rect 8310 2800 8350 2840
rect 8410 2800 8450 2840
rect 8510 2800 8550 2840
rect 8610 2800 8650 2840
rect 8710 2800 8750 2840
rect 8810 2800 8850 2840
rect 8910 2800 8950 2840
rect 9010 2800 9050 2840
rect 9110 2800 9150 2840
rect 9210 2800 9250 2840
rect 9310 2800 9350 2840
rect 9410 2800 9450 2840
rect 9510 2800 9550 2840
rect 9610 2800 9650 2840
rect 9710 2800 9750 2840
rect 9810 2800 9850 2840
rect 9910 2800 9950 2840
rect 10010 2800 10050 2840
rect 10110 2800 10150 2840
rect 10210 2800 10250 2840
rect 10310 2800 10350 2840
rect 10410 2800 10450 2840
rect 10510 2800 10550 2840
rect 10610 2800 10650 2840
rect 10710 2800 10750 2840
rect 10810 2800 10850 2840
rect 10910 2800 10950 2840
rect 11010 2800 11050 2840
rect 1750 2540 1790 2580
rect 5810 2640 5850 2680
rect 6450 2640 6490 2680
rect 11720 2640 11790 2710
rect 17110 2660 17180 2730
rect 17610 2660 17680 2730
rect 1880 2530 1920 2570
rect 1980 2530 2020 2570
rect 2080 2530 2120 2570
rect 2180 2530 2220 2570
rect 2280 2530 2320 2570
rect 2380 2530 2420 2570
rect 2480 2530 2520 2570
rect 2580 2530 2620 2570
rect 2680 2530 2720 2570
rect 2780 2530 2820 2570
rect 2880 2530 2920 2570
rect 2980 2530 3020 2570
rect 3080 2530 3120 2570
rect 3180 2530 3220 2570
rect 3280 2530 3320 2570
rect 3380 2530 3420 2570
rect 3480 2530 3520 2570
rect 3580 2530 3620 2570
rect 3680 2530 3720 2570
rect 3780 2530 3820 2570
rect 3880 2530 3920 2570
rect 3980 2530 4020 2570
rect 4080 2530 4120 2570
rect 4180 2530 4220 2570
rect 4280 2530 4320 2570
rect 4380 2530 4420 2570
rect 4480 2530 4520 2570
rect 4580 2530 4620 2570
rect 4680 2530 4720 2570
rect 4780 2530 4820 2570
rect 4880 2530 4920 2570
rect 4980 2530 5020 2570
rect 5080 2530 5120 2570
rect 5180 2530 5220 2570
rect 5280 2530 5320 2570
rect 5380 2530 5420 2570
rect 5480 2530 5520 2570
rect 5580 2530 5620 2570
rect 5680 2530 5720 2570
rect 5780 2530 5820 2570
rect 5880 2530 5920 2570
rect 5980 2530 6020 2570
rect 6080 2530 6120 2570
rect 6180 2530 6220 2570
rect 6280 2530 6320 2570
rect 6380 2530 6420 2570
rect 6480 2530 6520 2570
rect 6580 2530 6620 2570
rect 6680 2530 6720 2570
rect 6780 2530 6820 2570
rect 6880 2530 6920 2570
rect 14430 2460 14490 2520
rect 23110 2450 23160 2500
rect 25552 2450 25602 2500
rect 7200 2120 7240 2160
rect 7300 2120 7340 2160
rect 7400 2120 7440 2160
rect 7500 2120 7540 2160
rect 7600 2120 7640 2160
rect 7700 2120 7740 2160
rect 7800 2120 7840 2160
rect 7900 2120 7940 2160
rect 8000 2120 8040 2160
rect 8100 2120 8140 2160
rect 8200 2120 8240 2160
rect 8300 2120 8340 2160
rect 8400 2120 8440 2160
rect 8500 2120 8540 2160
rect 8600 2120 8640 2160
rect 8700 2120 8740 2160
rect 8800 2120 8840 2160
rect 8900 2120 8940 2160
rect 9000 2120 9040 2160
rect 9100 2120 9140 2160
rect 9200 2120 9240 2160
rect 9300 2120 9340 2160
rect 9400 2120 9440 2160
rect 9500 2120 9540 2160
rect 9600 2120 9640 2160
rect 9700 2120 9740 2160
rect 9800 2120 9840 2160
rect 9900 2120 9940 2160
rect 10000 2120 10040 2160
rect 10100 2120 10140 2160
rect 10200 2120 10240 2160
rect 10300 2120 10340 2160
rect 10400 2120 10440 2160
rect 10500 2120 10540 2160
rect 10600 2120 10640 2160
rect 10700 2120 10740 2160
rect 10800 2120 10840 2160
rect 10900 2120 10940 2160
rect 11000 2120 11040 2160
rect 11100 2120 11140 2160
rect 11200 2120 11240 2160
rect 11300 2120 11340 2160
rect 11400 2120 11440 2160
rect 11500 2120 11540 2160
rect 11600 2120 11640 2160
rect 11700 2120 11740 2160
rect 11800 2120 11840 2160
rect 11900 2120 11940 2160
rect 12000 2120 12040 2160
rect 12100 2120 12140 2160
rect 12190 2100 12250 2160
rect 12300 2120 12340 2160
rect 12400 2120 12440 2160
rect 12500 2120 12540 2160
rect 12600 2120 12640 2160
rect 12700 2120 12740 2160
rect 12800 2120 12840 2160
rect 12900 2120 12940 2160
rect 13000 2120 13040 2160
rect 13100 2120 13140 2160
rect 13200 2120 13240 2160
rect 13300 2120 13340 2160
rect 13400 2120 13440 2160
rect 13500 2120 13540 2160
rect 13600 2120 13640 2160
rect 13700 2120 13740 2160
rect 13800 2120 13840 2160
rect 13900 2120 13940 2160
rect 14000 2120 14040 2160
rect 14100 2120 14140 2160
rect 14200 2120 14240 2160
rect 14300 2120 14340 2160
rect 14400 2120 14440 2160
rect 14500 2120 14540 2160
rect 14600 2120 14640 2160
rect 14700 2120 14740 2160
rect 14800 2120 14840 2160
rect 14900 2120 14940 2160
rect 15000 2120 15040 2160
rect 15100 2120 15140 2160
rect 15200 2120 15240 2160
rect 15300 2120 15340 2160
rect 15400 2120 15440 2160
rect 15500 2120 15540 2160
rect 15600 2120 15640 2160
rect 15700 2120 15740 2160
rect 15800 2120 15840 2160
rect 15900 2120 15940 2160
rect 16000 2120 16040 2160
rect 16100 2120 16140 2160
rect 16200 2120 16240 2160
rect 16300 2120 16340 2160
rect 16400 2120 16440 2160
rect 16500 2120 16540 2160
rect 16600 2120 16640 2160
rect 16700 2120 16740 2160
rect 16800 2120 16840 2160
rect 16900 2120 16940 2160
rect 17000 2120 17040 2160
rect 17100 2120 17140 2160
rect 17200 2120 17240 2160
rect 17300 2120 17340 2160
rect 1770 1600 1810 1640
rect 1870 1600 1910 1640
rect 1970 1600 2010 1640
rect 2070 1600 2110 1640
rect 2170 1600 2210 1640
rect 2270 1600 2310 1640
rect 2370 1600 2410 1640
rect 2470 1600 2510 1640
rect 2570 1600 2610 1640
rect 2670 1600 2710 1640
rect 2770 1600 2810 1640
rect 2870 1600 2910 1640
rect 2970 1600 3010 1640
rect 3070 1600 3110 1640
rect 3170 1600 3210 1640
rect 3270 1600 3310 1640
rect 3370 1600 3410 1640
rect 3470 1600 3510 1640
rect 3570 1600 3610 1640
rect 3670 1600 3710 1640
rect 3770 1600 3810 1640
rect 3870 1600 3910 1640
rect 3970 1600 4010 1640
rect 4070 1600 4110 1640
rect 4170 1600 4210 1640
rect 4270 1600 4310 1640
rect 4370 1600 4410 1640
rect 4470 1600 4510 1640
rect 4570 1600 4610 1640
rect 4670 1600 4710 1640
rect 4770 1600 4810 1640
rect 4870 1600 4910 1640
rect 4970 1600 5010 1640
rect 5070 1600 5110 1640
rect 5170 1600 5210 1640
rect 5270 1600 5310 1640
rect 5370 1600 5410 1640
rect 5470 1600 5510 1640
rect 5570 1600 5610 1640
rect 5670 1600 5710 1640
rect 5770 1600 5810 1640
rect 5870 1600 5910 1640
rect 5970 1600 6010 1640
rect 6070 1600 6110 1640
rect 6170 1600 6210 1640
rect 6270 1600 6310 1640
rect 6370 1600 6410 1640
rect 6470 1600 6510 1640
rect 6570 1600 6610 1640
rect 6670 1600 6710 1640
rect 6770 1600 6810 1640
rect 6870 1600 6910 1640
rect 6970 1600 7010 1640
rect 7070 1600 7110 1640
rect 7170 1600 7210 1640
rect 7270 1600 7310 1640
rect 7370 1600 7410 1640
rect 7470 1600 7510 1640
rect 7570 1600 7610 1640
rect 7670 1600 7710 1640
rect 7770 1600 7810 1640
rect 7870 1600 7910 1640
rect 7970 1600 8010 1640
rect 8070 1600 8110 1640
rect 8170 1600 8210 1640
rect 8270 1600 8310 1640
rect 8370 1600 8410 1640
rect 8470 1600 8510 1640
rect 8570 1600 8610 1640
rect 8670 1600 8710 1640
rect 8770 1600 8810 1640
rect 8870 1600 8910 1640
rect 8970 1600 9010 1640
rect 9070 1600 9110 1640
rect 9170 1600 9210 1640
rect 9270 1600 9310 1640
rect 9370 1600 9410 1640
rect 9470 1600 9510 1640
rect 9570 1600 9610 1640
rect 9670 1600 9710 1640
rect 9770 1600 9810 1640
rect 9870 1600 9910 1640
rect 9970 1600 10010 1640
rect 10070 1600 10110 1640
rect 10170 1600 10210 1640
rect 10270 1600 10310 1640
rect 10370 1600 10410 1640
rect 10470 1600 10510 1640
rect 10570 1600 10610 1640
rect 10670 1600 10710 1640
rect 10770 1600 10810 1640
rect 10870 1600 10910 1640
rect 10970 1600 11010 1640
rect 11070 1600 11110 1640
rect 11170 1600 11210 1640
rect 11270 1600 11310 1640
rect 11370 1600 11410 1640
rect 11470 1600 11510 1640
rect 11570 1600 11610 1640
rect 11670 1600 11710 1640
rect 11770 1600 11810 1640
rect 11870 1600 11910 1640
rect 11970 1600 12010 1640
rect 12070 1600 12110 1640
rect 12190 1600 12250 1660
rect 1800 1490 1840 1530
rect 2750 1470 2790 1510
rect 2880 1480 2920 1520
rect 3820 1480 3860 1520
rect 5380 1480 5420 1520
rect 7984 1490 8024 1530
rect 1630 1220 1670 1260
rect 3410 1250 3450 1290
rect 3930 1250 3970 1290
rect 4150 1050 4190 1090
rect 5650 1240 5690 1280
rect 12530 1600 12570 1640
rect 12610 1600 12650 1640
rect 12650 1480 12690 1520
rect 13130 1600 13170 1640
rect 13210 1600 13250 1640
rect 13250 1480 13290 1520
rect 13730 1600 13770 1640
rect 13810 1600 13850 1640
rect 13850 1480 13890 1520
rect 12310 1250 12350 1290
rect 14080 1250 14120 1290
rect 1640 820 1700 880
rect 2440 930 2480 970
rect 2630 930 2670 970
rect 2750 950 2790 990
rect 3560 930 3600 970
rect 3690 930 3730 970
rect 4820 930 4860 970
rect 5040 930 5080 970
rect 6170 920 6210 960
rect 6580 920 6620 960
rect 8530 930 8570 970
rect 9110 930 9150 970
rect 9830 930 9870 970
rect 10410 930 10450 970
rect 11130 930 11170 970
rect 11710 930 11750 970
rect 1770 820 1810 860
rect 1870 820 1910 860
rect 1970 820 2010 860
rect 2070 820 2110 860
rect 2170 820 2210 860
rect 2270 820 2310 860
rect 2370 820 2410 860
rect 2470 820 2510 860
rect 2570 820 2610 860
rect 2670 820 2710 860
rect 2770 820 2810 860
rect 2870 820 2910 860
rect 2970 820 3010 860
rect 3070 820 3110 860
rect 3170 820 3210 860
rect 3270 820 3310 860
rect 3370 820 3410 860
rect 3470 820 3510 860
rect 3570 820 3610 860
rect 3670 820 3710 860
rect 3770 820 3810 860
rect 3870 820 3910 860
rect 3970 820 4010 860
rect 4070 820 4110 860
rect 4170 820 4210 860
rect 4270 820 4310 860
rect 4370 820 4410 860
rect 4470 820 4510 860
rect 4570 820 4610 860
rect 4670 820 4710 860
rect 4770 820 4810 860
rect 4870 820 4910 860
rect 4970 820 5010 860
rect 5070 820 5110 860
rect 5170 820 5210 860
rect 5270 820 5310 860
rect 5370 820 5410 860
rect 5470 820 5510 860
rect 5570 820 5610 860
rect 5670 820 5710 860
rect 5770 820 5810 860
rect 5870 820 5910 860
rect 5970 820 6010 860
rect 6070 820 6110 860
rect 6170 820 6210 860
rect 6270 820 6310 860
rect 6370 820 6410 860
rect 6470 820 6510 860
rect 6570 820 6610 860
rect 6670 820 6710 860
rect 6770 820 6810 860
rect 6870 820 6910 860
rect 6970 820 7010 860
rect 7070 820 7110 860
rect 7170 820 7210 860
rect 7270 820 7310 860
rect 7370 820 7410 860
rect 7470 820 7510 860
rect 7570 820 7610 860
rect 7670 820 7710 860
rect 7770 820 7810 860
rect 7870 820 7910 860
rect 7970 820 8010 860
rect 8070 820 8110 860
rect 8170 820 8210 860
rect 8270 820 8310 860
rect 8370 820 8410 860
rect 8470 820 8510 860
rect 8570 820 8610 860
rect 8670 820 8710 860
rect 8770 820 8810 860
rect 8870 820 8910 860
rect 8970 820 9010 860
rect 9070 820 9110 860
rect 9170 820 9210 860
rect 9270 820 9310 860
rect 9370 820 9410 860
rect 9470 820 9510 860
rect 9570 820 9610 860
rect 9670 820 9710 860
rect 9770 820 9810 860
rect 9870 820 9910 860
rect 9970 820 10010 860
rect 10070 820 10110 860
rect 10170 820 10210 860
rect 10270 820 10310 860
rect 10370 820 10410 860
rect 10470 820 10510 860
rect 10570 820 10610 860
rect 10670 820 10710 860
rect 10770 820 10810 860
rect 10870 820 10910 860
rect 10970 820 11010 860
rect 11070 820 11110 860
rect 11170 820 11210 860
rect 11270 820 11310 860
rect 11370 820 11410 860
rect 11470 820 11510 860
rect 11570 820 11610 860
rect 11670 820 11710 860
rect 11770 820 11810 860
rect 11870 820 11910 860
rect 11970 820 12010 860
rect 12070 820 12110 860
rect 12190 800 12250 860
rect 12720 930 12760 970
rect 12610 810 12650 850
rect 13320 930 13360 970
rect 12610 710 12650 750
rect 13210 810 13250 850
rect 13920 930 13960 970
rect 13210 710 13250 750
rect 13810 810 13850 850
rect 13810 710 13850 750
rect 14320 1770 14360 1810
rect 12190 20 12250 80
rect 12300 20 12340 60
rect 12400 20 12440 60
rect 12500 20 12540 60
rect 12600 20 12640 60
rect 12700 20 12740 60
rect 12800 20 12840 60
rect 12900 20 12940 60
rect 13000 20 13040 60
rect 13100 20 13140 60
rect 13200 20 13240 60
rect 13300 20 13340 60
rect 13400 20 13440 60
rect 13500 20 13540 60
rect 13600 20 13640 60
rect 13700 20 13740 60
rect 13800 20 13840 60
rect 13900 20 13940 60
rect 14000 20 14040 60
rect 14100 20 14140 60
rect 14200 20 14240 60
rect 14300 20 14340 60
rect 14400 20 14440 60
rect 14500 20 14540 60
<< metal1 >>
rect 110 15200 190 15210
rect 110 15140 120 15200
rect 180 15140 190 15200
rect 110 14198 190 15140
rect 480 15090 560 15100
rect 480 15030 490 15090
rect 550 15030 560 15090
rect 480 15010 560 15030
rect 480 14950 490 15010
rect 550 14950 560 15010
rect 480 14930 560 14950
rect 480 14870 490 14930
rect 550 14870 560 14930
rect 480 14408 560 14870
rect 910 15090 990 15100
rect 910 15030 920 15090
rect 980 15030 990 15090
rect 910 15010 990 15030
rect 910 14950 920 15010
rect 980 14950 990 15010
rect 910 14930 990 14950
rect 910 14870 920 14930
rect 980 14870 990 14930
rect 910 14560 990 14870
rect 910 14558 980 14560
rect 910 14478 980 14488
rect 480 14328 550 14338
rect 120 14118 190 14128
rect 120 12850 190 12870
rect 0 10220 80 10230
rect 0 10160 10 10220
rect 70 10160 80 10220
rect 0 7100 80 10160
rect 0 7040 10 7100
rect 70 7040 80 7100
rect 0 7030 80 7040
rect 110 7590 190 12780
rect 240 12800 310 12810
rect 240 12726 310 12730
rect 110 7530 120 7590
rect 180 7530 190 7590
rect 110 5770 190 7530
rect 230 8530 310 12726
rect 670 12420 740 12430
rect 670 12340 740 12350
rect 660 10730 740 12340
rect 660 10670 670 10730
rect 730 10670 740 10730
rect 660 10660 740 10670
rect 230 8470 240 8530
rect 300 8470 310 8530
rect 230 7210 310 8470
rect 230 7150 240 7210
rect 300 7150 310 7210
rect 230 7140 310 7150
rect 340 10500 420 10510
rect 340 10440 350 10500
rect 410 10440 420 10500
rect 340 8760 420 10440
rect 340 8700 350 8760
rect 410 8700 420 8760
rect 110 5710 120 5770
rect 180 5710 190 5770
rect 110 5700 190 5710
rect 340 5320 420 8700
rect 610 10390 690 10400
rect 610 10330 620 10390
rect 680 10330 690 10390
rect 610 8060 690 10330
rect 1020 10390 1100 15210
rect 7280 15200 7360 15210
rect 7280 15140 7290 15200
rect 7350 15140 7360 15200
rect 3230 15090 3310 15100
rect 3230 15030 3240 15090
rect 3300 15030 3310 15090
rect 3230 15010 3310 15030
rect 3230 14950 3240 15010
rect 3300 14950 3310 15010
rect 3230 14930 3310 14950
rect 3230 14870 3240 14930
rect 3300 14870 3310 14930
rect 3230 14860 3310 14870
rect 5430 15090 5510 15100
rect 5430 15030 5440 15090
rect 5500 15030 5510 15090
rect 5430 15010 5510 15030
rect 5430 14950 5440 15010
rect 5500 14950 5510 15010
rect 5430 14930 5510 14950
rect 5430 14870 5440 14930
rect 5500 14870 5510 14930
rect 5430 14860 5510 14870
rect 5790 15090 5870 15100
rect 5790 15030 5800 15090
rect 5860 15030 5870 15090
rect 5790 15010 5870 15030
rect 5790 14950 5800 15010
rect 5860 14950 5870 15010
rect 5790 14930 5870 14950
rect 5790 14870 5800 14930
rect 5860 14870 5870 14930
rect 5790 14860 5870 14870
rect 5440 14558 5510 14860
rect 1560 14424 4980 14500
rect 5440 14478 5510 14488
rect 1560 14390 1650 14424
rect 1684 14390 1750 14424
rect 1784 14390 1850 14424
rect 1884 14390 1950 14424
rect 1984 14390 2050 14424
rect 2084 14390 2150 14424
rect 2184 14390 3010 14424
rect 3044 14390 3110 14424
rect 3144 14390 3210 14424
rect 3244 14390 3310 14424
rect 3344 14390 3410 14424
rect 3444 14390 3510 14424
rect 3544 14390 4370 14424
rect 4404 14390 4470 14424
rect 4504 14390 4570 14424
rect 4604 14390 4670 14424
rect 4704 14390 4770 14424
rect 4804 14390 4870 14424
rect 4904 14390 4980 14424
rect 1560 14324 4980 14390
rect 5800 14408 5870 14860
rect 5800 14328 5870 14338
rect 5930 15090 6090 15100
rect 5930 15030 5940 15090
rect 6000 15030 6020 15090
rect 6080 15030 6090 15090
rect 5930 15010 6090 15030
rect 5930 14950 5940 15010
rect 6000 14950 6020 15010
rect 6080 14950 6090 15010
rect 5930 14930 6090 14950
rect 5930 14870 5940 14930
rect 6000 14870 6020 14930
rect 6080 14870 6090 14930
rect 1560 14290 1650 14324
rect 1684 14290 1750 14324
rect 1784 14290 1850 14324
rect 1884 14290 1950 14324
rect 1984 14290 2050 14324
rect 2084 14290 2150 14324
rect 2184 14290 3010 14324
rect 3044 14290 3110 14324
rect 3144 14290 3210 14324
rect 3244 14290 3310 14324
rect 3344 14290 3410 14324
rect 3444 14290 3510 14324
rect 3544 14290 4370 14324
rect 4404 14290 4470 14324
rect 4504 14290 4570 14324
rect 4604 14290 4670 14324
rect 4704 14290 4770 14324
rect 4804 14290 4870 14324
rect 4904 14290 4980 14324
rect 1560 14224 4980 14290
rect 1560 14190 1650 14224
rect 1684 14190 1750 14224
rect 1784 14190 1850 14224
rect 1884 14190 1950 14224
rect 1984 14190 2050 14224
rect 2084 14190 2150 14224
rect 2184 14190 3010 14224
rect 3044 14190 3110 14224
rect 3144 14190 3210 14224
rect 3244 14190 3310 14224
rect 3344 14190 3410 14224
rect 3444 14190 3510 14224
rect 3544 14190 4370 14224
rect 4404 14190 4470 14224
rect 4504 14190 4570 14224
rect 4604 14190 4670 14224
rect 4704 14190 4770 14224
rect 4804 14190 4870 14224
rect 4904 14190 4980 14224
rect 1560 14124 4980 14190
rect 1560 14090 1650 14124
rect 1684 14090 1750 14124
rect 1784 14090 1850 14124
rect 1884 14090 1950 14124
rect 1984 14090 2050 14124
rect 2084 14090 2150 14124
rect 2184 14090 3010 14124
rect 3044 14090 3110 14124
rect 3144 14090 3210 14124
rect 3244 14090 3310 14124
rect 3344 14090 3410 14124
rect 3444 14090 3510 14124
rect 3544 14090 4370 14124
rect 4404 14090 4470 14124
rect 4504 14090 4570 14124
rect 4604 14090 4670 14124
rect 4704 14090 4770 14124
rect 4804 14090 4870 14124
rect 4904 14090 4980 14124
rect 1560 14024 4980 14090
rect 1560 13990 1650 14024
rect 1684 13990 1750 14024
rect 1784 13990 1850 14024
rect 1884 13990 1950 14024
rect 1984 13990 2050 14024
rect 2084 13990 2150 14024
rect 2184 13990 3010 14024
rect 3044 13990 3110 14024
rect 3144 13990 3210 14024
rect 3244 13990 3310 14024
rect 3344 13990 3410 14024
rect 3444 13990 3510 14024
rect 3544 13990 4370 14024
rect 4404 13990 4470 14024
rect 4504 13990 4570 14024
rect 4604 13990 4670 14024
rect 4704 13990 4770 14024
rect 4804 13990 4870 14024
rect 4904 13990 4980 14024
rect 1560 13924 4980 13990
rect 1560 13890 1650 13924
rect 1684 13890 1750 13924
rect 1784 13890 1850 13924
rect 1884 13890 1950 13924
rect 1984 13890 2050 13924
rect 2084 13890 2150 13924
rect 2184 13890 3010 13924
rect 3044 13890 3110 13924
rect 3144 13890 3210 13924
rect 3244 13890 3310 13924
rect 3344 13890 3410 13924
rect 3444 13890 3510 13924
rect 3544 13890 4370 13924
rect 4404 13890 4470 13924
rect 4504 13890 4570 13924
rect 4604 13890 4670 13924
rect 4704 13890 4770 13924
rect 4804 13890 4870 13924
rect 4904 13890 4980 13924
rect 1560 13800 4980 13890
rect 1560 13064 2260 13800
rect 1560 13030 1650 13064
rect 1684 13030 1750 13064
rect 1784 13030 1850 13064
rect 1884 13030 1950 13064
rect 1984 13030 2050 13064
rect 2084 13030 2150 13064
rect 2184 13030 2260 13064
rect 1560 12964 2260 13030
rect 1560 12930 1650 12964
rect 1684 12930 1750 12964
rect 1784 12930 1850 12964
rect 1884 12930 1950 12964
rect 1984 12930 2050 12964
rect 2084 12930 2150 12964
rect 2184 12930 2260 12964
rect 1560 12864 2260 12930
rect 1560 12830 1650 12864
rect 1684 12830 1750 12864
rect 1784 12830 1850 12864
rect 1884 12830 1950 12864
rect 1984 12830 2050 12864
rect 2084 12830 2150 12864
rect 2184 12830 2260 12864
rect 1130 12820 1210 12830
rect 1130 12760 1140 12820
rect 1200 12760 1210 12820
rect 1130 10620 1210 12760
rect 1560 12820 2260 12830
rect 1560 12760 1570 12820
rect 1630 12764 2260 12820
rect 1630 12760 1650 12764
rect 1560 12730 1650 12760
rect 1684 12730 1750 12764
rect 1784 12730 1850 12764
rect 1884 12730 1950 12764
rect 1984 12730 2050 12764
rect 2084 12730 2150 12764
rect 2184 12730 2260 12764
rect 1560 12664 2260 12730
rect 1560 12630 1650 12664
rect 1684 12630 1750 12664
rect 1784 12630 1850 12664
rect 1884 12630 1950 12664
rect 1984 12630 2050 12664
rect 2084 12630 2150 12664
rect 2184 12630 2260 12664
rect 1560 12564 2260 12630
rect 1560 12530 1650 12564
rect 1684 12530 1750 12564
rect 1784 12530 1850 12564
rect 1884 12530 1950 12564
rect 1984 12530 2050 12564
rect 2084 12530 2150 12564
rect 2184 12530 2260 12564
rect 1560 11780 2260 12530
rect 2920 13064 3620 13140
rect 2920 13030 3010 13064
rect 3044 13030 3110 13064
rect 3144 13030 3210 13064
rect 3244 13030 3310 13064
rect 3344 13030 3410 13064
rect 3444 13030 3510 13064
rect 3544 13030 3620 13064
rect 2920 12964 3620 13030
rect 2920 12930 3010 12964
rect 3044 12930 3110 12964
rect 3144 12930 3210 12964
rect 3244 12930 3310 12964
rect 3344 12930 3410 12964
rect 3444 12930 3510 12964
rect 3544 12930 3620 12964
rect 2920 12864 3620 12930
rect 2920 12830 3010 12864
rect 3044 12830 3110 12864
rect 3144 12830 3210 12864
rect 3244 12830 3310 12864
rect 3344 12830 3410 12864
rect 3444 12830 3510 12864
rect 3544 12830 3620 12864
rect 2920 12820 3620 12830
rect 2920 12764 3240 12820
rect 3300 12764 3620 12820
rect 2920 12730 3010 12764
rect 3044 12730 3110 12764
rect 3144 12730 3210 12764
rect 3300 12760 3310 12764
rect 3244 12730 3310 12760
rect 3344 12730 3410 12764
rect 3444 12730 3510 12764
rect 3544 12730 3620 12764
rect 2920 12664 3620 12730
rect 2920 12630 3010 12664
rect 3044 12630 3110 12664
rect 3144 12630 3210 12664
rect 3244 12630 3310 12664
rect 3344 12630 3410 12664
rect 3444 12630 3510 12664
rect 3544 12630 3620 12664
rect 2920 12564 3620 12630
rect 2920 12530 3010 12564
rect 3044 12530 3110 12564
rect 3144 12530 3210 12564
rect 3244 12530 3310 12564
rect 3344 12530 3410 12564
rect 3444 12530 3510 12564
rect 3544 12530 3620 12564
rect 2920 12440 3620 12530
rect 4280 13064 4980 13800
rect 4280 13030 4370 13064
rect 4404 13030 4470 13064
rect 4504 13030 4570 13064
rect 4604 13030 4670 13064
rect 4704 13030 4770 13064
rect 4804 13030 4870 13064
rect 4904 13030 4980 13064
rect 4280 12964 4980 13030
rect 4280 12930 4370 12964
rect 4404 12930 4470 12964
rect 4504 12930 4570 12964
rect 4604 12930 4670 12964
rect 4704 12930 4770 12964
rect 4804 12930 4870 12964
rect 4904 12930 4980 12964
rect 4280 12864 4980 12930
rect 4280 12830 4370 12864
rect 4404 12830 4470 12864
rect 4504 12830 4570 12864
rect 4604 12830 4670 12864
rect 4704 12830 4770 12864
rect 4804 12830 4870 12864
rect 4904 12830 4980 12864
rect 5800 13270 5870 13280
rect 5800 13190 5870 13200
rect 4280 12764 4980 12830
rect 4280 12730 4370 12764
rect 4404 12730 4470 12764
rect 4504 12730 4570 12764
rect 4604 12730 4670 12764
rect 4704 12730 4770 12764
rect 4804 12730 4870 12764
rect 4904 12730 4980 12764
rect 5330 12820 5410 12830
rect 5330 12760 5340 12820
rect 5400 12760 5410 12820
rect 5330 12750 5410 12760
rect 4280 12664 4980 12730
rect 4280 12630 4370 12664
rect 4404 12630 4470 12664
rect 4504 12630 4570 12664
rect 4604 12630 4670 12664
rect 4704 12630 4770 12664
rect 4804 12630 4870 12664
rect 4904 12630 4980 12664
rect 4280 12564 4980 12630
rect 4280 12530 4370 12564
rect 4404 12530 4470 12564
rect 4504 12530 4570 12564
rect 4604 12530 4670 12564
rect 4704 12530 4770 12564
rect 4804 12530 4870 12564
rect 4904 12530 4980 12564
rect 4280 11780 4980 12530
rect 1560 11704 4980 11780
rect 1560 11670 1650 11704
rect 1684 11670 1750 11704
rect 1784 11670 1850 11704
rect 1884 11670 1950 11704
rect 1984 11670 2050 11704
rect 2084 11670 2150 11704
rect 2184 11670 3010 11704
rect 3044 11670 3110 11704
rect 3144 11670 3210 11704
rect 3244 11670 3310 11704
rect 3344 11670 3410 11704
rect 3444 11670 3510 11704
rect 3544 11670 4370 11704
rect 4404 11670 4470 11704
rect 4504 11670 4570 11704
rect 4604 11670 4670 11704
rect 4704 11670 4770 11704
rect 4804 11670 4870 11704
rect 4904 11670 4980 11704
rect 1560 11604 4980 11670
rect 1560 11570 1650 11604
rect 1684 11570 1750 11604
rect 1784 11570 1850 11604
rect 1884 11570 1950 11604
rect 1984 11570 2050 11604
rect 2084 11570 2150 11604
rect 2184 11570 3010 11604
rect 3044 11570 3110 11604
rect 3144 11570 3210 11604
rect 3244 11570 3310 11604
rect 3344 11570 3410 11604
rect 3444 11570 3510 11604
rect 3544 11570 4370 11604
rect 4404 11570 4470 11604
rect 4504 11570 4570 11604
rect 4604 11570 4670 11604
rect 4704 11570 4770 11604
rect 4804 11570 4870 11604
rect 4904 11570 4980 11604
rect 1560 11504 4980 11570
rect 1560 11470 1650 11504
rect 1684 11470 1750 11504
rect 1784 11470 1850 11504
rect 1884 11470 1950 11504
rect 1984 11470 2050 11504
rect 2084 11470 2150 11504
rect 2184 11470 3010 11504
rect 3044 11470 3110 11504
rect 3144 11470 3210 11504
rect 3244 11470 3310 11504
rect 3344 11470 3410 11504
rect 3444 11470 3510 11504
rect 3544 11470 4370 11504
rect 4404 11470 4470 11504
rect 4504 11470 4570 11504
rect 4604 11470 4670 11504
rect 4704 11470 4770 11504
rect 4804 11470 4870 11504
rect 4904 11470 4980 11504
rect 1560 11404 4980 11470
rect 1560 11370 1650 11404
rect 1684 11370 1750 11404
rect 1784 11370 1850 11404
rect 1884 11370 1950 11404
rect 1984 11370 2050 11404
rect 2084 11370 2150 11404
rect 2184 11370 3010 11404
rect 3044 11370 3110 11404
rect 3144 11370 3210 11404
rect 3244 11370 3310 11404
rect 3344 11370 3410 11404
rect 3444 11370 3510 11404
rect 3544 11370 4370 11404
rect 4404 11370 4470 11404
rect 4504 11370 4570 11404
rect 4604 11370 4670 11404
rect 4704 11370 4770 11404
rect 4804 11370 4870 11404
rect 4904 11370 4980 11404
rect 1560 11304 4980 11370
rect 1560 11270 1650 11304
rect 1684 11270 1750 11304
rect 1784 11270 1850 11304
rect 1884 11270 1950 11304
rect 1984 11270 2050 11304
rect 2084 11270 2150 11304
rect 2184 11270 3010 11304
rect 3044 11270 3110 11304
rect 3144 11270 3210 11304
rect 3244 11270 3310 11304
rect 3344 11270 3410 11304
rect 3444 11270 3510 11304
rect 3544 11270 4370 11304
rect 4404 11270 4470 11304
rect 4504 11270 4570 11304
rect 4604 11270 4670 11304
rect 4704 11270 4770 11304
rect 4804 11270 4870 11304
rect 4904 11270 4980 11304
rect 1560 11204 4980 11270
rect 1560 11170 1650 11204
rect 1684 11170 1750 11204
rect 1784 11170 1850 11204
rect 1884 11170 1950 11204
rect 1984 11170 2050 11204
rect 2084 11170 2150 11204
rect 2184 11170 3010 11204
rect 3044 11170 3110 11204
rect 3144 11170 3210 11204
rect 3244 11170 3310 11204
rect 3344 11170 3410 11204
rect 3444 11170 3510 11204
rect 3544 11170 4370 11204
rect 4404 11170 4470 11204
rect 4504 11170 4570 11204
rect 4604 11170 4670 11204
rect 4704 11170 4770 11204
rect 4804 11170 4870 11204
rect 4904 11170 4980 11204
rect 1560 11080 4980 11170
rect 5350 10820 5390 12750
rect 5680 12420 5750 12430
rect 5680 12340 5750 12350
rect 5700 10820 5740 12340
rect 5330 10810 5410 10820
rect 5330 10750 5340 10810
rect 5400 10750 5410 10810
rect 5330 10740 5410 10750
rect 5680 10810 5760 10820
rect 5680 10750 5690 10810
rect 5750 10750 5760 10810
rect 5680 10740 5760 10750
rect 3940 10730 4020 10740
rect 3940 10670 3950 10730
rect 4010 10670 4020 10730
rect 3940 10620 4020 10670
rect 1130 10560 1140 10620
rect 1200 10560 1210 10620
rect 1130 10550 1210 10560
rect 2532 10550 2542 10620
rect 2612 10550 2622 10620
rect 3930 10550 3940 10620
rect 4010 10550 4020 10620
rect 5800 10500 5880 13190
rect 5800 10440 5810 10500
rect 5870 10440 5880 10500
rect 5800 10430 5880 10440
rect 1020 10330 1030 10390
rect 1090 10330 1100 10390
rect 1020 10320 1100 10330
rect 5460 10260 5540 10270
rect 1070 10220 1150 10230
rect 1070 10160 1080 10220
rect 1140 10160 1150 10220
rect 1070 10150 1150 10160
rect 5460 10200 5470 10260
rect 5530 10200 5540 10260
rect 5460 10180 5540 10200
rect 5460 10120 5470 10180
rect 5530 10120 5540 10180
rect 5460 10110 5540 10120
rect 5930 10260 6090 14870
rect 7280 14860 7360 15140
rect 7280 14800 7290 14860
rect 7350 14800 7360 14860
rect 7280 14790 7360 14800
rect 6460 14408 6530 14420
rect 6460 14328 6530 14338
rect 6830 14410 6920 14420
rect 6830 14340 6840 14410
rect 6910 14340 6920 14410
rect 6830 14330 6920 14340
rect 6460 13062 6530 13072
rect 6460 12980 6530 12992
rect 6460 12760 6540 12980
rect 6460 12700 6470 12760
rect 6530 12700 6540 12760
rect 6230 10810 6310 10820
rect 6230 10750 6240 10810
rect 6300 10750 6310 10810
rect 6230 10740 6310 10750
rect 6140 10610 6220 10620
rect 6140 10550 6150 10610
rect 6210 10550 6220 10610
rect 6140 10540 6220 10550
rect 5930 10200 5940 10260
rect 6000 10200 6020 10260
rect 6080 10200 6090 10260
rect 5930 10180 6090 10200
rect 5930 10120 5940 10180
rect 6000 10120 6020 10180
rect 6080 10120 6090 10180
rect 5930 10110 6090 10120
rect 1150 10050 1230 10060
rect 1150 9990 1160 10050
rect 1220 9990 1230 10050
rect 1150 9980 1230 9990
rect 1310 10050 1390 10060
rect 1310 9990 1320 10050
rect 1380 9990 1390 10050
rect 1310 9980 1390 9990
rect 1470 10050 1550 10060
rect 1470 9990 1480 10050
rect 1540 9990 1550 10050
rect 1470 9980 1550 9990
rect 1630 10050 1710 10060
rect 1630 9990 1640 10050
rect 1700 9990 1710 10050
rect 1630 9980 1710 9990
rect 1790 10050 1870 10060
rect 1790 9990 1800 10050
rect 1860 9990 1870 10050
rect 1790 9980 1870 9990
rect 1950 10050 2030 10060
rect 1950 9990 1960 10050
rect 2020 9990 2030 10050
rect 1950 9980 2030 9990
rect 2110 10050 2190 10060
rect 2110 9990 2120 10050
rect 2180 9990 2190 10050
rect 2110 9980 2190 9990
rect 2270 10050 2350 10060
rect 2270 9990 2280 10050
rect 2340 9990 2350 10050
rect 2270 9980 2350 9990
rect 2430 10050 2510 10060
rect 2430 9990 2440 10050
rect 2500 9990 2510 10050
rect 2430 9980 2510 9990
rect 2590 10050 2670 10060
rect 2590 9990 2600 10050
rect 2660 9990 2670 10050
rect 2590 9980 2670 9990
rect 2750 10050 2830 10060
rect 2750 9990 2760 10050
rect 2820 9990 2830 10050
rect 2750 9980 2830 9990
rect 2910 10050 2990 10060
rect 2910 9990 2920 10050
rect 2980 9990 2990 10050
rect 2910 9980 2990 9990
rect 3070 10050 3150 10060
rect 3070 9990 3080 10050
rect 3140 9990 3150 10050
rect 3070 9980 3150 9990
rect 3230 10050 3310 10060
rect 3230 9990 3240 10050
rect 3300 9990 3310 10050
rect 3230 9980 3310 9990
rect 3390 10050 3470 10060
rect 3390 9990 3400 10050
rect 3460 9990 3470 10050
rect 3390 9980 3470 9990
rect 3550 10050 3630 10060
rect 3550 9990 3560 10050
rect 3620 9990 3630 10050
rect 3550 9980 3630 9990
rect 3710 10050 3790 10060
rect 3710 9990 3720 10050
rect 3780 9990 3790 10050
rect 3710 9980 3790 9990
rect 3870 10050 3950 10060
rect 3870 9990 3880 10050
rect 3940 9990 3950 10050
rect 3870 9980 3950 9990
rect 4030 10050 4110 10060
rect 4030 9990 4040 10050
rect 4100 9990 4110 10050
rect 4030 9980 4110 9990
rect 4190 10050 4270 10060
rect 4190 9990 4200 10050
rect 4260 9990 4270 10050
rect 4190 9980 4270 9990
rect 4350 10050 4430 10060
rect 4350 9990 4360 10050
rect 4420 9990 4430 10050
rect 4350 9980 4430 9990
rect 4510 10050 4590 10060
rect 4510 9990 4520 10050
rect 4580 9990 4590 10050
rect 4510 9980 4590 9990
rect 4670 10050 4750 10060
rect 4670 9990 4680 10050
rect 4740 9990 4750 10050
rect 4670 9980 4750 9990
rect 4830 10050 4910 10060
rect 4830 9990 4840 10050
rect 4900 9990 4910 10050
rect 4830 9980 4910 9990
rect 4990 10050 5070 10060
rect 4990 9990 5000 10050
rect 5060 9990 5070 10050
rect 4990 9980 5070 9990
rect 5150 10050 5230 10060
rect 5150 9990 5160 10050
rect 5220 9990 5230 10050
rect 5150 9980 5230 9990
rect 1890 9940 1970 9950
rect 1890 9880 1900 9940
rect 1960 9880 1970 9940
rect 1890 9860 1970 9880
rect 1890 9800 1900 9860
rect 1960 9800 1970 9860
rect 1890 9780 1970 9800
rect 1890 9720 1900 9780
rect 1960 9720 1970 9780
rect 1890 9710 1970 9720
rect 3150 9940 3390 9950
rect 3150 9880 3160 9940
rect 3220 9880 3240 9940
rect 3300 9880 3320 9940
rect 3380 9880 3390 9940
rect 3150 9860 3390 9880
rect 3150 9800 3160 9860
rect 3220 9800 3240 9860
rect 3300 9800 3320 9860
rect 3380 9800 3390 9860
rect 3150 9780 3390 9800
rect 3150 9720 3160 9780
rect 3220 9720 3240 9780
rect 3300 9720 3320 9780
rect 3380 9720 3390 9780
rect 730 9170 810 9190
rect 730 9130 750 9170
rect 790 9130 810 9170
rect 3060 9160 3120 9180
rect 730 9110 810 9130
rect 910 9140 990 9150
rect 750 8880 790 9110
rect 910 9080 920 9140
rect 980 9080 990 9140
rect 910 9060 990 9080
rect 910 9000 920 9060
rect 980 9000 990 9060
rect 910 8980 990 9000
rect 910 8920 920 8980
rect 980 8920 990 8980
rect 910 8910 990 8920
rect 1150 9140 1230 9150
rect 1150 9080 1160 9140
rect 1220 9080 1230 9140
rect 1150 9060 1230 9080
rect 1150 9000 1160 9060
rect 1220 9000 1230 9060
rect 1150 8980 1230 9000
rect 1150 8920 1160 8980
rect 1220 8920 1230 8980
rect 1150 8910 1230 8920
rect 1390 9140 1470 9150
rect 1390 9080 1400 9140
rect 1460 9080 1470 9140
rect 1390 9060 1470 9080
rect 1390 9000 1400 9060
rect 1460 9000 1470 9060
rect 1390 8980 1470 9000
rect 1390 8920 1400 8980
rect 1460 8920 1470 8980
rect 1390 8910 1470 8920
rect 1630 9140 1710 9150
rect 1630 9080 1640 9140
rect 1700 9080 1710 9140
rect 1630 9060 1710 9080
rect 1630 9000 1640 9060
rect 1700 9000 1710 9060
rect 1630 8980 1710 9000
rect 1630 8920 1640 8980
rect 1700 8920 1710 8980
rect 1630 8910 1710 8920
rect 2270 9140 2350 9150
rect 2270 9080 2280 9140
rect 2340 9080 2350 9140
rect 2270 9060 2350 9080
rect 2270 9000 2280 9060
rect 2340 9000 2350 9060
rect 2270 8980 2350 9000
rect 2270 8920 2280 8980
rect 2340 8920 2350 8980
rect 2270 8910 2350 8920
rect 2510 9140 2590 9150
rect 2510 9080 2520 9140
rect 2580 9080 2590 9140
rect 2510 9060 2590 9080
rect 2510 9000 2520 9060
rect 2580 9000 2590 9060
rect 2510 8980 2590 9000
rect 2510 8920 2520 8980
rect 2580 8920 2590 8980
rect 2510 8910 2590 8920
rect 2750 9140 2830 9150
rect 2750 9080 2760 9140
rect 2820 9080 2830 9140
rect 2750 9060 2830 9080
rect 2750 9000 2760 9060
rect 2820 9000 2830 9060
rect 2750 8980 2830 9000
rect 2750 8920 2760 8980
rect 2820 8920 2830 8980
rect 2750 8910 2830 8920
rect 3060 9120 3070 9160
rect 3110 9120 3120 9160
rect 730 8870 810 8880
rect 730 8810 740 8870
rect 800 8810 810 8870
rect 730 8800 810 8810
rect 1480 8870 1560 8880
rect 1480 8810 1490 8870
rect 1550 8810 1560 8870
rect 1480 8800 1560 8810
rect 1700 8870 1780 8880
rect 1700 8810 1710 8870
rect 1770 8810 1780 8870
rect 1700 8800 1780 8810
rect 1960 8870 2040 8880
rect 1960 8810 1970 8870
rect 2030 8810 2040 8870
rect 1960 8800 2040 8810
rect 2180 8870 2260 8880
rect 2180 8810 2190 8870
rect 2250 8810 2260 8870
rect 2180 8800 2260 8810
rect 2440 8870 2520 8880
rect 2440 8810 2450 8870
rect 2510 8810 2520 8870
rect 2440 8800 2520 8810
rect 1421 8760 1479 8770
rect 1421 8708 1423 8760
rect 1475 8708 1479 8760
rect 1421 8700 1479 8708
rect 1510 8660 1540 8800
rect 1720 8660 1750 8800
rect 1781 8760 1839 8770
rect 1781 8708 1783 8760
rect 1835 8708 1839 8760
rect 1781 8700 1839 8708
rect 1901 8760 1959 8770
rect 1901 8708 1903 8760
rect 1955 8708 1959 8760
rect 1901 8700 1959 8708
rect 1990 8660 2020 8800
rect 2200 8660 2230 8800
rect 2261 8760 2319 8770
rect 2261 8708 2263 8760
rect 2315 8708 2319 8760
rect 2261 8700 2319 8708
rect 2381 8760 2439 8770
rect 2381 8708 2383 8760
rect 2435 8708 2439 8760
rect 2381 8700 2439 8708
rect 2470 8660 2500 8800
rect 2790 8740 2870 8750
rect 2790 8680 2800 8740
rect 2860 8680 2870 8740
rect 2790 8660 2870 8680
rect 1360 8640 1420 8660
rect 1360 8600 1370 8640
rect 1410 8600 1420 8640
rect 1360 8330 1420 8600
rect 1480 8640 1540 8660
rect 1480 8600 1490 8640
rect 1530 8600 1540 8640
rect 1480 8580 1540 8600
rect 1600 8640 1660 8660
rect 1600 8600 1610 8640
rect 1650 8600 1660 8640
rect 1600 8580 1660 8600
rect 1720 8640 1780 8660
rect 1720 8600 1730 8640
rect 1770 8600 1780 8640
rect 1720 8580 1780 8600
rect 1840 8640 1900 8660
rect 1840 8600 1850 8640
rect 1890 8600 1900 8640
rect 1840 8580 1900 8600
rect 1960 8640 2020 8660
rect 1960 8600 1970 8640
rect 2010 8600 2020 8640
rect 1960 8580 2020 8600
rect 2080 8640 2140 8660
rect 2080 8600 2090 8640
rect 2130 8600 2140 8640
rect 2080 8580 2140 8600
rect 2200 8640 2260 8660
rect 2200 8600 2210 8640
rect 2250 8600 2260 8640
rect 2200 8580 2260 8600
rect 2320 8640 2380 8660
rect 2320 8600 2330 8640
rect 2370 8600 2380 8640
rect 2320 8580 2380 8600
rect 2440 8640 2500 8660
rect 2440 8600 2450 8640
rect 2490 8600 2500 8640
rect 2440 8580 2500 8600
rect 2560 8640 2620 8660
rect 2560 8600 2570 8640
rect 2610 8600 2620 8640
rect 2560 8580 2620 8600
rect 2790 8600 2800 8660
rect 2860 8600 2870 8660
rect 2790 8580 2870 8600
rect 1522 8532 1580 8540
rect 1522 8480 1526 8532
rect 1578 8480 1580 8532
rect 1522 8470 1580 8480
rect 1610 8440 1650 8580
rect 1680 8532 1738 8540
rect 1680 8480 1684 8532
rect 1736 8480 1738 8532
rect 1680 8470 1738 8480
rect 1590 8430 1670 8440
rect 1590 8370 1600 8430
rect 1660 8370 1670 8430
rect 1350 8320 1430 8330
rect 1350 8260 1360 8320
rect 1420 8260 1430 8320
rect 610 8050 770 8060
rect 610 7990 620 8050
rect 680 7990 700 8050
rect 760 7990 770 8050
rect 610 7980 770 7990
rect 1110 8050 1190 8060
rect 1110 7990 1120 8050
rect 1180 7990 1190 8050
rect 1110 7980 1190 7990
rect 1350 8050 1430 8260
rect 1350 7990 1360 8050
rect 1420 7990 1430 8050
rect 1350 7980 1430 7990
rect 700 7930 760 7980
rect 700 7890 710 7930
rect 750 7890 760 7930
rect 700 7870 760 7890
rect 870 7930 950 7940
rect 870 7870 880 7930
rect 940 7870 950 7930
rect 870 7860 950 7870
rect 520 7800 580 7820
rect 520 7760 530 7800
rect 570 7760 580 7800
rect 520 7700 580 7760
rect 520 7660 530 7700
rect 570 7660 580 7700
rect 520 7580 580 7660
rect 640 7800 700 7820
rect 640 7760 650 7800
rect 690 7760 700 7800
rect 640 7700 700 7760
rect 640 7660 650 7700
rect 690 7660 700 7700
rect 640 7600 700 7660
rect 760 7800 820 7820
rect 760 7760 770 7800
rect 810 7760 820 7800
rect 760 7700 820 7760
rect 760 7660 770 7700
rect 810 7660 820 7700
rect 520 7540 530 7580
rect 570 7540 580 7580
rect 520 7490 580 7540
rect 630 7590 710 7600
rect 630 7530 640 7590
rect 700 7530 710 7590
rect 630 7520 710 7530
rect 760 7490 820 7660
rect 880 7800 940 7860
rect 880 7760 890 7800
rect 930 7760 940 7800
rect 880 7700 940 7760
rect 880 7660 890 7700
rect 930 7660 940 7700
rect 880 7640 940 7660
rect 1000 7800 1060 7820
rect 1000 7760 1010 7800
rect 1050 7760 1060 7800
rect 1000 7700 1060 7760
rect 1000 7660 1010 7700
rect 1050 7660 1060 7700
rect 1000 7490 1060 7660
rect 1120 7800 1180 7980
rect 1360 7920 1420 7980
rect 1360 7880 1370 7920
rect 1410 7880 1420 7920
rect 1360 7860 1420 7880
rect 1590 7930 1670 8370
rect 1850 8330 1890 8580
rect 2004 8532 2062 8540
rect 2004 8480 2008 8532
rect 2060 8480 2062 8532
rect 2004 8470 2062 8480
rect 2090 8440 2130 8580
rect 2158 8532 2216 8540
rect 2158 8480 2162 8532
rect 2214 8480 2216 8532
rect 2158 8470 2216 8480
rect 2070 8430 2150 8440
rect 2070 8370 2080 8430
rect 2140 8370 2150 8430
rect 2070 8360 2150 8370
rect 2330 8330 2370 8580
rect 2482 8532 2540 8540
rect 2482 8480 2486 8532
rect 2538 8480 2540 8532
rect 2482 8470 2540 8480
rect 2570 8440 2610 8580
rect 2790 8520 2800 8580
rect 2860 8520 2870 8580
rect 2790 8510 2870 8520
rect 2550 8430 2630 8440
rect 2550 8370 2560 8430
rect 2620 8370 2630 8430
rect 2550 8360 2630 8370
rect 1830 8320 1910 8330
rect 1830 8260 1840 8320
rect 1900 8260 1910 8320
rect 1830 8250 1910 8260
rect 2310 8320 2390 8330
rect 2310 8260 2320 8320
rect 2380 8260 2390 8320
rect 2310 8250 2390 8260
rect 1830 8050 1910 8060
rect 1830 7990 1840 8050
rect 1900 7990 1910 8050
rect 1830 7980 1910 7990
rect 2070 8050 2150 8060
rect 2070 7990 2080 8050
rect 2140 7990 2150 8050
rect 2070 7980 2150 7990
rect 2550 8050 2630 8060
rect 2550 7990 2560 8050
rect 2620 7990 2630 8050
rect 2550 7980 2630 7990
rect 2730 8050 2810 8060
rect 2730 7990 2740 8050
rect 2800 7990 2810 8050
rect 2730 7980 2810 7990
rect 1590 7870 1600 7930
rect 1660 7870 1670 7930
rect 1590 7860 1670 7870
rect 1120 7760 1130 7800
rect 1170 7760 1180 7800
rect 1120 7700 1180 7760
rect 1120 7660 1130 7700
rect 1170 7660 1180 7700
rect 1120 7640 1180 7660
rect 1240 7800 1300 7820
rect 1240 7760 1250 7800
rect 1290 7760 1300 7800
rect 1240 7700 1300 7760
rect 1240 7660 1250 7700
rect 1290 7660 1300 7700
rect 1240 7490 1300 7660
rect 1360 7800 1420 7820
rect 1360 7760 1370 7800
rect 1410 7760 1420 7800
rect 1360 7700 1420 7760
rect 1360 7660 1370 7700
rect 1410 7660 1420 7700
rect 1360 7600 1420 7660
rect 1480 7800 1540 7820
rect 1480 7760 1490 7800
rect 1530 7760 1540 7800
rect 1480 7700 1540 7760
rect 1480 7660 1490 7700
rect 1530 7660 1540 7700
rect 1350 7590 1430 7600
rect 1350 7530 1360 7590
rect 1420 7530 1430 7590
rect 1350 7520 1430 7530
rect 1480 7490 1540 7660
rect 1600 7800 1660 7860
rect 1600 7760 1610 7800
rect 1650 7760 1660 7800
rect 1600 7700 1660 7760
rect 1600 7660 1610 7700
rect 1650 7660 1660 7700
rect 1600 7640 1660 7660
rect 1720 7800 1780 7820
rect 1720 7760 1730 7800
rect 1770 7760 1780 7800
rect 1720 7700 1780 7760
rect 1720 7660 1730 7700
rect 1770 7660 1780 7700
rect 1720 7490 1780 7660
rect 1840 7800 1900 7980
rect 2080 7920 2140 7980
rect 2080 7880 2090 7920
rect 2130 7880 2140 7920
rect 2080 7860 2140 7880
rect 2310 7930 2390 7940
rect 2310 7870 2320 7930
rect 2380 7870 2390 7930
rect 2310 7860 2390 7870
rect 1840 7760 1850 7800
rect 1890 7760 1900 7800
rect 1840 7700 1900 7760
rect 1840 7660 1850 7700
rect 1890 7660 1900 7700
rect 1840 7640 1900 7660
rect 1960 7800 2020 7820
rect 1960 7760 1970 7800
rect 2010 7760 2020 7800
rect 1960 7700 2020 7760
rect 1960 7660 1970 7700
rect 2010 7660 2020 7700
rect 1960 7490 2020 7660
rect 2080 7800 2140 7820
rect 2080 7760 2090 7800
rect 2130 7760 2140 7800
rect 2080 7700 2140 7760
rect 2080 7660 2090 7700
rect 2130 7660 2140 7700
rect 2080 7600 2140 7660
rect 2200 7800 2260 7820
rect 2200 7760 2210 7800
rect 2250 7760 2260 7800
rect 2200 7700 2260 7760
rect 2200 7660 2210 7700
rect 2250 7660 2260 7700
rect 2070 7590 2150 7600
rect 2070 7530 2080 7590
rect 2140 7530 2150 7590
rect 2070 7520 2150 7530
rect 2200 7490 2260 7660
rect 2320 7800 2380 7860
rect 2320 7760 2330 7800
rect 2370 7760 2380 7800
rect 2320 7700 2380 7760
rect 2320 7660 2330 7700
rect 2370 7660 2380 7700
rect 2320 7640 2380 7660
rect 2440 7800 2500 7820
rect 2440 7760 2450 7800
rect 2490 7760 2500 7800
rect 2440 7700 2500 7760
rect 2440 7660 2450 7700
rect 2490 7660 2500 7700
rect 2440 7490 2500 7660
rect 2560 7800 2620 7980
rect 2740 7920 2800 7980
rect 2740 7880 2750 7920
rect 2790 7880 2800 7920
rect 2740 7860 2800 7880
rect 2560 7760 2570 7800
rect 2610 7760 2620 7800
rect 2560 7700 2620 7760
rect 2560 7660 2570 7700
rect 2610 7660 2620 7700
rect 2560 7640 2620 7660
rect 2680 7800 2740 7820
rect 2680 7760 2690 7800
rect 2730 7760 2740 7800
rect 2680 7700 2740 7760
rect 2680 7660 2690 7700
rect 2730 7660 2740 7700
rect 2680 7490 2740 7660
rect 2800 7800 2860 7820
rect 2800 7760 2810 7800
rect 2850 7760 2860 7800
rect 2800 7700 2860 7760
rect 2800 7660 2810 7700
rect 2850 7660 2860 7700
rect 2800 7600 2860 7660
rect 2920 7800 2980 7820
rect 2920 7760 2930 7800
rect 2970 7760 2980 7800
rect 2920 7700 2980 7760
rect 2920 7660 2930 7700
rect 2970 7660 2980 7700
rect 2790 7590 2870 7600
rect 2790 7530 2800 7590
rect 2860 7530 2870 7590
rect 2790 7520 2870 7530
rect 2920 7580 2980 7660
rect 3060 7600 3120 9120
rect 3150 8740 3390 9720
rect 4570 9940 4650 9950
rect 4570 9880 4580 9940
rect 4640 9880 4650 9940
rect 4570 9860 4650 9880
rect 4570 9800 4580 9860
rect 4640 9800 4650 9860
rect 4570 9780 4650 9800
rect 4570 9720 4580 9780
rect 4640 9720 4650 9780
rect 4570 9710 4650 9720
rect 5740 9650 5800 9670
rect 5740 9610 5750 9650
rect 5790 9610 5800 9650
rect 5740 9550 5800 9610
rect 5740 9510 5750 9550
rect 5790 9510 5800 9550
rect 5740 9450 5800 9510
rect 5740 9410 5750 9450
rect 5790 9410 5800 9450
rect 5740 9350 5800 9410
rect 5740 9310 5750 9350
rect 5790 9310 5800 9350
rect 5740 9250 5800 9310
rect 5740 9210 5750 9250
rect 5790 9210 5800 9250
rect 3150 8680 3160 8740
rect 3220 8680 3240 8740
rect 3300 8680 3320 8740
rect 3380 8680 3390 8740
rect 3150 8660 3390 8680
rect 3150 8600 3160 8660
rect 3220 8600 3240 8660
rect 3300 8600 3320 8660
rect 3380 8600 3390 8660
rect 3150 8580 3390 8600
rect 3150 8520 3160 8580
rect 3220 8520 3240 8580
rect 3300 8520 3320 8580
rect 3380 8520 3390 8580
rect 3150 8510 3390 8520
rect 3420 9160 3480 9180
rect 3420 9120 3430 9160
rect 3470 9120 3480 9160
rect 3420 7600 3480 9120
rect 3710 9140 3790 9150
rect 3710 9080 3720 9140
rect 3780 9080 3790 9140
rect 3710 9060 3790 9080
rect 3710 9000 3720 9060
rect 3780 9000 3790 9060
rect 3710 8980 3790 9000
rect 3710 8920 3720 8980
rect 3780 8920 3790 8980
rect 3710 8910 3790 8920
rect 3950 9140 4030 9150
rect 3950 9080 3960 9140
rect 4020 9080 4030 9140
rect 3950 9060 4030 9080
rect 3950 9000 3960 9060
rect 4020 9000 4030 9060
rect 3950 8980 4030 9000
rect 3950 8920 3960 8980
rect 4020 8920 4030 8980
rect 3950 8910 4030 8920
rect 4190 9140 4270 9150
rect 4190 9080 4200 9140
rect 4260 9080 4270 9140
rect 4190 9060 4270 9080
rect 4190 9000 4200 9060
rect 4260 9000 4270 9060
rect 4190 8980 4270 9000
rect 4190 8920 4200 8980
rect 4260 8920 4270 8980
rect 4190 8910 4270 8920
rect 4830 9140 4910 9150
rect 4830 9080 4840 9140
rect 4900 9080 4910 9140
rect 4830 9060 4910 9080
rect 4830 9000 4840 9060
rect 4900 9000 4910 9060
rect 4830 8980 4910 9000
rect 4830 8920 4840 8980
rect 4900 8920 4910 8980
rect 4830 8910 4910 8920
rect 5070 9140 5150 9150
rect 5070 9080 5080 9140
rect 5140 9080 5150 9140
rect 5070 9060 5150 9080
rect 5070 9000 5080 9060
rect 5140 9000 5150 9060
rect 5070 8980 5150 9000
rect 5070 8920 5080 8980
rect 5140 8920 5150 8980
rect 5070 8910 5150 8920
rect 5310 9140 5390 9150
rect 5310 9080 5320 9140
rect 5380 9080 5390 9140
rect 5310 9060 5390 9080
rect 5310 9000 5320 9060
rect 5380 9000 5390 9060
rect 5310 8980 5390 9000
rect 5310 8920 5320 8980
rect 5380 8920 5390 8980
rect 5310 8910 5390 8920
rect 5550 9140 5630 9150
rect 5550 9080 5560 9140
rect 5620 9080 5630 9140
rect 5550 9060 5630 9080
rect 5550 9000 5560 9060
rect 5620 9000 5630 9060
rect 5550 8980 5630 9000
rect 5550 8920 5560 8980
rect 5620 8920 5630 8980
rect 5550 8910 5630 8920
rect 5740 8880 5800 9210
rect 4020 8870 4100 8880
rect 4020 8810 4030 8870
rect 4090 8810 4100 8870
rect 4020 8800 4100 8810
rect 4280 8870 4360 8880
rect 4280 8810 4290 8870
rect 4350 8810 4360 8870
rect 4280 8800 4360 8810
rect 4500 8870 4580 8880
rect 4500 8810 4510 8870
rect 4570 8810 4580 8870
rect 4500 8800 4580 8810
rect 4760 8870 4840 8880
rect 4760 8810 4770 8870
rect 4830 8810 4840 8870
rect 4760 8800 4840 8810
rect 4980 8870 5060 8880
rect 4980 8810 4990 8870
rect 5050 8810 5060 8870
rect 4980 8800 5060 8810
rect 5730 8870 5810 8880
rect 5730 8810 5740 8870
rect 5800 8810 5810 8870
rect 5730 8800 5810 8810
rect 3670 8740 3750 8750
rect 3670 8680 3680 8740
rect 3740 8680 3750 8740
rect 3670 8660 3750 8680
rect 4040 8660 4070 8800
rect 4101 8760 4159 8770
rect 4101 8708 4105 8760
rect 4157 8708 4159 8760
rect 4101 8700 4159 8708
rect 4221 8760 4279 8770
rect 4221 8708 4225 8760
rect 4277 8708 4279 8760
rect 4221 8700 4279 8708
rect 4310 8660 4340 8800
rect 4520 8660 4550 8800
rect 4581 8760 4639 8770
rect 4581 8708 4585 8760
rect 4637 8708 4639 8760
rect 4581 8700 4639 8708
rect 4701 8760 4759 8770
rect 4701 8708 4705 8760
rect 4757 8708 4759 8760
rect 4701 8700 4759 8708
rect 4790 8660 4820 8800
rect 5000 8660 5030 8800
rect 6160 8770 6200 10540
rect 5061 8760 5119 8770
rect 5061 8708 5065 8760
rect 5117 8708 5119 8760
rect 5061 8700 5119 8708
rect 6140 8760 6220 8770
rect 6140 8700 6150 8760
rect 6210 8700 6220 8760
rect 6140 8690 6220 8700
rect 3670 8600 3680 8660
rect 3740 8600 3750 8660
rect 3670 8580 3750 8600
rect 3920 8640 3980 8660
rect 3920 8600 3930 8640
rect 3970 8600 3980 8640
rect 3920 8580 3980 8600
rect 4040 8640 4100 8660
rect 4040 8600 4050 8640
rect 4090 8600 4100 8640
rect 4040 8580 4100 8600
rect 4160 8640 4220 8660
rect 4160 8600 4170 8640
rect 4210 8600 4220 8640
rect 4160 8580 4220 8600
rect 4280 8640 4340 8660
rect 4280 8600 4290 8640
rect 4330 8600 4340 8640
rect 4280 8580 4340 8600
rect 4400 8640 4460 8660
rect 4400 8600 4410 8640
rect 4450 8600 4460 8640
rect 4400 8580 4460 8600
rect 4520 8640 4580 8660
rect 4520 8600 4530 8640
rect 4570 8600 4580 8640
rect 4520 8580 4580 8600
rect 4640 8640 4700 8660
rect 4640 8600 4650 8640
rect 4690 8600 4700 8640
rect 4640 8580 4700 8600
rect 4760 8640 4820 8660
rect 4760 8600 4770 8640
rect 4810 8600 4820 8640
rect 4760 8580 4820 8600
rect 4880 8640 4940 8660
rect 4880 8600 4890 8640
rect 4930 8600 4940 8640
rect 4880 8580 4940 8600
rect 5000 8640 5060 8660
rect 5000 8600 5010 8640
rect 5050 8600 5060 8640
rect 5000 8580 5060 8600
rect 5120 8640 5180 8660
rect 5120 8600 5130 8640
rect 5170 8600 5180 8640
rect 3670 8520 3680 8580
rect 3740 8520 3750 8580
rect 3670 8510 3750 8520
rect 3930 8440 3970 8580
rect 4000 8532 4058 8540
rect 4000 8480 4002 8532
rect 4054 8480 4058 8532
rect 4000 8470 4058 8480
rect 3910 8430 3990 8440
rect 3910 8370 3920 8430
rect 3980 8370 3990 8430
rect 3910 8360 3990 8370
rect 4170 8330 4210 8580
rect 4324 8532 4382 8540
rect 4324 8480 4326 8532
rect 4378 8480 4382 8532
rect 4324 8470 4382 8480
rect 4410 8440 4450 8580
rect 4478 8532 4536 8540
rect 4478 8480 4480 8532
rect 4532 8480 4536 8532
rect 4478 8470 4536 8480
rect 4390 8430 4470 8440
rect 4390 8370 4400 8430
rect 4460 8370 4470 8430
rect 4390 8360 4470 8370
rect 4650 8330 4690 8580
rect 4802 8532 4860 8540
rect 4802 8480 4804 8532
rect 4856 8480 4860 8532
rect 4802 8470 4860 8480
rect 4890 8440 4930 8580
rect 4960 8532 5018 8540
rect 4960 8480 4962 8532
rect 5014 8480 5018 8532
rect 4960 8470 5018 8480
rect 4870 8430 4950 8440
rect 4870 8370 4880 8430
rect 4940 8370 4950 8430
rect 4150 8320 4230 8330
rect 4150 8260 4160 8320
rect 4220 8260 4230 8320
rect 4150 8250 4230 8260
rect 4630 8320 4710 8330
rect 4630 8260 4640 8320
rect 4700 8260 4710 8320
rect 4630 8250 4710 8260
rect 3730 8210 3810 8220
rect 3730 8150 3740 8210
rect 3800 8150 3810 8210
rect 3730 8130 3810 8150
rect 3730 8070 3740 8130
rect 3800 8070 3810 8130
rect 3730 8050 3810 8070
rect 3730 7990 3740 8050
rect 3800 7990 3810 8050
rect 3730 7980 3810 7990
rect 3910 8210 3990 8220
rect 3910 8150 3920 8210
rect 3980 8150 3990 8210
rect 3910 8130 3990 8150
rect 3910 8070 3920 8130
rect 3980 8070 3990 8130
rect 3910 8050 3990 8070
rect 3910 7990 3920 8050
rect 3980 7990 3990 8050
rect 3910 7980 3990 7990
rect 4150 8210 4230 8220
rect 4150 8150 4160 8210
rect 4220 8150 4230 8210
rect 4150 8130 4230 8150
rect 4150 8070 4160 8130
rect 4220 8070 4230 8130
rect 4150 8050 4230 8070
rect 4150 7990 4160 8050
rect 4220 7990 4230 8050
rect 4150 7980 4230 7990
rect 4390 8210 4470 8220
rect 4390 8150 4400 8210
rect 4460 8150 4470 8210
rect 4390 8130 4470 8150
rect 4390 8070 4400 8130
rect 4460 8070 4470 8130
rect 4390 8050 4470 8070
rect 4390 7990 4400 8050
rect 4460 7990 4470 8050
rect 4390 7980 4470 7990
rect 4630 8210 4710 8220
rect 4630 8150 4640 8210
rect 4700 8150 4710 8210
rect 4630 8130 4710 8150
rect 4630 8070 4640 8130
rect 4700 8070 4710 8130
rect 4630 8050 4710 8070
rect 4630 7990 4640 8050
rect 4700 7990 4710 8050
rect 4630 7980 4710 7990
rect 3740 7920 3800 7980
rect 3740 7880 3750 7920
rect 3790 7880 3800 7920
rect 3740 7860 3800 7880
rect 3560 7800 3620 7820
rect 3560 7760 3570 7800
rect 3610 7760 3620 7800
rect 3560 7700 3620 7760
rect 3560 7660 3570 7700
rect 3610 7660 3620 7700
rect 2920 7540 2930 7580
rect 2970 7540 2980 7580
rect 2920 7490 2980 7540
rect 3050 7590 3130 7600
rect 3050 7530 3060 7590
rect 3120 7530 3130 7590
rect 3050 7520 3130 7530
rect 3410 7590 3490 7600
rect 3410 7530 3420 7590
rect 3480 7530 3490 7590
rect 510 7480 590 7490
rect 510 7420 520 7480
rect 580 7420 590 7480
rect 510 7400 590 7420
rect 510 7340 520 7400
rect 580 7340 590 7400
rect 510 7320 590 7340
rect 510 7260 520 7320
rect 580 7260 590 7320
rect 510 7250 590 7260
rect 750 7480 830 7490
rect 750 7420 760 7480
rect 820 7420 830 7480
rect 750 7400 830 7420
rect 750 7340 760 7400
rect 820 7340 830 7400
rect 750 7320 830 7340
rect 750 7260 760 7320
rect 820 7260 830 7320
rect 750 7250 830 7260
rect 990 7480 1070 7490
rect 990 7420 1000 7480
rect 1060 7420 1070 7480
rect 990 7400 1070 7420
rect 990 7340 1000 7400
rect 1060 7340 1070 7400
rect 990 7320 1070 7340
rect 990 7260 1000 7320
rect 1060 7260 1070 7320
rect 990 7250 1070 7260
rect 1230 7480 1310 7490
rect 1230 7420 1240 7480
rect 1300 7420 1310 7480
rect 1230 7400 1310 7420
rect 1230 7340 1240 7400
rect 1300 7340 1310 7400
rect 1230 7320 1310 7340
rect 1230 7260 1240 7320
rect 1300 7260 1310 7320
rect 1230 7250 1310 7260
rect 1470 7480 1550 7490
rect 1470 7420 1480 7480
rect 1540 7420 1550 7480
rect 1470 7400 1550 7420
rect 1470 7340 1480 7400
rect 1540 7340 1550 7400
rect 1470 7320 1550 7340
rect 1470 7260 1480 7320
rect 1540 7260 1550 7320
rect 1470 7250 1550 7260
rect 1710 7480 1790 7490
rect 1710 7420 1720 7480
rect 1780 7420 1790 7480
rect 1710 7400 1790 7420
rect 1710 7340 1720 7400
rect 1780 7340 1790 7400
rect 1710 7320 1790 7340
rect 1710 7260 1720 7320
rect 1780 7260 1790 7320
rect 1710 7250 1790 7260
rect 1950 7480 2030 7490
rect 1950 7420 1960 7480
rect 2020 7420 2030 7480
rect 1950 7400 2030 7420
rect 1950 7340 1960 7400
rect 2020 7340 2030 7400
rect 1950 7320 2030 7340
rect 1950 7260 1960 7320
rect 2020 7260 2030 7320
rect 1950 7250 2030 7260
rect 2190 7480 2270 7490
rect 2190 7420 2200 7480
rect 2260 7420 2270 7480
rect 2190 7400 2270 7420
rect 2190 7340 2200 7400
rect 2260 7340 2270 7400
rect 2190 7320 2270 7340
rect 2190 7260 2200 7320
rect 2260 7260 2270 7320
rect 2190 7250 2270 7260
rect 2430 7480 2510 7490
rect 2430 7420 2440 7480
rect 2500 7420 2510 7480
rect 2430 7400 2510 7420
rect 2430 7340 2440 7400
rect 2500 7340 2510 7400
rect 2430 7320 2510 7340
rect 2430 7260 2440 7320
rect 2500 7260 2510 7320
rect 2430 7250 2510 7260
rect 2670 7480 2750 7490
rect 2670 7420 2680 7480
rect 2740 7420 2750 7480
rect 2670 7400 2750 7420
rect 2670 7340 2680 7400
rect 2740 7340 2750 7400
rect 2670 7320 2750 7340
rect 2670 7260 2680 7320
rect 2740 7260 2750 7320
rect 2670 7250 2750 7260
rect 2910 7480 2990 7490
rect 2910 7420 2920 7480
rect 2980 7420 2990 7480
rect 2910 7400 2990 7420
rect 2910 7340 2920 7400
rect 2980 7340 2990 7400
rect 2910 7320 2990 7340
rect 2910 7260 2920 7320
rect 2980 7260 2990 7320
rect 2910 7250 2990 7260
rect 1790 7210 1870 7220
rect 1790 7150 1800 7210
rect 1860 7150 1870 7210
rect 1790 7140 1870 7150
rect 3230 7210 3310 7220
rect 3230 7150 3240 7210
rect 3300 7150 3310 7210
rect 3230 7140 3310 7150
rect 1620 6640 1680 6660
rect 1620 6600 1630 6640
rect 1670 6600 1680 6640
rect 1620 6540 1680 6600
rect 1620 6500 1630 6540
rect 1670 6500 1680 6540
rect 1620 6440 1680 6500
rect 1620 6400 1630 6440
rect 1670 6400 1680 6440
rect 1620 6340 1680 6400
rect 1620 6300 1630 6340
rect 1670 6300 1680 6340
rect 1620 6240 1680 6300
rect 1620 6200 1630 6240
rect 1670 6200 1680 6240
rect 1620 6140 1680 6200
rect 1620 6100 1630 6140
rect 1670 6100 1680 6140
rect 1620 6080 1680 6100
rect 1800 6640 1860 7140
rect 2150 7100 2230 7110
rect 2150 7040 2160 7100
rect 2220 7040 2230 7100
rect 2150 7030 2230 7040
rect 1890 6770 1960 6780
rect 1950 6710 1960 6770
rect 1890 6700 1960 6710
rect 2060 6770 2140 6780
rect 2060 6710 2070 6770
rect 2130 6710 2140 6770
rect 2060 6700 2140 6710
rect 2170 6660 2210 7030
rect 2510 6990 2590 7000
rect 2510 6930 2520 6990
rect 2580 6930 2590 6990
rect 2510 6920 2590 6930
rect 2240 6770 2320 6780
rect 2240 6710 2250 6770
rect 2310 6710 2320 6770
rect 2240 6700 2320 6710
rect 2420 6770 2500 6780
rect 2420 6710 2430 6770
rect 2490 6710 2500 6770
rect 2420 6700 2500 6710
rect 2530 6660 2570 6920
rect 2870 6880 2950 6890
rect 2870 6820 2880 6880
rect 2940 6820 2950 6880
rect 2870 6810 2950 6820
rect 2600 6770 2680 6780
rect 2600 6710 2610 6770
rect 2670 6710 2680 6770
rect 2600 6700 2680 6710
rect 2780 6770 2860 6780
rect 2780 6710 2790 6770
rect 2850 6710 2860 6770
rect 2780 6700 2860 6710
rect 2890 6660 2930 6810
rect 2960 6770 3040 6780
rect 2960 6710 2970 6770
rect 3030 6710 3040 6770
rect 2960 6700 3040 6710
rect 3140 6770 3210 6780
rect 3140 6710 3150 6770
rect 3140 6700 3210 6710
rect 1800 6600 1810 6640
rect 1850 6600 1860 6640
rect 1800 6540 1860 6600
rect 1800 6500 1810 6540
rect 1850 6500 1860 6540
rect 1800 6440 1860 6500
rect 1800 6400 1810 6440
rect 1850 6400 1860 6440
rect 1800 6340 1860 6400
rect 1800 6300 1810 6340
rect 1850 6300 1860 6340
rect 1800 6240 1860 6300
rect 1800 6200 1810 6240
rect 1850 6200 1860 6240
rect 1800 6140 1860 6200
rect 1800 6100 1810 6140
rect 1850 6100 1860 6140
rect 1800 6080 1860 6100
rect 1980 6640 2040 6660
rect 1980 6600 1990 6640
rect 2030 6600 2040 6640
rect 1980 6540 2040 6600
rect 1980 6500 1990 6540
rect 2030 6500 2040 6540
rect 1980 6440 2040 6500
rect 1980 6400 1990 6440
rect 2030 6400 2040 6440
rect 1980 6340 2040 6400
rect 1980 6300 1990 6340
rect 2030 6300 2040 6340
rect 1980 6240 2040 6300
rect 1980 6200 1990 6240
rect 2030 6200 2040 6240
rect 1980 6140 2040 6200
rect 1980 6100 1990 6140
rect 2030 6100 2040 6140
rect 1980 6080 2040 6100
rect 2160 6640 2220 6660
rect 2160 6600 2170 6640
rect 2210 6600 2220 6640
rect 2160 6540 2220 6600
rect 2160 6500 2170 6540
rect 2210 6500 2220 6540
rect 2160 6440 2220 6500
rect 2160 6400 2170 6440
rect 2210 6400 2220 6440
rect 2160 6340 2220 6400
rect 2160 6300 2170 6340
rect 2210 6300 2220 6340
rect 2160 6240 2220 6300
rect 2160 6200 2170 6240
rect 2210 6200 2220 6240
rect 2160 6140 2220 6200
rect 2160 6100 2170 6140
rect 2210 6100 2220 6140
rect 2160 6080 2220 6100
rect 2340 6640 2400 6660
rect 2340 6600 2350 6640
rect 2390 6600 2400 6640
rect 2340 6540 2400 6600
rect 2340 6500 2350 6540
rect 2390 6500 2400 6540
rect 2340 6440 2400 6500
rect 2340 6400 2350 6440
rect 2390 6400 2400 6440
rect 2340 6340 2400 6400
rect 2340 6300 2350 6340
rect 2390 6300 2400 6340
rect 2340 6240 2400 6300
rect 2340 6200 2350 6240
rect 2390 6200 2400 6240
rect 2340 6140 2400 6200
rect 2340 6100 2350 6140
rect 2390 6100 2400 6140
rect 2340 6080 2400 6100
rect 2520 6640 2580 6660
rect 2520 6600 2530 6640
rect 2570 6600 2580 6640
rect 2520 6540 2580 6600
rect 2520 6500 2530 6540
rect 2570 6500 2580 6540
rect 2520 6440 2580 6500
rect 2520 6400 2530 6440
rect 2570 6400 2580 6440
rect 2520 6340 2580 6400
rect 2520 6300 2530 6340
rect 2570 6300 2580 6340
rect 2520 6240 2580 6300
rect 2520 6200 2530 6240
rect 2570 6200 2580 6240
rect 2520 6140 2580 6200
rect 2520 6100 2530 6140
rect 2570 6100 2580 6140
rect 2520 6080 2580 6100
rect 2700 6640 2760 6660
rect 2700 6600 2710 6640
rect 2750 6600 2760 6640
rect 2700 6540 2760 6600
rect 2700 6500 2710 6540
rect 2750 6500 2760 6540
rect 2700 6440 2760 6500
rect 2700 6400 2710 6440
rect 2750 6400 2760 6440
rect 2700 6340 2760 6400
rect 2700 6300 2710 6340
rect 2750 6300 2760 6340
rect 2700 6240 2760 6300
rect 2700 6200 2710 6240
rect 2750 6200 2760 6240
rect 2700 6140 2760 6200
rect 2700 6100 2710 6140
rect 2750 6100 2760 6140
rect 2700 6080 2760 6100
rect 2880 6640 2940 6660
rect 2880 6600 2890 6640
rect 2930 6600 2940 6640
rect 2880 6540 2940 6600
rect 2880 6500 2890 6540
rect 2930 6500 2940 6540
rect 2880 6440 2940 6500
rect 2880 6400 2890 6440
rect 2930 6400 2940 6440
rect 2880 6340 2940 6400
rect 2880 6300 2890 6340
rect 2930 6300 2940 6340
rect 2880 6240 2940 6300
rect 2880 6200 2890 6240
rect 2930 6200 2940 6240
rect 2880 6140 2940 6200
rect 2880 6100 2890 6140
rect 2930 6100 2940 6140
rect 2880 6080 2940 6100
rect 3060 6640 3120 6660
rect 3060 6600 3070 6640
rect 3110 6600 3120 6640
rect 3060 6540 3120 6600
rect 3060 6500 3070 6540
rect 3110 6500 3120 6540
rect 3060 6440 3120 6500
rect 3060 6400 3070 6440
rect 3110 6400 3120 6440
rect 3060 6340 3120 6400
rect 3060 6300 3070 6340
rect 3110 6300 3120 6340
rect 3060 6240 3120 6300
rect 3060 6200 3070 6240
rect 3110 6200 3120 6240
rect 3060 6140 3120 6200
rect 3060 6100 3070 6140
rect 3110 6100 3120 6140
rect 3060 6080 3120 6100
rect 3240 6640 3300 7140
rect 3410 6780 3490 7530
rect 3560 7580 3620 7660
rect 3680 7800 3740 7820
rect 3680 7760 3690 7800
rect 3730 7760 3740 7800
rect 3680 7700 3740 7760
rect 3680 7660 3690 7700
rect 3730 7660 3740 7700
rect 3680 7600 3740 7660
rect 3800 7800 3860 7820
rect 3800 7760 3810 7800
rect 3850 7760 3860 7800
rect 3800 7700 3860 7760
rect 3800 7660 3810 7700
rect 3850 7660 3860 7700
rect 3560 7540 3570 7580
rect 3610 7540 3620 7580
rect 3560 7490 3620 7540
rect 3670 7590 3750 7600
rect 3670 7530 3680 7590
rect 3740 7530 3750 7590
rect 3670 7520 3750 7530
rect 3800 7490 3860 7660
rect 3920 7800 3980 7980
rect 4150 7930 4230 7940
rect 4150 7870 4160 7930
rect 4220 7870 4230 7930
rect 4150 7860 4230 7870
rect 4400 7920 4460 7980
rect 4400 7880 4410 7920
rect 4450 7880 4460 7920
rect 4400 7860 4460 7880
rect 3920 7760 3930 7800
rect 3970 7760 3980 7800
rect 3920 7700 3980 7760
rect 3920 7660 3930 7700
rect 3970 7660 3980 7700
rect 3920 7640 3980 7660
rect 4040 7800 4100 7820
rect 4040 7760 4050 7800
rect 4090 7760 4100 7800
rect 4040 7700 4100 7760
rect 4040 7660 4050 7700
rect 4090 7660 4100 7700
rect 4040 7490 4100 7660
rect 4160 7800 4220 7860
rect 4160 7760 4170 7800
rect 4210 7760 4220 7800
rect 4160 7700 4220 7760
rect 4160 7660 4170 7700
rect 4210 7660 4220 7700
rect 4160 7640 4220 7660
rect 4280 7800 4340 7820
rect 4280 7760 4290 7800
rect 4330 7760 4340 7800
rect 4280 7700 4340 7760
rect 4280 7660 4290 7700
rect 4330 7660 4340 7700
rect 4280 7490 4340 7660
rect 4400 7800 4460 7820
rect 4400 7760 4410 7800
rect 4450 7760 4460 7800
rect 4400 7700 4460 7760
rect 4400 7660 4410 7700
rect 4450 7660 4460 7700
rect 4400 7600 4460 7660
rect 4520 7800 4580 7820
rect 4520 7760 4530 7800
rect 4570 7760 4580 7800
rect 4520 7700 4580 7760
rect 4520 7660 4530 7700
rect 4570 7660 4580 7700
rect 4390 7590 4470 7600
rect 4390 7530 4400 7590
rect 4460 7530 4470 7590
rect 4390 7520 4470 7530
rect 4520 7490 4580 7660
rect 4640 7800 4700 7980
rect 4870 7930 4950 8370
rect 5120 8330 5180 8600
rect 5110 8320 5190 8330
rect 5110 8260 5120 8320
rect 5180 8260 5190 8320
rect 5110 8210 5190 8260
rect 5110 8150 5120 8210
rect 5180 8150 5190 8210
rect 5110 8130 5190 8150
rect 5110 8070 5120 8130
rect 5180 8070 5190 8130
rect 5110 8050 5190 8070
rect 5110 7990 5120 8050
rect 5180 7990 5190 8050
rect 5110 7980 5190 7990
rect 5350 8210 5430 8220
rect 5350 8150 5360 8210
rect 5420 8150 5430 8210
rect 5350 8130 5430 8150
rect 5350 8070 5360 8130
rect 5420 8070 5430 8130
rect 5350 8050 5430 8070
rect 5350 7990 5360 8050
rect 5420 7990 5430 8050
rect 5350 7980 5430 7990
rect 5770 8210 5850 8220
rect 5770 8150 5780 8210
rect 5840 8150 5850 8210
rect 5770 8130 5850 8150
rect 5770 8070 5780 8130
rect 5840 8070 5850 8130
rect 5770 8050 5850 8070
rect 5770 7990 5780 8050
rect 5840 7990 5850 8050
rect 5770 7980 5850 7990
rect 4870 7870 4880 7930
rect 4940 7870 4950 7930
rect 4870 7860 4950 7870
rect 5120 7920 5180 7980
rect 5120 7880 5130 7920
rect 5170 7880 5180 7920
rect 5120 7860 5180 7880
rect 4640 7760 4650 7800
rect 4690 7760 4700 7800
rect 4640 7700 4700 7760
rect 4640 7660 4650 7700
rect 4690 7660 4700 7700
rect 4640 7640 4700 7660
rect 4760 7800 4820 7820
rect 4760 7760 4770 7800
rect 4810 7760 4820 7800
rect 4760 7700 4820 7760
rect 4760 7660 4770 7700
rect 4810 7660 4820 7700
rect 4760 7490 4820 7660
rect 4880 7800 4940 7860
rect 4880 7760 4890 7800
rect 4930 7760 4940 7800
rect 4880 7700 4940 7760
rect 4880 7660 4890 7700
rect 4930 7660 4940 7700
rect 4880 7640 4940 7660
rect 5000 7800 5060 7820
rect 5000 7760 5010 7800
rect 5050 7760 5060 7800
rect 5000 7700 5060 7760
rect 5000 7660 5010 7700
rect 5050 7660 5060 7700
rect 5000 7490 5060 7660
rect 5120 7800 5180 7820
rect 5120 7760 5130 7800
rect 5170 7760 5180 7800
rect 5120 7700 5180 7760
rect 5120 7660 5130 7700
rect 5170 7660 5180 7700
rect 5120 7600 5180 7660
rect 5240 7800 5300 7820
rect 5240 7760 5250 7800
rect 5290 7760 5300 7800
rect 5240 7700 5300 7760
rect 5240 7660 5250 7700
rect 5290 7660 5300 7700
rect 5110 7590 5190 7600
rect 5110 7530 5120 7590
rect 5180 7530 5190 7590
rect 5110 7520 5190 7530
rect 5240 7490 5300 7660
rect 5360 7800 5420 7980
rect 5590 7930 5670 7940
rect 5590 7870 5600 7930
rect 5660 7870 5670 7930
rect 5780 7930 5840 7980
rect 5780 7890 5790 7930
rect 5830 7890 5840 7930
rect 5780 7870 5840 7890
rect 5590 7860 5670 7870
rect 5360 7760 5370 7800
rect 5410 7760 5420 7800
rect 5360 7700 5420 7760
rect 5360 7660 5370 7700
rect 5410 7660 5420 7700
rect 5360 7640 5420 7660
rect 5480 7800 5540 7820
rect 5480 7760 5490 7800
rect 5530 7760 5540 7800
rect 5480 7700 5540 7760
rect 5480 7660 5490 7700
rect 5530 7660 5540 7700
rect 5480 7490 5540 7660
rect 5600 7800 5660 7860
rect 5600 7760 5610 7800
rect 5650 7760 5660 7800
rect 5600 7700 5660 7760
rect 5600 7660 5610 7700
rect 5650 7660 5660 7700
rect 5600 7640 5660 7660
rect 5720 7800 5780 7820
rect 5720 7760 5730 7800
rect 5770 7760 5780 7800
rect 5720 7700 5780 7760
rect 5720 7660 5730 7700
rect 5770 7660 5780 7700
rect 5720 7490 5780 7660
rect 5840 7800 5900 7820
rect 5840 7760 5850 7800
rect 5890 7760 5900 7800
rect 5840 7700 5900 7760
rect 5840 7660 5850 7700
rect 5890 7660 5900 7700
rect 5840 7600 5900 7660
rect 5960 7800 6020 7820
rect 5960 7760 5970 7800
rect 6010 7760 6020 7800
rect 5960 7700 6020 7760
rect 5960 7660 5970 7700
rect 6010 7660 6020 7700
rect 5830 7590 5910 7600
rect 5830 7530 5840 7590
rect 5900 7530 5910 7590
rect 3550 7480 3630 7490
rect 3550 7420 3560 7480
rect 3620 7420 3630 7480
rect 3550 7400 3630 7420
rect 3550 7340 3560 7400
rect 3620 7340 3630 7400
rect 3550 7320 3630 7340
rect 3550 7260 3560 7320
rect 3620 7260 3630 7320
rect 3550 7250 3630 7260
rect 3790 7480 3870 7490
rect 3790 7420 3800 7480
rect 3860 7420 3870 7480
rect 3790 7400 3870 7420
rect 3790 7340 3800 7400
rect 3860 7340 3870 7400
rect 3790 7320 3870 7340
rect 3790 7260 3800 7320
rect 3860 7260 3870 7320
rect 3790 7250 3870 7260
rect 4030 7480 4110 7490
rect 4030 7420 4040 7480
rect 4100 7420 4110 7480
rect 4030 7400 4110 7420
rect 4030 7340 4040 7400
rect 4100 7340 4110 7400
rect 4030 7320 4110 7340
rect 4030 7260 4040 7320
rect 4100 7260 4110 7320
rect 4030 7250 4110 7260
rect 4270 7480 4350 7490
rect 4270 7420 4280 7480
rect 4340 7420 4350 7480
rect 4270 7400 4350 7420
rect 4270 7340 4280 7400
rect 4340 7340 4350 7400
rect 4270 7320 4350 7340
rect 4270 7260 4280 7320
rect 4340 7260 4350 7320
rect 4270 7250 4350 7260
rect 4510 7480 4590 7490
rect 4510 7420 4520 7480
rect 4580 7420 4590 7480
rect 4510 7400 4590 7420
rect 4510 7340 4520 7400
rect 4580 7340 4590 7400
rect 4510 7320 4590 7340
rect 4510 7260 4520 7320
rect 4580 7260 4590 7320
rect 4510 7250 4590 7260
rect 4750 7480 4830 7490
rect 4750 7420 4760 7480
rect 4820 7420 4830 7480
rect 4750 7400 4830 7420
rect 4750 7340 4760 7400
rect 4820 7340 4830 7400
rect 4750 7320 4830 7340
rect 4750 7260 4760 7320
rect 4820 7260 4830 7320
rect 4750 7250 4830 7260
rect 4990 7480 5070 7490
rect 4990 7420 5000 7480
rect 5060 7420 5070 7480
rect 4990 7400 5070 7420
rect 4990 7340 5000 7400
rect 5060 7340 5070 7400
rect 4990 7320 5070 7340
rect 4990 7260 5000 7320
rect 5060 7260 5070 7320
rect 4990 7250 5070 7260
rect 5230 7480 5310 7490
rect 5230 7420 5240 7480
rect 5300 7420 5310 7480
rect 5230 7400 5310 7420
rect 5230 7340 5240 7400
rect 5300 7340 5310 7400
rect 5230 7320 5310 7340
rect 5230 7260 5240 7320
rect 5300 7260 5310 7320
rect 5230 7250 5310 7260
rect 5470 7480 5550 7490
rect 5470 7420 5480 7480
rect 5540 7420 5550 7480
rect 5470 7400 5550 7420
rect 5470 7340 5480 7400
rect 5540 7340 5550 7400
rect 5470 7320 5550 7340
rect 5470 7260 5480 7320
rect 5540 7260 5550 7320
rect 5470 7250 5550 7260
rect 5710 7480 5790 7490
rect 5710 7420 5720 7480
rect 5780 7420 5790 7480
rect 5710 7400 5790 7420
rect 5710 7340 5720 7400
rect 5780 7340 5790 7400
rect 5710 7320 5790 7340
rect 5710 7260 5720 7320
rect 5780 7260 5790 7320
rect 5710 7250 5790 7260
rect 4670 7210 4750 7220
rect 4670 7150 4680 7210
rect 4740 7150 4750 7210
rect 4670 7140 4750 7150
rect 4310 7100 4390 7110
rect 4310 7040 4320 7100
rect 4380 7040 4390 7100
rect 4310 7030 4390 7040
rect 3950 6990 4030 7000
rect 3950 6930 3960 6990
rect 4020 6930 4030 6990
rect 3950 6920 4030 6930
rect 3590 6880 3670 6890
rect 3590 6820 3600 6880
rect 3660 6820 3670 6880
rect 3590 6810 3670 6820
rect 3330 6770 3580 6780
rect 3390 6710 3420 6770
rect 3480 6710 3510 6770
rect 3570 6710 3580 6770
rect 3330 6700 3580 6710
rect 3610 6660 3650 6810
rect 3680 6770 3760 6780
rect 3680 6710 3690 6770
rect 3750 6710 3760 6770
rect 3680 6700 3760 6710
rect 3860 6770 3940 6780
rect 3860 6710 3870 6770
rect 3930 6710 3940 6770
rect 3860 6700 3940 6710
rect 3970 6660 4010 6920
rect 4040 6770 4120 6780
rect 4040 6710 4050 6770
rect 4110 6710 4120 6770
rect 4040 6700 4120 6710
rect 4220 6770 4300 6780
rect 4220 6710 4230 6770
rect 4290 6710 4300 6770
rect 4220 6700 4300 6710
rect 4330 6660 4370 7030
rect 4400 6770 4480 6780
rect 4400 6710 4410 6770
rect 4470 6710 4480 6770
rect 4400 6700 4480 6710
rect 4580 6770 4650 6780
rect 4580 6710 4590 6770
rect 4580 6700 4650 6710
rect 3240 6600 3250 6640
rect 3290 6600 3300 6640
rect 3240 6540 3300 6600
rect 3240 6500 3250 6540
rect 3290 6500 3300 6540
rect 3240 6440 3300 6500
rect 3240 6400 3250 6440
rect 3290 6400 3300 6440
rect 3240 6340 3300 6400
rect 3240 6300 3250 6340
rect 3290 6300 3300 6340
rect 3240 6240 3300 6300
rect 3240 6200 3250 6240
rect 3290 6200 3300 6240
rect 3240 6140 3300 6200
rect 3240 6100 3250 6140
rect 3290 6100 3300 6140
rect 3240 6080 3300 6100
rect 3420 6640 3480 6660
rect 3420 6600 3430 6640
rect 3470 6600 3480 6640
rect 3420 6540 3480 6600
rect 3420 6500 3430 6540
rect 3470 6500 3480 6540
rect 3420 6440 3480 6500
rect 3420 6400 3430 6440
rect 3470 6400 3480 6440
rect 3420 6340 3480 6400
rect 3420 6300 3430 6340
rect 3470 6300 3480 6340
rect 3420 6240 3480 6300
rect 3420 6200 3430 6240
rect 3470 6200 3480 6240
rect 3420 6140 3480 6200
rect 3420 6100 3430 6140
rect 3470 6100 3480 6140
rect 3420 6080 3480 6100
rect 3600 6640 3660 6660
rect 3600 6600 3610 6640
rect 3650 6600 3660 6640
rect 3600 6540 3660 6600
rect 3600 6500 3610 6540
rect 3650 6500 3660 6540
rect 3600 6440 3660 6500
rect 3600 6400 3610 6440
rect 3650 6400 3660 6440
rect 3600 6340 3660 6400
rect 3600 6300 3610 6340
rect 3650 6300 3660 6340
rect 3600 6240 3660 6300
rect 3600 6200 3610 6240
rect 3650 6200 3660 6240
rect 3600 6140 3660 6200
rect 3600 6100 3610 6140
rect 3650 6100 3660 6140
rect 3600 6080 3660 6100
rect 3780 6640 3840 6660
rect 3780 6600 3790 6640
rect 3830 6600 3840 6640
rect 3780 6540 3840 6600
rect 3780 6500 3790 6540
rect 3830 6500 3840 6540
rect 3780 6440 3840 6500
rect 3780 6400 3790 6440
rect 3830 6400 3840 6440
rect 3780 6340 3840 6400
rect 3780 6300 3790 6340
rect 3830 6300 3840 6340
rect 3780 6240 3840 6300
rect 3780 6200 3790 6240
rect 3830 6200 3840 6240
rect 3780 6140 3840 6200
rect 3780 6100 3790 6140
rect 3830 6100 3840 6140
rect 3780 6080 3840 6100
rect 3960 6640 4020 6660
rect 3960 6600 3970 6640
rect 4010 6600 4020 6640
rect 3960 6540 4020 6600
rect 3960 6500 3970 6540
rect 4010 6500 4020 6540
rect 3960 6440 4020 6500
rect 3960 6400 3970 6440
rect 4010 6400 4020 6440
rect 3960 6340 4020 6400
rect 3960 6300 3970 6340
rect 4010 6300 4020 6340
rect 3960 6240 4020 6300
rect 3960 6200 3970 6240
rect 4010 6200 4020 6240
rect 3960 6140 4020 6200
rect 3960 6100 3970 6140
rect 4010 6100 4020 6140
rect 3960 6080 4020 6100
rect 4140 6640 4200 6660
rect 4140 6600 4150 6640
rect 4190 6600 4200 6640
rect 4140 6540 4200 6600
rect 4140 6500 4150 6540
rect 4190 6500 4200 6540
rect 4140 6440 4200 6500
rect 4140 6400 4150 6440
rect 4190 6400 4200 6440
rect 4140 6340 4200 6400
rect 4140 6300 4150 6340
rect 4190 6300 4200 6340
rect 4140 6240 4200 6300
rect 4140 6200 4150 6240
rect 4190 6200 4200 6240
rect 4140 6140 4200 6200
rect 4140 6100 4150 6140
rect 4190 6100 4200 6140
rect 4140 6080 4200 6100
rect 4320 6640 4380 6660
rect 4320 6600 4330 6640
rect 4370 6600 4380 6640
rect 4320 6540 4380 6600
rect 4320 6500 4330 6540
rect 4370 6500 4380 6540
rect 4320 6440 4380 6500
rect 4320 6400 4330 6440
rect 4370 6400 4380 6440
rect 4320 6340 4380 6400
rect 4320 6300 4330 6340
rect 4370 6300 4380 6340
rect 4320 6240 4380 6300
rect 4320 6200 4330 6240
rect 4370 6200 4380 6240
rect 4320 6140 4380 6200
rect 4320 6100 4330 6140
rect 4370 6100 4380 6140
rect 4320 6080 4380 6100
rect 4500 6640 4560 6660
rect 4500 6600 4510 6640
rect 4550 6600 4560 6640
rect 4500 6540 4560 6600
rect 4500 6500 4510 6540
rect 4550 6500 4560 6540
rect 4500 6440 4560 6500
rect 4500 6400 4510 6440
rect 4550 6400 4560 6440
rect 4500 6340 4560 6400
rect 4500 6300 4510 6340
rect 4550 6300 4560 6340
rect 4500 6240 4560 6300
rect 4500 6200 4510 6240
rect 4550 6200 4560 6240
rect 4500 6140 4560 6200
rect 4500 6100 4510 6140
rect 4550 6100 4560 6140
rect 4500 6080 4560 6100
rect 4680 6640 4740 7140
rect 5700 7100 5780 7110
rect 5700 7040 5710 7100
rect 5770 7040 5780 7100
rect 5230 6990 5310 7000
rect 5230 6930 5240 6990
rect 5300 6930 5310 6990
rect 5230 6920 5310 6930
rect 4680 6600 4690 6640
rect 4730 6600 4740 6640
rect 4680 6540 4740 6600
rect 4680 6500 4690 6540
rect 4730 6500 4740 6540
rect 4680 6440 4740 6500
rect 4680 6400 4690 6440
rect 4730 6400 4740 6440
rect 4680 6340 4740 6400
rect 4680 6300 4690 6340
rect 4730 6300 4740 6340
rect 4680 6240 4740 6300
rect 4680 6200 4690 6240
rect 4730 6200 4740 6240
rect 4680 6140 4740 6200
rect 4680 6100 4690 6140
rect 4730 6100 4740 6140
rect 4680 6080 4740 6100
rect 4860 6640 4920 6660
rect 4860 6600 4870 6640
rect 4910 6600 4920 6640
rect 4860 6540 4920 6600
rect 4860 6500 4870 6540
rect 4910 6500 4920 6540
rect 4860 6440 4920 6500
rect 4860 6400 4870 6440
rect 4910 6400 4920 6440
rect 4860 6340 4920 6400
rect 4860 6300 4870 6340
rect 4910 6300 4920 6340
rect 4860 6240 4920 6300
rect 5250 6240 5290 6920
rect 5580 6570 5660 6580
rect 5580 6510 5590 6570
rect 5650 6510 5660 6570
rect 5580 6500 5660 6510
rect 5700 6560 5780 7040
rect 5830 6580 5910 7530
rect 5960 7580 6020 7660
rect 5960 7540 5970 7580
rect 6010 7540 6020 7580
rect 5960 7490 6020 7540
rect 5950 7480 6030 7490
rect 5950 7420 5960 7480
rect 6020 7420 6030 7480
rect 5950 7400 6030 7420
rect 5950 7340 5960 7400
rect 6020 7340 6030 7400
rect 5950 7320 6030 7340
rect 5950 7260 5960 7320
rect 6020 7260 6030 7320
rect 5950 7250 6030 7260
rect 6160 6890 6200 8690
rect 6250 8540 6290 10740
rect 6230 8530 6310 8540
rect 6230 8470 6240 8530
rect 6300 8470 6310 8530
rect 6230 8460 6310 8470
rect 6250 7000 6290 8460
rect 6460 7590 6540 12700
rect 6840 12060 6920 14330
rect 6950 14160 7050 14180
rect 6950 14100 6970 14160
rect 7030 14100 7050 14160
rect 6950 14080 7050 14100
rect 6840 12000 6850 12060
rect 6910 12000 6920 12060
rect 6840 11990 6920 12000
rect 6570 11360 6810 11380
rect 6570 11300 6580 11360
rect 6640 11300 6660 11360
rect 6720 11300 6740 11360
rect 6800 11300 6810 11360
rect 6570 8210 6810 11300
rect 6960 10390 7040 14080
rect 7210 13460 7290 13470
rect 7210 13400 7220 13460
rect 7280 13400 7290 13460
rect 7070 12760 7170 12780
rect 7070 12700 7090 12760
rect 7150 12700 7170 12760
rect 7070 12680 7170 12700
rect 7070 11360 7170 11380
rect 7070 11300 7090 11360
rect 7150 11300 7170 11360
rect 7070 11280 7170 11300
rect 6960 10330 6970 10390
rect 7030 10330 7040 10390
rect 6960 10320 7040 10330
rect 7210 9150 7290 13400
rect 11750 9810 11850 9830
rect 11750 9750 11770 9810
rect 11830 9750 11850 9810
rect 11750 9730 11850 9750
rect 7200 9110 7300 9150
rect 7200 9050 7220 9110
rect 7280 9050 7300 9110
rect 7200 9010 7300 9050
rect 7200 8950 7220 9010
rect 7280 8950 7300 9010
rect 7200 8910 7300 8950
rect 8410 8580 8490 8600
rect 8410 8530 8430 8580
rect 8470 8530 8490 8580
rect 8410 8440 8490 8530
rect 8410 8390 8430 8440
rect 8470 8390 8490 8440
rect 8410 8370 8490 8390
rect 8810 8580 8890 8600
rect 8810 8530 8830 8580
rect 8870 8530 8890 8580
rect 8810 8440 8890 8530
rect 8810 8390 8830 8440
rect 8870 8390 8890 8440
rect 8810 8370 8890 8390
rect 9210 8580 9290 8600
rect 9210 8530 9230 8580
rect 9270 8530 9290 8580
rect 9210 8440 9290 8530
rect 9210 8390 9230 8440
rect 9270 8390 9290 8440
rect 9210 8370 9290 8390
rect 9610 8580 9690 8600
rect 9610 8530 9630 8580
rect 9670 8530 9690 8580
rect 9610 8440 9690 8530
rect 9610 8390 9630 8440
rect 9670 8390 9690 8440
rect 9610 8370 9690 8390
rect 10010 8580 10090 8600
rect 10010 8530 10030 8580
rect 10070 8530 10090 8580
rect 10010 8440 10090 8530
rect 10010 8390 10030 8440
rect 10070 8390 10090 8440
rect 10010 8370 10090 8390
rect 8210 8310 8290 8330
rect 8210 8270 8230 8310
rect 8270 8270 8290 8310
rect 8210 8250 8290 8270
rect 6570 8150 6580 8210
rect 6640 8150 6660 8210
rect 6720 8150 6740 8210
rect 6800 8150 6810 8210
rect 8230 8180 8270 8250
rect 8430 8180 8470 8370
rect 8830 8180 8870 8370
rect 9230 8180 9270 8370
rect 9630 8180 9670 8370
rect 9790 8280 9870 8290
rect 9790 8220 9800 8280
rect 9860 8220 9870 8280
rect 9790 8210 9870 8220
rect 10030 8180 10070 8370
rect 10210 8310 10290 8330
rect 10210 8270 10230 8310
rect 10270 8270 10290 8310
rect 10210 8250 10290 8270
rect 10230 8180 10270 8250
rect 6570 8130 6810 8150
rect 6570 8070 6580 8130
rect 6640 8070 6660 8130
rect 6720 8070 6740 8130
rect 6800 8070 6810 8130
rect 7830 8160 10990 8180
rect 7830 8100 7850 8160
rect 7910 8120 7990 8160
rect 8030 8120 8090 8160
rect 8130 8120 8190 8160
rect 8230 8120 8290 8160
rect 8330 8120 8390 8160
rect 8430 8120 8490 8160
rect 8530 8120 8590 8160
rect 8630 8120 8690 8160
rect 8730 8120 8790 8160
rect 8830 8120 8890 8160
rect 8930 8120 8990 8160
rect 9030 8120 9090 8160
rect 9130 8120 9190 8160
rect 9230 8120 9290 8160
rect 9330 8120 9390 8160
rect 9430 8120 9490 8160
rect 9530 8120 9590 8160
rect 9630 8120 9690 8160
rect 9730 8120 9790 8160
rect 9830 8120 9890 8160
rect 9930 8120 9990 8160
rect 10030 8120 10090 8160
rect 10130 8120 10190 8160
rect 10230 8120 10290 8160
rect 10330 8120 10390 8160
rect 10430 8120 10490 8160
rect 10530 8120 10590 8160
rect 10630 8120 10690 8160
rect 10730 8120 10790 8160
rect 10830 8120 10890 8160
rect 10930 8120 10990 8160
rect 7910 8100 10990 8120
rect 7830 8080 7930 8100
rect 6570 8050 6810 8070
rect 6570 7990 6580 8050
rect 6640 7990 6660 8050
rect 6720 7990 6740 8050
rect 6800 7990 6810 8050
rect 9790 8060 9870 8070
rect 9790 8000 9800 8060
rect 9860 8000 9870 8060
rect 9790 7990 9870 8000
rect 6570 7980 6810 7990
rect 11750 7880 11860 7900
rect 11750 7810 11770 7880
rect 11840 7810 11860 7880
rect 11750 7790 11860 7810
rect 9570 7780 9650 7790
rect 8890 7720 8970 7730
rect 7550 7710 7630 7720
rect 7550 7650 7560 7710
rect 7620 7650 7630 7710
rect 7550 7640 7630 7650
rect 8070 7700 8150 7710
rect 8070 7640 8080 7700
rect 8140 7680 8150 7700
rect 8890 7680 8900 7720
rect 8140 7660 8900 7680
rect 8960 7680 8970 7720
rect 9570 7720 9580 7780
rect 9640 7720 9650 7780
rect 9570 7710 9650 7720
rect 10010 7750 10090 7770
rect 10010 7710 10030 7750
rect 10070 7710 10090 7750
rect 10010 7680 10090 7710
rect 8960 7660 10090 7680
rect 8140 7650 10090 7660
rect 10710 7650 10790 7670
rect 8140 7640 8150 7650
rect 6460 7530 6470 7590
rect 6530 7530 6540 7590
rect 6460 7520 6540 7530
rect 7440 7540 7520 7550
rect 7440 7480 7450 7540
rect 7510 7480 7520 7540
rect 7440 7470 7520 7480
rect 6230 6990 6310 7000
rect 6230 6930 6240 6990
rect 6300 6930 6310 6990
rect 6230 6920 6310 6930
rect 6140 6880 6220 6890
rect 6140 6820 6150 6880
rect 6210 6820 6220 6880
rect 6140 6810 6220 6820
rect 5700 6520 5720 6560
rect 5760 6520 5780 6560
rect 5700 6500 5780 6520
rect 5820 6570 5900 6580
rect 5820 6510 5830 6570
rect 5890 6510 5900 6570
rect 5820 6500 5900 6510
rect 5490 6440 5550 6460
rect 5490 6400 5500 6440
rect 5540 6400 5550 6440
rect 5490 6340 5550 6400
rect 5490 6300 5500 6340
rect 5540 6300 5550 6340
rect 5490 6240 5550 6300
rect 5600 6440 5660 6500
rect 5600 6400 5610 6440
rect 5650 6400 5660 6440
rect 5600 6340 5660 6400
rect 5600 6300 5610 6340
rect 5650 6300 5660 6340
rect 5600 6280 5660 6300
rect 5710 6440 5770 6460
rect 5710 6400 5720 6440
rect 5760 6400 5770 6440
rect 5710 6340 5770 6400
rect 5710 6300 5720 6340
rect 5760 6300 5770 6340
rect 5710 6240 5770 6300
rect 5820 6440 5880 6500
rect 5820 6400 5830 6440
rect 5870 6400 5880 6440
rect 5820 6340 5880 6400
rect 5820 6300 5830 6340
rect 5870 6300 5880 6340
rect 5820 6280 5880 6300
rect 5930 6440 5990 6460
rect 5930 6400 5940 6440
rect 5980 6400 5990 6440
rect 5930 6340 5990 6400
rect 5930 6300 5940 6340
rect 5980 6300 5990 6340
rect 5930 6240 5990 6300
rect 4860 6200 4870 6240
rect 4910 6200 4920 6240
rect 4860 6140 4920 6200
rect 5230 6230 5310 6240
rect 5230 6170 5240 6230
rect 5300 6170 5310 6230
rect 5230 6160 5310 6170
rect 5480 6220 5560 6240
rect 5480 6180 5500 6220
rect 5540 6180 5560 6220
rect 5480 6160 5560 6180
rect 5700 6230 5780 6240
rect 5700 6170 5710 6230
rect 5770 6170 5780 6230
rect 5700 6160 5780 6170
rect 5920 6220 6000 6240
rect 5920 6180 5940 6220
rect 5980 6180 6000 6220
rect 5920 6160 6000 6180
rect 4860 6100 4870 6140
rect 4910 6100 4920 6140
rect 4860 6080 4920 6100
rect 5490 6040 5550 6160
rect 5930 6040 5990 6160
rect 1610 6030 1690 6040
rect 1610 5970 1620 6030
rect 1680 5970 1690 6030
rect 1610 5950 1690 5970
rect 1610 5890 1620 5950
rect 1680 5890 1690 5950
rect 1610 5870 1690 5890
rect 1610 5810 1620 5870
rect 1680 5810 1690 5870
rect 1610 5800 1690 5810
rect 1970 6030 2050 6040
rect 1970 5970 1980 6030
rect 2040 5970 2050 6030
rect 1970 5950 2050 5970
rect 1970 5890 1980 5950
rect 2040 5890 2050 5950
rect 1970 5870 2050 5890
rect 1970 5810 1980 5870
rect 2040 5810 2050 5870
rect 1970 5800 2050 5810
rect 2330 6030 2410 6040
rect 2330 5970 2340 6030
rect 2400 5970 2410 6030
rect 2330 5950 2410 5970
rect 2330 5890 2340 5950
rect 2400 5890 2410 5950
rect 2330 5870 2410 5890
rect 2330 5810 2340 5870
rect 2400 5810 2410 5870
rect 2330 5800 2410 5810
rect 2690 6030 2770 6040
rect 2690 5970 2700 6030
rect 2760 5970 2770 6030
rect 2690 5950 2770 5970
rect 2690 5890 2700 5950
rect 2760 5890 2770 5950
rect 2690 5870 2770 5890
rect 2690 5810 2700 5870
rect 2760 5810 2770 5870
rect 2690 5800 2770 5810
rect 3050 6030 3130 6040
rect 3050 5970 3060 6030
rect 3120 5970 3130 6030
rect 3050 5950 3130 5970
rect 3050 5890 3060 5950
rect 3120 5890 3130 5950
rect 3050 5870 3130 5890
rect 3050 5810 3060 5870
rect 3120 5810 3130 5870
rect 3050 5800 3130 5810
rect 3410 6030 3490 6040
rect 3410 5970 3420 6030
rect 3480 5970 3490 6030
rect 3410 5950 3490 5970
rect 3410 5890 3420 5950
rect 3480 5890 3490 5950
rect 3410 5870 3490 5890
rect 3410 5810 3420 5870
rect 3480 5810 3490 5870
rect 3410 5800 3490 5810
rect 3770 6030 3850 6040
rect 3770 5970 3780 6030
rect 3840 5970 3850 6030
rect 3770 5950 3850 5970
rect 3770 5890 3780 5950
rect 3840 5890 3850 5950
rect 3770 5870 3850 5890
rect 3770 5810 3780 5870
rect 3840 5810 3850 5870
rect 3770 5800 3850 5810
rect 4130 6030 4210 6040
rect 4130 5970 4140 6030
rect 4200 5970 4210 6030
rect 4130 5950 4210 5970
rect 4130 5890 4140 5950
rect 4200 5890 4210 5950
rect 4130 5870 4210 5890
rect 4130 5810 4140 5870
rect 4200 5810 4210 5870
rect 4130 5800 4210 5810
rect 4490 6030 4570 6040
rect 4490 5970 4500 6030
rect 4560 5970 4570 6030
rect 4490 5950 4570 5970
rect 4490 5890 4500 5950
rect 4560 5890 4570 5950
rect 4490 5870 4570 5890
rect 4490 5810 4500 5870
rect 4560 5810 4570 5870
rect 4490 5800 4570 5810
rect 4850 6030 4930 6040
rect 4850 5970 4860 6030
rect 4920 5970 4930 6030
rect 4850 5950 4930 5970
rect 4850 5890 4860 5950
rect 4920 5890 4930 5950
rect 4850 5870 4930 5890
rect 4850 5810 4860 5870
rect 4920 5810 4930 5870
rect 4850 5800 4930 5810
rect 5480 6030 5560 6040
rect 5480 5970 5490 6030
rect 5550 5970 5560 6030
rect 5480 5950 5560 5970
rect 5480 5890 5490 5950
rect 5550 5890 5560 5950
rect 5480 5870 5560 5890
rect 5480 5810 5490 5870
rect 5550 5810 5560 5870
rect 5480 5800 5560 5810
rect 5920 6030 6000 6040
rect 5920 5970 5930 6030
rect 5990 5970 6000 6030
rect 5920 5950 6000 5970
rect 5920 5890 5930 5950
rect 5990 5890 6000 5950
rect 5920 5870 6000 5890
rect 5920 5810 5930 5870
rect 5990 5810 6000 5870
rect 5920 5800 6000 5810
rect 1796 5760 1854 5770
rect 1796 5708 1798 5760
rect 1850 5708 1854 5760
rect 1796 5700 1854 5708
rect 1906 5760 1964 5770
rect 1906 5708 1908 5760
rect 1960 5708 1964 5760
rect 1906 5700 1964 5708
rect 2016 5760 2074 5770
rect 2016 5708 2018 5760
rect 2070 5708 2074 5760
rect 2016 5700 2074 5708
rect 2126 5760 2184 5770
rect 2126 5708 2128 5760
rect 2180 5708 2184 5760
rect 2126 5700 2184 5708
rect 2236 5760 2294 5770
rect 2236 5708 2238 5760
rect 2290 5708 2294 5760
rect 2236 5700 2294 5708
rect 2346 5760 2404 5770
rect 2346 5708 2348 5760
rect 2400 5708 2404 5760
rect 2346 5700 2404 5708
rect 2456 5760 2514 5770
rect 2456 5708 2458 5760
rect 2510 5708 2514 5760
rect 2456 5700 2514 5708
rect 2566 5760 2624 5770
rect 2566 5708 2568 5760
rect 2620 5708 2624 5760
rect 2566 5700 2624 5708
rect 2676 5760 2734 5770
rect 2676 5708 2678 5760
rect 2730 5708 2734 5760
rect 2676 5700 2734 5708
rect 2786 5760 2844 5770
rect 2786 5708 2788 5760
rect 2840 5708 2844 5760
rect 2786 5700 2844 5708
rect 3696 5760 3754 5770
rect 3696 5708 3698 5760
rect 3750 5708 3754 5760
rect 3696 5700 3754 5708
rect 3806 5760 3864 5770
rect 3806 5708 3808 5760
rect 3860 5708 3864 5760
rect 3806 5700 3864 5708
rect 3916 5760 3974 5770
rect 3916 5708 3918 5760
rect 3970 5708 3974 5760
rect 3916 5700 3974 5708
rect 4026 5760 4084 5770
rect 4026 5708 4028 5760
rect 4080 5708 4084 5760
rect 4026 5700 4084 5708
rect 4136 5760 4194 5770
rect 4136 5708 4138 5760
rect 4190 5708 4194 5760
rect 4136 5700 4194 5708
rect 4246 5760 4304 5770
rect 4246 5708 4248 5760
rect 4300 5708 4304 5760
rect 4246 5700 4304 5708
rect 4356 5760 4414 5770
rect 4356 5708 4358 5760
rect 4410 5708 4414 5760
rect 4356 5700 4414 5708
rect 4466 5760 4524 5770
rect 4466 5708 4468 5760
rect 4520 5708 4524 5760
rect 4466 5700 4524 5708
rect 4576 5760 4634 5770
rect 4576 5708 4578 5760
rect 4630 5708 4634 5760
rect 4576 5700 4634 5708
rect 4686 5760 4744 5770
rect 4686 5708 4688 5760
rect 4740 5708 4744 5760
rect 4686 5700 4744 5708
rect 1550 5640 1690 5660
rect 1550 5600 1560 5640
rect 1600 5600 1640 5640
rect 1680 5600 1690 5640
rect 1550 5540 1690 5600
rect 1550 5500 1560 5540
rect 1600 5500 1640 5540
rect 1680 5500 1690 5540
rect 1550 5480 1690 5500
rect 1630 5440 1690 5480
rect 1740 5640 1800 5660
rect 1740 5600 1750 5640
rect 1790 5600 1800 5640
rect 1740 5540 1800 5600
rect 1740 5500 1750 5540
rect 1790 5500 1800 5540
rect 1620 5430 1700 5440
rect 1620 5370 1630 5430
rect 1690 5370 1700 5430
rect 1620 5360 1700 5370
rect 1740 5330 1800 5500
rect 1850 5640 1910 5660
rect 1850 5600 1860 5640
rect 1900 5600 1910 5640
rect 1850 5540 1910 5600
rect 1850 5500 1860 5540
rect 1900 5500 1910 5540
rect 1850 5440 1910 5500
rect 1960 5640 2020 5660
rect 1960 5600 1970 5640
rect 2010 5600 2020 5640
rect 1960 5540 2020 5600
rect 1960 5500 1970 5540
rect 2010 5500 2020 5540
rect 1840 5430 1920 5440
rect 1840 5370 1850 5430
rect 1910 5370 1920 5430
rect 1840 5360 1920 5370
rect 1960 5330 2020 5500
rect 2070 5640 2130 5660
rect 2070 5600 2080 5640
rect 2120 5600 2130 5640
rect 2070 5540 2130 5600
rect 2070 5500 2080 5540
rect 2120 5500 2130 5540
rect 2070 5440 2130 5500
rect 2180 5640 2240 5660
rect 2180 5600 2190 5640
rect 2230 5600 2240 5640
rect 2180 5540 2240 5600
rect 2180 5500 2190 5540
rect 2230 5500 2240 5540
rect 2060 5430 2140 5440
rect 2060 5370 2070 5430
rect 2130 5370 2140 5430
rect 2060 5360 2140 5370
rect 2180 5330 2240 5500
rect 2290 5640 2350 5660
rect 2290 5600 2300 5640
rect 2340 5600 2350 5640
rect 2290 5540 2350 5600
rect 2290 5500 2300 5540
rect 2340 5500 2350 5540
rect 2290 5440 2350 5500
rect 2400 5640 2460 5660
rect 2400 5600 2410 5640
rect 2450 5600 2460 5640
rect 2400 5540 2460 5600
rect 2400 5500 2410 5540
rect 2450 5500 2460 5540
rect 2280 5430 2360 5440
rect 2280 5370 2290 5430
rect 2350 5370 2360 5430
rect 2280 5360 2360 5370
rect 2400 5330 2460 5500
rect 2510 5640 2570 5660
rect 2510 5600 2520 5640
rect 2560 5600 2570 5640
rect 2510 5540 2570 5600
rect 2510 5500 2520 5540
rect 2560 5500 2570 5540
rect 2510 5440 2570 5500
rect 2620 5640 2680 5660
rect 2620 5600 2630 5640
rect 2670 5600 2680 5640
rect 2620 5540 2680 5600
rect 2620 5500 2630 5540
rect 2670 5500 2680 5540
rect 2500 5430 2580 5440
rect 2500 5370 2510 5430
rect 2570 5370 2580 5430
rect 2500 5360 2580 5370
rect 2620 5330 2680 5500
rect 2730 5640 2790 5660
rect 2730 5600 2740 5640
rect 2780 5600 2790 5640
rect 2730 5540 2790 5600
rect 2730 5500 2740 5540
rect 2780 5500 2790 5540
rect 2730 5440 2790 5500
rect 2840 5640 2900 5660
rect 2840 5600 2850 5640
rect 2890 5600 2900 5640
rect 2840 5540 2900 5600
rect 2840 5500 2850 5540
rect 2890 5500 2900 5540
rect 2720 5430 2800 5440
rect 2720 5370 2730 5430
rect 2790 5370 2800 5430
rect 2720 5360 2800 5370
rect 2840 5330 2900 5500
rect 2950 5640 3090 5660
rect 2950 5600 2960 5640
rect 3000 5600 3040 5640
rect 3080 5600 3090 5640
rect 2950 5540 3090 5600
rect 2950 5500 2960 5540
rect 3000 5500 3040 5540
rect 3080 5500 3090 5540
rect 2950 5480 3090 5500
rect 3450 5640 3590 5660
rect 3450 5600 3460 5640
rect 3500 5600 3540 5640
rect 3580 5600 3590 5640
rect 3450 5540 3590 5600
rect 3450 5500 3460 5540
rect 3500 5500 3540 5540
rect 3580 5500 3590 5540
rect 3450 5480 3590 5500
rect 2950 5440 3010 5480
rect 3530 5440 3590 5480
rect 3640 5640 3700 5660
rect 3640 5600 3650 5640
rect 3690 5600 3700 5640
rect 3640 5540 3700 5600
rect 3640 5500 3650 5540
rect 3690 5500 3700 5540
rect 2940 5430 3020 5440
rect 2940 5370 2950 5430
rect 3010 5370 3020 5430
rect 2940 5360 3020 5370
rect 3520 5430 3600 5440
rect 3520 5370 3530 5430
rect 3590 5370 3600 5430
rect 3520 5360 3600 5370
rect 3640 5330 3700 5500
rect 3750 5640 3810 5660
rect 3750 5600 3760 5640
rect 3800 5600 3810 5640
rect 3750 5540 3810 5600
rect 3750 5500 3760 5540
rect 3800 5500 3810 5540
rect 3750 5440 3810 5500
rect 3860 5640 3920 5660
rect 3860 5600 3870 5640
rect 3910 5600 3920 5640
rect 3860 5540 3920 5600
rect 3860 5500 3870 5540
rect 3910 5500 3920 5540
rect 3740 5430 3820 5440
rect 3740 5370 3750 5430
rect 3810 5370 3820 5430
rect 3740 5360 3820 5370
rect 3860 5330 3920 5500
rect 3970 5640 4030 5660
rect 3970 5600 3980 5640
rect 4020 5600 4030 5640
rect 3970 5540 4030 5600
rect 3970 5500 3980 5540
rect 4020 5500 4030 5540
rect 3970 5440 4030 5500
rect 4080 5640 4140 5660
rect 4080 5600 4090 5640
rect 4130 5600 4140 5640
rect 4080 5540 4140 5600
rect 4080 5500 4090 5540
rect 4130 5500 4140 5540
rect 3960 5430 4040 5440
rect 3960 5370 3970 5430
rect 4030 5370 4040 5430
rect 3960 5360 4040 5370
rect 4080 5330 4140 5500
rect 4190 5640 4250 5660
rect 4190 5600 4200 5640
rect 4240 5600 4250 5640
rect 4190 5540 4250 5600
rect 4190 5500 4200 5540
rect 4240 5500 4250 5540
rect 4190 5440 4250 5500
rect 4300 5640 4360 5660
rect 4300 5600 4310 5640
rect 4350 5600 4360 5640
rect 4300 5540 4360 5600
rect 4300 5500 4310 5540
rect 4350 5500 4360 5540
rect 4180 5430 4260 5440
rect 4180 5370 4190 5430
rect 4250 5370 4260 5430
rect 4180 5360 4260 5370
rect 4300 5330 4360 5500
rect 4410 5640 4470 5660
rect 4410 5600 4420 5640
rect 4460 5600 4470 5640
rect 4410 5540 4470 5600
rect 4410 5500 4420 5540
rect 4460 5500 4470 5540
rect 4410 5440 4470 5500
rect 4520 5640 4580 5660
rect 4520 5600 4530 5640
rect 4570 5600 4580 5640
rect 4520 5540 4580 5600
rect 4520 5500 4530 5540
rect 4570 5500 4580 5540
rect 4400 5430 4480 5440
rect 4400 5370 4410 5430
rect 4470 5370 4480 5430
rect 4400 5360 4480 5370
rect 4520 5330 4580 5500
rect 4630 5640 4690 5660
rect 4630 5600 4640 5640
rect 4680 5600 4690 5640
rect 4630 5540 4690 5600
rect 4630 5500 4640 5540
rect 4680 5500 4690 5540
rect 4630 5440 4690 5500
rect 4740 5640 4800 5660
rect 4740 5600 4750 5640
rect 4790 5600 4800 5640
rect 4740 5540 4800 5600
rect 4740 5500 4750 5540
rect 4790 5500 4800 5540
rect 4620 5430 4700 5440
rect 4620 5370 4630 5430
rect 4690 5370 4700 5430
rect 4620 5360 4700 5370
rect 4740 5330 4800 5500
rect 4850 5640 4990 5660
rect 4850 5600 4860 5640
rect 4900 5600 4940 5640
rect 4980 5600 4990 5640
rect 4850 5540 4990 5600
rect 4850 5500 4860 5540
rect 4900 5500 4940 5540
rect 4980 5500 4990 5540
rect 4850 5480 4990 5500
rect 4850 5440 4910 5480
rect 4840 5430 4920 5440
rect 4840 5370 4850 5430
rect 4910 5370 4920 5430
rect 4840 5360 4920 5370
rect 340 5260 350 5320
rect 410 5260 420 5320
rect 340 5250 420 5260
rect 1730 5320 1810 5330
rect 1730 5260 1740 5320
rect 1800 5260 1810 5320
rect 1730 5250 1810 5260
rect 1950 5320 2030 5330
rect 1950 5260 1960 5320
rect 2020 5260 2030 5320
rect 1950 5250 2030 5260
rect 2170 5320 2250 5330
rect 2170 5260 2180 5320
rect 2240 5260 2250 5320
rect 2170 5250 2250 5260
rect 2390 5320 2470 5330
rect 2390 5260 2400 5320
rect 2460 5260 2470 5320
rect 2390 5250 2470 5260
rect 2610 5320 2690 5330
rect 2610 5260 2620 5320
rect 2680 5260 2690 5320
rect 2610 5250 2690 5260
rect 2830 5320 2910 5330
rect 2830 5260 2840 5320
rect 2900 5260 2910 5320
rect 2830 5250 2910 5260
rect 3630 5320 3710 5330
rect 3630 5260 3640 5320
rect 3700 5260 3710 5320
rect 1150 5210 1390 5220
rect 1150 5150 1160 5210
rect 1220 5150 1240 5210
rect 1300 5150 1320 5210
rect 1380 5150 1390 5210
rect 1150 5130 1390 5150
rect 1150 5070 1160 5130
rect 1220 5070 1240 5130
rect 1300 5070 1320 5130
rect 1380 5070 1390 5130
rect 1150 5050 1390 5070
rect 1150 4990 1160 5050
rect 1220 4990 1240 5050
rect 1300 4990 1320 5050
rect 1380 4990 1390 5050
rect 1150 2460 1390 4990
rect 3630 5210 3710 5260
rect 3630 5150 3640 5210
rect 3700 5150 3710 5210
rect 3630 5130 3710 5150
rect 3630 5070 3640 5130
rect 3700 5070 3710 5130
rect 3630 5050 3710 5070
rect 3630 4990 3640 5050
rect 3700 4990 3710 5050
rect 3630 4980 3710 4990
rect 3850 5320 3930 5330
rect 3850 5260 3860 5320
rect 3920 5260 3930 5320
rect 3850 5210 3930 5260
rect 3850 5150 3860 5210
rect 3920 5150 3930 5210
rect 3850 5130 3930 5150
rect 3850 5070 3860 5130
rect 3920 5070 3930 5130
rect 3850 5050 3930 5070
rect 3850 4990 3860 5050
rect 3920 4990 3930 5050
rect 3850 4980 3930 4990
rect 4070 5320 4150 5330
rect 4070 5260 4080 5320
rect 4140 5260 4150 5320
rect 4070 5210 4150 5260
rect 4070 5150 4080 5210
rect 4140 5150 4150 5210
rect 4070 5130 4150 5150
rect 4070 5070 4080 5130
rect 4140 5070 4150 5130
rect 4070 5050 4150 5070
rect 4070 4990 4080 5050
rect 4140 4990 4150 5050
rect 4070 4980 4150 4990
rect 4290 5320 4370 5330
rect 4290 5260 4300 5320
rect 4360 5260 4370 5320
rect 4290 5210 4370 5260
rect 4290 5150 4300 5210
rect 4360 5150 4370 5210
rect 4290 5130 4370 5150
rect 4290 5070 4300 5130
rect 4360 5070 4370 5130
rect 4290 5050 4370 5070
rect 4290 4990 4300 5050
rect 4360 4990 4370 5050
rect 4290 4980 4370 4990
rect 4510 5320 4590 5330
rect 4510 5260 4520 5320
rect 4580 5260 4590 5320
rect 4510 5210 4590 5260
rect 4510 5150 4520 5210
rect 4580 5150 4590 5210
rect 4510 5130 4590 5150
rect 4510 5070 4520 5130
rect 4580 5070 4590 5130
rect 4510 5050 4590 5070
rect 4510 4990 4520 5050
rect 4580 4990 4590 5050
rect 4510 4980 4590 4990
rect 4730 5320 4810 5330
rect 4730 5260 4740 5320
rect 4800 5260 4810 5320
rect 4730 5210 4810 5260
rect 4730 5150 4740 5210
rect 4800 5150 4810 5210
rect 7460 5200 7500 7470
rect 4730 5130 4810 5150
rect 4730 5070 4740 5130
rect 4800 5070 4810 5130
rect 7440 5190 7520 5200
rect 7440 5130 7450 5190
rect 7510 5130 7520 5190
rect 7440 5120 7520 5130
rect 4730 5050 4810 5070
rect 4730 4990 4740 5050
rect 4800 4990 4810 5050
rect 7350 5080 7430 5090
rect 7350 5020 7360 5080
rect 7420 5020 7430 5080
rect 7350 5010 7430 5020
rect 4730 4980 4810 4990
rect 7040 4950 7140 4960
rect 1720 4940 7140 4950
rect 1720 4930 7060 4940
rect 1720 4870 1740 4930
rect 1800 4890 1880 4930
rect 1920 4890 1980 4930
rect 2020 4890 2080 4930
rect 2120 4890 2180 4930
rect 2220 4890 2280 4930
rect 2320 4890 2380 4930
rect 2420 4890 2480 4930
rect 2520 4890 2580 4930
rect 2620 4890 2680 4930
rect 2720 4890 2780 4930
rect 2820 4890 2880 4930
rect 2920 4890 2980 4930
rect 3020 4890 3080 4930
rect 3120 4890 3180 4930
rect 3220 4890 3280 4930
rect 3320 4890 3380 4930
rect 3420 4890 3480 4930
rect 3520 4890 3580 4930
rect 3620 4890 3680 4930
rect 3720 4890 3780 4930
rect 3820 4890 3880 4930
rect 3920 4890 3980 4930
rect 4020 4890 4080 4930
rect 4120 4890 4180 4930
rect 4220 4890 4280 4930
rect 4320 4890 4380 4930
rect 4420 4890 4480 4930
rect 4520 4890 4580 4930
rect 4620 4890 4680 4930
rect 4720 4890 4780 4930
rect 4820 4890 4880 4930
rect 4920 4890 4980 4930
rect 5020 4890 5080 4930
rect 5120 4890 5180 4930
rect 5220 4890 5280 4930
rect 5320 4890 5380 4930
rect 5420 4890 5480 4930
rect 5520 4890 5580 4930
rect 5620 4890 5680 4930
rect 5720 4890 5780 4930
rect 5820 4890 5880 4930
rect 5920 4890 5980 4930
rect 6020 4890 6080 4930
rect 6120 4890 6180 4930
rect 6220 4890 6280 4930
rect 6320 4890 6380 4930
rect 6420 4890 6480 4930
rect 6520 4890 6580 4930
rect 6620 4890 6680 4930
rect 6720 4890 6780 4930
rect 6820 4890 6880 4930
rect 6920 4890 7060 4930
rect 1800 4880 7060 4890
rect 7120 4880 7140 4940
rect 1800 4870 7140 4880
rect 1720 4850 1820 4870
rect 7040 4860 7140 4870
rect 2550 4820 2630 4840
rect 2550 4780 2570 4820
rect 2610 4800 2630 4820
rect 4270 4820 4350 4840
rect 4270 4800 4290 4820
rect 2610 4780 4290 4800
rect 4330 4800 4350 4820
rect 6340 4830 6420 4840
rect 4330 4780 5180 4800
rect 2550 4760 5180 4780
rect 6340 4770 6350 4830
rect 6410 4770 6420 4830
rect 6340 4760 6420 4770
rect 1930 4480 2010 4490
rect 1930 4420 1940 4480
rect 2000 4420 2010 4480
rect 1930 4410 2010 4420
rect 3840 4480 3920 4490
rect 3840 4420 3850 4480
rect 3910 4420 3920 4480
rect 5140 4480 5180 4760
rect 7370 4710 7410 5010
rect 7440 4830 7520 4840
rect 7440 4770 7450 4830
rect 7510 4770 7520 4830
rect 7440 4760 7520 4770
rect 6640 4700 6720 4710
rect 6640 4640 6650 4700
rect 6710 4640 6720 4700
rect 6640 4630 6720 4640
rect 7350 4700 7430 4710
rect 7350 4640 7360 4700
rect 7420 4640 7430 4700
rect 7350 4630 7430 4640
rect 5140 4460 5220 4480
rect 3840 4410 3920 4420
rect 5010 4440 5090 4450
rect 5010 4380 5020 4440
rect 5080 4380 5090 4440
rect 5140 4420 5160 4460
rect 5200 4420 5220 4460
rect 6660 4420 6700 4630
rect 5140 4400 5220 4420
rect 6640 4410 6720 4420
rect 5010 4370 5090 4380
rect 6640 4350 6650 4410
rect 6710 4350 6720 4410
rect 6640 4340 6720 4350
rect 6880 4410 6960 4420
rect 6880 4350 6890 4410
rect 6950 4350 6960 4410
rect 6880 4340 6960 4350
rect 7350 4410 7430 4420
rect 7350 4350 7360 4410
rect 7420 4350 7430 4410
rect 7350 4340 7430 4350
rect 4140 3870 4220 3880
rect 4140 3810 4150 3870
rect 4210 3810 4220 3870
rect 4140 3800 4220 3810
rect 1900 3770 2000 3780
rect 7200 3770 7300 3790
rect 1900 3760 7220 3770
rect 1900 3700 1920 3760
rect 1980 3750 7220 3760
rect 1980 3710 2080 3750
rect 2120 3710 2180 3750
rect 2220 3710 2280 3750
rect 2320 3710 2380 3750
rect 2420 3710 2480 3750
rect 2520 3710 2580 3750
rect 2620 3710 2680 3750
rect 2720 3710 2780 3750
rect 2820 3710 2880 3750
rect 2920 3710 2980 3750
rect 3020 3710 3080 3750
rect 3120 3710 3180 3750
rect 3220 3710 3280 3750
rect 3320 3710 3380 3750
rect 3420 3710 3480 3750
rect 3520 3710 3580 3750
rect 3620 3710 3680 3750
rect 3720 3710 3780 3750
rect 3820 3710 3880 3750
rect 3920 3710 3980 3750
rect 4020 3710 4080 3750
rect 4120 3710 4180 3750
rect 4220 3710 4280 3750
rect 4320 3710 4380 3750
rect 4420 3710 4480 3750
rect 4520 3710 4580 3750
rect 4620 3710 4680 3750
rect 4720 3710 4780 3750
rect 4820 3710 4880 3750
rect 4920 3710 4980 3750
rect 5020 3710 5080 3750
rect 5120 3710 5180 3750
rect 5220 3710 5280 3750
rect 5320 3710 5380 3750
rect 5420 3710 5480 3750
rect 5520 3710 5580 3750
rect 5620 3710 5680 3750
rect 5720 3710 5780 3750
rect 5820 3710 5880 3750
rect 5920 3710 5980 3750
rect 6020 3710 6080 3750
rect 6120 3710 6180 3750
rect 6220 3710 6280 3750
rect 6320 3710 6380 3750
rect 6420 3710 6480 3750
rect 6520 3710 6580 3750
rect 6620 3710 6680 3750
rect 6720 3710 6780 3750
rect 6820 3710 6880 3750
rect 6920 3710 6980 3750
rect 7020 3710 7080 3750
rect 7120 3710 7220 3750
rect 7280 3710 7300 3770
rect 7370 3740 7410 4340
rect 7460 3900 7500 4760
rect 7440 3890 7520 3900
rect 7440 3830 7450 3890
rect 7510 3830 7520 3890
rect 7440 3820 7520 3830
rect 7570 3810 7610 7640
rect 8070 7630 8150 7640
rect 10710 7620 10730 7650
rect 9330 7610 10730 7620
rect 10770 7610 10790 7650
rect 9330 7600 10790 7610
rect 8430 7560 8510 7570
rect 8070 7540 8150 7550
rect 8070 7480 8080 7540
rect 8140 7520 8150 7540
rect 8430 7520 8440 7560
rect 8140 7500 8440 7520
rect 8500 7520 8510 7560
rect 9330 7560 9350 7600
rect 9390 7590 10790 7600
rect 11920 7600 12000 7620
rect 14230 7610 14310 7620
rect 14230 7600 14240 7610
rect 9390 7560 9410 7590
rect 11920 7560 11940 7600
rect 11980 7570 14240 7600
rect 11980 7560 12000 7570
rect 9330 7550 9410 7560
rect 9570 7550 9650 7560
rect 9570 7520 9580 7550
rect 8500 7500 9580 7520
rect 8140 7490 9580 7500
rect 9640 7490 9650 7550
rect 11920 7540 12000 7560
rect 14230 7550 14240 7570
rect 14300 7550 14310 7610
rect 14230 7540 14310 7550
rect 8140 7480 8150 7490
rect 9570 7480 9650 7490
rect 8070 7470 8150 7480
rect 8430 7450 8510 7460
rect 8430 7390 8440 7450
rect 8500 7390 8510 7450
rect 8430 7380 8510 7390
rect 8870 7450 8950 7460
rect 8870 7390 8880 7450
rect 8940 7390 8950 7450
rect 8870 7380 8950 7390
rect 11750 7380 11860 7400
rect 11750 7310 11770 7380
rect 11840 7310 11860 7380
rect 11750 7290 11860 7310
rect 8750 7070 8830 7080
rect 8750 7010 8760 7070
rect 8820 7010 8830 7070
rect 8750 7000 8830 7010
rect 7830 6970 7930 6990
rect 7830 6910 7850 6970
rect 7910 6950 10990 6970
rect 7910 6910 7990 6950
rect 8030 6910 8090 6950
rect 8130 6910 8190 6950
rect 8230 6910 8290 6950
rect 8330 6910 8390 6950
rect 8430 6910 8490 6950
rect 8530 6910 8590 6950
rect 8630 6910 8690 6950
rect 8730 6910 8790 6950
rect 8830 6910 8890 6950
rect 8930 6910 8990 6950
rect 9030 6910 9090 6950
rect 9130 6910 9190 6950
rect 9230 6910 9290 6950
rect 9330 6910 9390 6950
rect 9430 6910 9490 6950
rect 9530 6910 9590 6950
rect 9630 6910 9690 6950
rect 9730 6910 9790 6950
rect 9830 6910 9890 6950
rect 9930 6910 9990 6950
rect 10030 6910 10090 6950
rect 10130 6910 10190 6950
rect 10230 6910 10290 6950
rect 10330 6910 10390 6950
rect 10430 6910 10490 6950
rect 10530 6910 10590 6950
rect 10630 6910 10690 6950
rect 10730 6910 10790 6950
rect 10830 6910 10890 6950
rect 10930 6910 10990 6950
rect 7830 6890 10990 6910
rect 8350 6810 8390 6890
rect 8330 6790 8410 6810
rect 8330 6750 8350 6790
rect 8390 6750 8410 6790
rect 8330 6730 8410 6750
rect 8550 6690 8590 6890
rect 8750 6850 8830 6860
rect 8750 6790 8760 6850
rect 8820 6790 8830 6850
rect 8750 6780 8830 6790
rect 8950 6690 8990 6890
rect 9350 6690 9390 6890
rect 9750 6690 9790 6890
rect 10150 6690 10190 6890
rect 10350 6810 10390 6890
rect 10330 6730 10410 6810
rect 8530 6670 8610 6690
rect 8530 6630 8550 6670
rect 8590 6630 8610 6670
rect 8530 6570 8610 6630
rect 8530 6530 8550 6570
rect 8590 6530 8610 6570
rect 8530 6470 8610 6530
rect 8530 6430 8550 6470
rect 8590 6430 8610 6470
rect 8530 6370 8610 6430
rect 8530 6330 8550 6370
rect 8590 6330 8610 6370
rect 8530 6270 8610 6330
rect 8530 6230 8550 6270
rect 8590 6230 8610 6270
rect 8530 6210 8610 6230
rect 8930 6670 9010 6690
rect 8930 6630 8950 6670
rect 8990 6630 9010 6670
rect 8930 6570 9010 6630
rect 8930 6530 8950 6570
rect 8990 6530 9010 6570
rect 8930 6470 9010 6530
rect 8930 6430 8950 6470
rect 8990 6430 9010 6470
rect 8930 6370 9010 6430
rect 8930 6330 8950 6370
rect 8990 6330 9010 6370
rect 8930 6270 9010 6330
rect 8930 6230 8950 6270
rect 8990 6230 9010 6270
rect 8930 6210 9010 6230
rect 9330 6670 9410 6690
rect 9330 6630 9350 6670
rect 9390 6630 9410 6670
rect 9330 6570 9410 6630
rect 9330 6530 9350 6570
rect 9390 6530 9410 6570
rect 9330 6470 9410 6530
rect 9330 6430 9350 6470
rect 9390 6430 9410 6470
rect 9330 6370 9410 6430
rect 9330 6330 9350 6370
rect 9390 6330 9410 6370
rect 9330 6270 9410 6330
rect 9330 6230 9350 6270
rect 9390 6230 9410 6270
rect 9330 6210 9410 6230
rect 9730 6670 9810 6690
rect 9730 6630 9750 6670
rect 9790 6630 9810 6670
rect 9730 6570 9810 6630
rect 9730 6530 9750 6570
rect 9790 6530 9810 6570
rect 9730 6470 9810 6530
rect 9730 6430 9750 6470
rect 9790 6430 9810 6470
rect 9730 6370 9810 6430
rect 9730 6330 9750 6370
rect 9790 6330 9810 6370
rect 9730 6270 9810 6330
rect 9730 6230 9750 6270
rect 9790 6230 9810 6270
rect 9730 6210 9810 6230
rect 10130 6670 10210 6690
rect 10130 6630 10150 6670
rect 10190 6630 10210 6670
rect 10130 6570 10210 6630
rect 10130 6530 10150 6570
rect 10190 6530 10210 6570
rect 10130 6470 10210 6530
rect 10130 6430 10150 6470
rect 10190 6430 10210 6470
rect 10130 6370 10210 6430
rect 10130 6330 10150 6370
rect 10190 6330 10210 6370
rect 10130 6270 10210 6330
rect 10130 6230 10150 6270
rect 10190 6230 10210 6270
rect 10130 6210 10210 6230
rect 11750 5440 11850 5460
rect 11750 5380 11770 5440
rect 11830 5380 11850 5440
rect 11750 5360 11850 5380
rect 7660 5300 7740 5310
rect 7660 5240 7670 5300
rect 7730 5240 7740 5300
rect 7660 5230 7740 5240
rect 14230 5290 14310 5300
rect 14230 5230 14240 5290
rect 14300 5230 14310 5290
rect 7680 3900 7720 5230
rect 14230 5220 14310 5230
rect 13180 5190 13260 5200
rect 13180 5130 13190 5190
rect 13250 5130 13260 5190
rect 13180 5120 13260 5130
rect 11590 5090 11700 5110
rect 11590 5020 11610 5090
rect 11680 5020 11700 5090
rect 11590 5000 11700 5020
rect 7750 4560 11070 4580
rect 7750 4500 7770 4560
rect 7830 4520 7900 4560
rect 7940 4520 8000 4560
rect 8040 4520 8100 4560
rect 8140 4520 8200 4560
rect 8240 4520 8300 4560
rect 8340 4520 8400 4560
rect 8440 4520 8500 4560
rect 8540 4520 8600 4560
rect 8640 4520 8700 4560
rect 8740 4520 8800 4560
rect 8840 4520 8900 4560
rect 8940 4520 9000 4560
rect 9040 4520 9100 4560
rect 9140 4520 9200 4560
rect 9240 4520 9300 4560
rect 9340 4520 9400 4560
rect 9440 4520 9500 4560
rect 9540 4520 9600 4560
rect 9640 4520 9700 4560
rect 9740 4520 9800 4560
rect 9840 4520 9900 4560
rect 9940 4520 10000 4560
rect 10040 4520 10100 4560
rect 10140 4520 10200 4560
rect 10240 4520 10300 4560
rect 10340 4520 10400 4560
rect 10440 4520 10500 4560
rect 10540 4520 10600 4560
rect 10640 4520 10700 4560
rect 10740 4520 10800 4560
rect 10840 4520 10900 4560
rect 10940 4520 11000 4560
rect 11040 4520 11070 4560
rect 7830 4500 11070 4520
rect 7750 4480 7850 4500
rect 11350 3910 11460 3930
rect 7660 3890 7740 3900
rect 7660 3830 7670 3890
rect 7730 3830 7740 3890
rect 7660 3820 7740 3830
rect 8460 3890 8540 3900
rect 8460 3830 8470 3890
rect 8530 3830 8540 3890
rect 8460 3820 8540 3830
rect 9980 3880 10060 3900
rect 9980 3840 10000 3880
rect 10040 3840 10060 3880
rect 7550 3800 7630 3810
rect 7550 3740 7560 3800
rect 7620 3740 7630 3800
rect 1980 3700 7300 3710
rect 1900 3690 7300 3700
rect 7350 3730 7430 3740
rect 7550 3730 7630 3740
rect 8590 3800 8670 3810
rect 8590 3740 8600 3800
rect 8660 3740 8670 3800
rect 8590 3730 8670 3740
rect 1900 3680 2000 3690
rect 5830 3660 5870 3690
rect 7350 3670 7360 3730
rect 7420 3670 7430 3730
rect 7350 3660 7430 3670
rect 9980 3710 10060 3840
rect 11350 3840 11370 3910
rect 11440 3840 11460 3910
rect 11350 3820 11460 3840
rect 13200 3730 13240 5120
rect 2590 3640 2670 3660
rect 2590 3600 2610 3640
rect 2650 3630 2670 3640
rect 4120 3650 4200 3660
rect 4120 3630 4130 3650
rect 2650 3600 4130 3630
rect 2590 3590 4130 3600
rect 4190 3630 4200 3650
rect 5710 3650 5790 3660
rect 4190 3590 5180 3630
rect 2590 3580 2670 3590
rect 4120 3580 4200 3590
rect 3860 3080 3940 3090
rect 1610 3040 1690 3050
rect 1610 2980 1620 3040
rect 1680 3030 1690 3040
rect 2020 3030 2100 3050
rect 1680 3000 2040 3030
rect 1680 2980 1690 3000
rect 1610 2970 1690 2980
rect 2020 2990 2040 3000
rect 2080 2990 2100 3030
rect 3860 3020 3870 3080
rect 3930 3020 3940 3080
rect 3860 3010 3940 3020
rect 4940 3080 5020 3090
rect 4940 3020 4950 3080
rect 5010 3020 5020 3080
rect 4940 3010 5020 3020
rect 5140 3080 5180 3590
rect 5710 3590 5720 3650
rect 5780 3590 5790 3650
rect 5710 3580 5790 3590
rect 5830 3650 5910 3660
rect 5830 3590 5840 3650
rect 5900 3590 5910 3650
rect 9980 3650 9990 3710
rect 10050 3650 10060 3710
rect 11180 3720 11260 3730
rect 11180 3660 11190 3720
rect 11250 3660 11260 3720
rect 11180 3650 11260 3660
rect 13180 3720 13260 3730
rect 13180 3660 13190 3720
rect 13250 3660 13260 3720
rect 13180 3650 13260 3660
rect 9980 3640 10060 3650
rect 5830 3580 5910 3590
rect 6640 3620 6720 3630
rect 6640 3560 6650 3620
rect 6710 3560 6720 3620
rect 6640 3550 6720 3560
rect 7270 3620 7510 3630
rect 7270 3560 7280 3620
rect 7340 3560 7360 3620
rect 7420 3560 7440 3620
rect 7500 3560 7510 3620
rect 6890 3080 6970 3090
rect 5140 3060 5220 3080
rect 5140 3020 5160 3060
rect 5200 3020 5220 3060
rect 5140 3000 5220 3020
rect 6890 3020 6900 3080
rect 6960 3020 6970 3080
rect 6890 3010 6970 3020
rect 2020 2970 2100 2990
rect 1150 2400 1160 2460
rect 1220 2400 1240 2460
rect 1300 2400 1320 2460
rect 1380 2400 1390 2460
rect 1150 2380 1390 2400
rect 1150 2320 1160 2380
rect 1220 2320 1240 2380
rect 1300 2320 1320 2380
rect 1380 2320 1390 2380
rect 1150 2300 1390 2320
rect 1150 2240 1160 2300
rect 1220 2240 1240 2300
rect 1300 2240 1320 2300
rect 1380 2240 1390 2300
rect 1150 2230 1390 2240
rect 1630 1280 1670 2970
rect 5670 2690 5750 2700
rect 5670 2630 5680 2690
rect 5740 2630 5750 2690
rect 5670 2620 5750 2630
rect 5790 2690 5870 2700
rect 5790 2630 5800 2690
rect 5860 2630 5870 2690
rect 5790 2620 5870 2630
rect 6430 2690 6510 2700
rect 6430 2630 6440 2690
rect 6500 2630 6510 2690
rect 6430 2620 6510 2630
rect 1720 2590 1820 2610
rect 5710 2590 5750 2620
rect 7040 2590 7140 2600
rect 1720 2530 1740 2590
rect 1800 2580 7140 2590
rect 1800 2570 7060 2580
rect 1800 2530 1880 2570
rect 1920 2530 1980 2570
rect 2020 2530 2080 2570
rect 2120 2530 2180 2570
rect 2220 2530 2280 2570
rect 2320 2530 2380 2570
rect 2420 2530 2480 2570
rect 2520 2530 2580 2570
rect 2620 2530 2680 2570
rect 2720 2530 2780 2570
rect 2820 2530 2880 2570
rect 2920 2530 2980 2570
rect 3020 2530 3080 2570
rect 3120 2530 3180 2570
rect 3220 2530 3280 2570
rect 3320 2530 3380 2570
rect 3420 2530 3480 2570
rect 3520 2530 3580 2570
rect 3620 2530 3680 2570
rect 3720 2530 3780 2570
rect 3820 2530 3880 2570
rect 3920 2530 3980 2570
rect 4020 2530 4080 2570
rect 4120 2530 4180 2570
rect 4220 2530 4280 2570
rect 4320 2530 4380 2570
rect 4420 2530 4480 2570
rect 4520 2530 4580 2570
rect 4620 2530 4680 2570
rect 4720 2530 4780 2570
rect 4820 2530 4880 2570
rect 4920 2530 4980 2570
rect 5020 2530 5080 2570
rect 5120 2530 5180 2570
rect 5220 2530 5280 2570
rect 5320 2530 5380 2570
rect 5420 2530 5480 2570
rect 5520 2530 5580 2570
rect 5620 2530 5680 2570
rect 5720 2530 5780 2570
rect 5820 2530 5880 2570
rect 5920 2530 5980 2570
rect 6020 2530 6080 2570
rect 6120 2530 6180 2570
rect 6220 2530 6280 2570
rect 6320 2530 6380 2570
rect 6420 2530 6480 2570
rect 6520 2530 6580 2570
rect 6620 2530 6680 2570
rect 6720 2530 6780 2570
rect 6820 2530 6880 2570
rect 6920 2530 7060 2570
rect 1720 2520 7060 2530
rect 7120 2520 7140 2580
rect 1720 2510 7140 2520
rect 7040 2500 7140 2510
rect 7270 2460 7510 3560
rect 8390 3620 8470 3630
rect 8390 3560 8400 3620
rect 8460 3560 8470 3620
rect 8390 3550 8470 3560
rect 10420 3510 10500 3520
rect 7750 3500 7830 3510
rect 7750 3440 7760 3500
rect 7820 3440 7830 3500
rect 10420 3450 10430 3510
rect 10490 3450 10500 3510
rect 10420 3440 10500 3450
rect 11350 3500 11460 3520
rect 7750 3430 7830 3440
rect 11350 3430 11370 3500
rect 11440 3430 11460 3500
rect 7770 3090 7810 3430
rect 11350 3410 11460 3430
rect 7750 3080 7830 3090
rect 7750 3020 7760 3080
rect 7820 3020 7830 3080
rect 7750 3010 7830 3020
rect 7750 2860 7850 2880
rect 7750 2800 7770 2860
rect 7830 2840 11070 2860
rect 7830 2800 7910 2840
rect 7950 2800 8010 2840
rect 8050 2800 8110 2840
rect 8150 2800 8210 2840
rect 8250 2800 8310 2840
rect 8350 2800 8410 2840
rect 8450 2800 8510 2840
rect 8550 2800 8610 2840
rect 8650 2800 8710 2840
rect 8750 2800 8810 2840
rect 8850 2800 8910 2840
rect 8950 2800 9010 2840
rect 9050 2800 9110 2840
rect 9150 2800 9210 2840
rect 9250 2800 9310 2840
rect 9350 2800 9410 2840
rect 9450 2800 9510 2840
rect 9550 2800 9610 2840
rect 9650 2800 9710 2840
rect 9750 2800 9810 2840
rect 9850 2800 9910 2840
rect 9950 2800 10010 2840
rect 10050 2800 10110 2840
rect 10150 2800 10210 2840
rect 10250 2800 10310 2840
rect 10350 2800 10410 2840
rect 10450 2800 10510 2840
rect 10550 2800 10610 2840
rect 10650 2800 10710 2840
rect 10750 2800 10810 2840
rect 10850 2800 10910 2840
rect 10950 2800 11010 2840
rect 11050 2800 11070 2840
rect 7750 2780 11070 2800
rect 11700 2710 11810 2730
rect 11700 2640 11720 2710
rect 11790 2640 11810 2710
rect 11700 2620 11810 2640
rect 13200 2520 13240 3650
rect 17090 2730 17200 2750
rect 17090 2660 17110 2730
rect 17180 2660 17200 2730
rect 17090 2640 17200 2660
rect 17590 2730 17700 2750
rect 17590 2660 17610 2730
rect 17680 2660 17700 2730
rect 17590 2640 17700 2660
rect 14410 2520 14510 2540
rect 7270 2400 7280 2460
rect 7340 2400 7360 2460
rect 7420 2400 7440 2460
rect 7500 2400 7510 2460
rect 13180 2510 13260 2520
rect 13180 2450 13190 2510
rect 13250 2450 13260 2510
rect 13180 2440 13260 2450
rect 14300 2510 14430 2520
rect 14300 2450 14310 2510
rect 14370 2460 14430 2510
rect 14490 2510 14510 2520
rect 31480 2520 31580 2540
rect 31480 2510 31500 2520
rect 14490 2500 23180 2510
rect 14490 2460 23110 2500
rect 14370 2450 23110 2460
rect 23160 2450 23180 2500
rect 14300 2440 23180 2450
rect 25530 2500 31500 2510
rect 25530 2450 25552 2500
rect 25602 2460 31500 2500
rect 31560 2460 31580 2520
rect 25602 2450 31580 2460
rect 25530 2440 31580 2450
rect 7270 2380 7510 2400
rect 7270 2320 7280 2380
rect 7340 2320 7360 2380
rect 7420 2320 7440 2380
rect 7500 2320 7510 2380
rect 7270 2300 7510 2320
rect 7270 2240 7280 2300
rect 7340 2240 7360 2300
rect 7420 2240 7440 2300
rect 7500 2240 7510 2300
rect 7270 2230 7510 2240
rect 7040 2180 7140 2200
rect 7040 2120 7060 2180
rect 7120 2160 17420 2180
rect 7120 2120 7200 2160
rect 7240 2120 7300 2160
rect 7340 2120 7400 2160
rect 7440 2120 7500 2160
rect 7540 2120 7600 2160
rect 7640 2120 7700 2160
rect 7740 2120 7800 2160
rect 7840 2120 7900 2160
rect 7940 2120 8000 2160
rect 8040 2120 8100 2160
rect 8140 2120 8200 2160
rect 8240 2120 8300 2160
rect 8340 2120 8400 2160
rect 8440 2120 8500 2160
rect 8540 2120 8600 2160
rect 8640 2120 8700 2160
rect 8740 2120 8800 2160
rect 8840 2120 8900 2160
rect 8940 2120 9000 2160
rect 9040 2120 9100 2160
rect 9140 2120 9200 2160
rect 9240 2120 9300 2160
rect 9340 2120 9400 2160
rect 9440 2120 9500 2160
rect 9540 2120 9600 2160
rect 9640 2120 9700 2160
rect 9740 2120 9800 2160
rect 9840 2120 9900 2160
rect 9940 2120 10000 2160
rect 10040 2120 10100 2160
rect 10140 2120 10200 2160
rect 10240 2120 10300 2160
rect 10340 2120 10400 2160
rect 10440 2120 10500 2160
rect 10540 2120 10600 2160
rect 10640 2120 10700 2160
rect 10740 2120 10800 2160
rect 10840 2120 10900 2160
rect 10940 2120 11000 2160
rect 11040 2120 11100 2160
rect 11140 2120 11200 2160
rect 11240 2120 11300 2160
rect 11340 2120 11400 2160
rect 11440 2120 11500 2160
rect 11540 2120 11600 2160
rect 11640 2120 11700 2160
rect 11740 2120 11800 2160
rect 11840 2120 11900 2160
rect 11940 2120 12000 2160
rect 12040 2120 12100 2160
rect 12140 2120 12190 2160
rect 7040 2100 12190 2120
rect 12250 2120 12300 2160
rect 12340 2120 12400 2160
rect 12440 2120 12500 2160
rect 12540 2120 12600 2160
rect 12640 2120 12700 2160
rect 12740 2120 12800 2160
rect 12840 2120 12900 2160
rect 12940 2120 13000 2160
rect 13040 2120 13100 2160
rect 13140 2120 13200 2160
rect 13240 2120 13300 2160
rect 13340 2120 13400 2160
rect 13440 2120 13500 2160
rect 13540 2120 13600 2160
rect 13640 2120 13700 2160
rect 13740 2120 13800 2160
rect 13840 2120 13900 2160
rect 13940 2120 14000 2160
rect 14040 2120 14100 2160
rect 14140 2120 14200 2160
rect 14240 2120 14300 2160
rect 14340 2120 14400 2160
rect 14440 2120 14500 2160
rect 14540 2120 14600 2160
rect 14640 2120 14700 2160
rect 14740 2120 14800 2160
rect 14840 2120 14900 2160
rect 14940 2120 15000 2160
rect 15040 2120 15100 2160
rect 15140 2120 15200 2160
rect 15240 2120 15300 2160
rect 15340 2120 15400 2160
rect 15440 2120 15500 2160
rect 15540 2120 15600 2160
rect 15640 2120 15700 2160
rect 15740 2120 15800 2160
rect 15840 2120 15900 2160
rect 15940 2120 16000 2160
rect 16040 2120 16100 2160
rect 16140 2120 16200 2160
rect 16240 2120 16300 2160
rect 16340 2120 16400 2160
rect 16440 2120 16500 2160
rect 16540 2120 16600 2160
rect 16640 2120 16700 2160
rect 16740 2120 16800 2160
rect 16840 2120 16900 2160
rect 16940 2120 17000 2160
rect 17040 2120 17100 2160
rect 17140 2120 17200 2160
rect 17240 2120 17300 2160
rect 17340 2120 17420 2160
rect 12250 2100 17420 2120
rect 12170 2080 12270 2100
rect 12330 2030 14140 2070
rect 12170 1660 12270 1680
rect 1720 1640 12190 1660
rect 1720 1600 1770 1640
rect 1810 1600 1870 1640
rect 1910 1600 1970 1640
rect 2010 1600 2070 1640
rect 2110 1600 2170 1640
rect 2210 1600 2270 1640
rect 2310 1600 2370 1640
rect 2410 1600 2470 1640
rect 2510 1600 2570 1640
rect 2610 1600 2670 1640
rect 2710 1600 2770 1640
rect 2810 1600 2870 1640
rect 2910 1600 2970 1640
rect 3010 1600 3070 1640
rect 3110 1600 3170 1640
rect 3210 1600 3270 1640
rect 3310 1600 3370 1640
rect 3410 1600 3470 1640
rect 3510 1600 3570 1640
rect 3610 1600 3670 1640
rect 3710 1600 3770 1640
rect 3810 1600 3870 1640
rect 3910 1600 3970 1640
rect 4010 1600 4070 1640
rect 4110 1600 4170 1640
rect 4210 1600 4270 1640
rect 4310 1600 4370 1640
rect 4410 1600 4470 1640
rect 4510 1600 4570 1640
rect 4610 1600 4670 1640
rect 4710 1600 4770 1640
rect 4810 1600 4870 1640
rect 4910 1600 4970 1640
rect 5010 1600 5070 1640
rect 5110 1600 5170 1640
rect 5210 1600 5270 1640
rect 5310 1600 5370 1640
rect 5410 1600 5470 1640
rect 5510 1600 5570 1640
rect 5610 1600 5670 1640
rect 5710 1600 5770 1640
rect 5810 1600 5870 1640
rect 5910 1600 5970 1640
rect 6010 1600 6070 1640
rect 6110 1600 6170 1640
rect 6210 1600 6270 1640
rect 6310 1600 6370 1640
rect 6410 1600 6470 1640
rect 6510 1600 6570 1640
rect 6610 1600 6670 1640
rect 6710 1600 6770 1640
rect 6810 1600 6870 1640
rect 6910 1600 6970 1640
rect 7010 1600 7070 1640
rect 7110 1600 7170 1640
rect 7210 1600 7270 1640
rect 7310 1600 7370 1640
rect 7410 1600 7470 1640
rect 7510 1600 7570 1640
rect 7610 1600 7670 1640
rect 7710 1600 7770 1640
rect 7810 1600 7870 1640
rect 7910 1600 7970 1640
rect 8010 1600 8070 1640
rect 8110 1600 8170 1640
rect 8210 1600 8270 1640
rect 8310 1600 8370 1640
rect 8410 1600 8470 1640
rect 8510 1600 8570 1640
rect 8610 1600 8670 1640
rect 8710 1600 8770 1640
rect 8810 1600 8870 1640
rect 8910 1600 8970 1640
rect 9010 1600 9070 1640
rect 9110 1600 9170 1640
rect 9210 1600 9270 1640
rect 9310 1600 9370 1640
rect 9410 1600 9470 1640
rect 9510 1600 9570 1640
rect 9610 1600 9670 1640
rect 9710 1600 9770 1640
rect 9810 1600 9870 1640
rect 9910 1600 9970 1640
rect 10010 1600 10070 1640
rect 10110 1600 10170 1640
rect 10210 1600 10270 1640
rect 10310 1600 10370 1640
rect 10410 1600 10470 1640
rect 10510 1600 10570 1640
rect 10610 1600 10670 1640
rect 10710 1600 10770 1640
rect 10810 1600 10870 1640
rect 10910 1600 10970 1640
rect 11010 1600 11070 1640
rect 11110 1600 11170 1640
rect 11210 1600 11270 1640
rect 11310 1600 11370 1640
rect 11410 1600 11470 1640
rect 11510 1600 11570 1640
rect 11610 1600 11670 1640
rect 11710 1600 11770 1640
rect 11810 1600 11870 1640
rect 11910 1600 11970 1640
rect 12010 1600 12070 1640
rect 12110 1600 12190 1640
rect 12250 1600 12270 1660
rect 1720 1580 12270 1600
rect 1780 1530 1860 1550
rect 1780 1490 1800 1530
rect 1840 1510 2810 1530
rect 1840 1490 2750 1510
rect 1780 1470 1860 1490
rect 2730 1470 2750 1490
rect 2790 1470 2810 1510
rect 2860 1520 5440 1540
rect 2860 1480 2880 1520
rect 2920 1500 3820 1520
rect 2920 1480 2940 1500
rect 2860 1470 2940 1480
rect 3800 1480 3820 1500
rect 3860 1500 5380 1520
rect 3860 1480 3880 1500
rect 3800 1470 3880 1480
rect 5360 1480 5380 1500
rect 5420 1480 5440 1520
rect 7974 1530 8040 1550
rect 7974 1510 7984 1530
rect 5360 1470 5440 1480
rect 5630 1490 7984 1510
rect 8024 1490 8040 1530
rect 5630 1470 8040 1490
rect 2730 1450 2810 1470
rect 3390 1290 3470 1310
rect 1610 1270 1690 1280
rect 1610 1210 1620 1270
rect 1680 1210 1690 1270
rect 3390 1250 3410 1290
rect 3450 1280 3470 1290
rect 3910 1290 3990 1310
rect 3910 1280 3930 1290
rect 3450 1250 3930 1280
rect 3970 1250 3990 1290
rect 3390 1240 3990 1250
rect 5630 1300 5670 1470
rect 12330 1310 12370 2030
rect 12520 1640 12780 1660
rect 12520 1600 12530 1640
rect 12570 1600 12610 1640
rect 12650 1600 12780 1640
rect 12520 1580 12780 1600
rect 13120 1640 13380 1660
rect 13120 1600 13130 1640
rect 13170 1600 13210 1640
rect 13250 1600 13380 1640
rect 13120 1580 13380 1600
rect 13720 1640 13980 1660
rect 13720 1600 13730 1640
rect 13770 1600 13810 1640
rect 13850 1600 13980 1640
rect 13720 1580 13980 1600
rect 5630 1280 5710 1300
rect 5630 1240 5650 1280
rect 5690 1240 5710 1280
rect 5630 1220 5710 1240
rect 12290 1290 12370 1310
rect 12290 1250 12310 1290
rect 12350 1250 12370 1290
rect 12290 1230 12370 1250
rect 12630 1520 12710 1540
rect 12630 1480 12650 1520
rect 12690 1480 12710 1520
rect 12630 1460 12710 1480
rect 1610 1200 1690 1210
rect 4130 1090 4210 1110
rect 4130 1050 4150 1090
rect 4190 1050 4210 1090
rect 4130 1030 4210 1050
rect 2730 990 2810 1010
rect 4130 990 4170 1030
rect 8550 990 8590 1030
rect 9850 990 9890 1030
rect 11150 990 11190 1030
rect 2420 970 2690 990
rect 2420 930 2440 970
rect 2480 950 2630 970
rect 2480 930 2500 950
rect 2420 910 2500 930
rect 2620 930 2630 950
rect 2670 930 2690 970
rect 2730 950 2750 990
rect 2790 970 3620 990
rect 2790 950 3560 970
rect 2730 930 2810 950
rect 3540 930 3560 950
rect 3600 930 3620 970
rect 2620 910 2690 930
rect 3540 910 3620 930
rect 3680 970 4170 990
rect 3680 930 3690 970
rect 3730 950 4170 970
rect 4800 970 5100 990
rect 3730 930 3740 950
rect 3680 910 3740 930
rect 4800 930 4820 970
rect 4860 950 5040 970
rect 4860 930 4880 950
rect 4800 910 4880 930
rect 5020 930 5040 950
rect 5080 930 5100 970
rect 5020 910 5100 930
rect 6150 960 6640 980
rect 6150 920 6170 960
rect 6210 940 6580 960
rect 6210 920 6230 940
rect 6150 910 6230 920
rect 6560 920 6580 940
rect 6620 920 6640 960
rect 6560 910 6640 920
rect 8510 970 9170 990
rect 8510 930 8530 970
rect 8570 950 9110 970
rect 8570 930 8590 950
rect 8510 910 8590 930
rect 9090 930 9110 950
rect 9150 930 9170 970
rect 9090 910 9170 930
rect 9810 970 10470 990
rect 9810 930 9830 970
rect 9870 950 10410 970
rect 9870 930 9890 950
rect 9810 910 9890 930
rect 10390 930 10410 950
rect 10450 930 10470 970
rect 10390 910 10470 930
rect 11110 970 11770 990
rect 11110 930 11130 970
rect 11170 950 11710 970
rect 11170 930 11190 950
rect 11110 910 11190 930
rect 11690 930 11710 950
rect 11750 930 11770 970
rect 11690 910 11770 930
rect 1620 880 1720 900
rect 1620 820 1640 880
rect 1700 860 12270 880
rect 12630 870 12670 1460
rect 12740 990 12780 1580
rect 12700 970 12780 990
rect 12700 930 12720 970
rect 12760 930 12780 970
rect 12700 910 12780 930
rect 13230 1520 13310 1540
rect 13230 1480 13250 1520
rect 13290 1480 13310 1520
rect 13230 1460 13310 1480
rect 13230 870 13270 1460
rect 13340 990 13380 1580
rect 13300 970 13380 990
rect 13300 930 13320 970
rect 13360 930 13380 970
rect 13300 910 13380 930
rect 13830 1520 13910 1540
rect 13830 1480 13850 1520
rect 13890 1480 13910 1520
rect 13830 1460 13910 1480
rect 13830 870 13870 1460
rect 13940 990 13980 1580
rect 14100 1310 14140 2030
rect 14300 1820 14380 1830
rect 14300 1760 14310 1820
rect 14370 1760 14380 1820
rect 14300 1750 14380 1760
rect 14060 1290 14140 1310
rect 14060 1250 14080 1290
rect 14120 1250 14140 1290
rect 14060 1230 14140 1250
rect 13900 970 13980 990
rect 13900 930 13920 970
rect 13960 930 13980 970
rect 13900 910 13980 930
rect 1700 820 1770 860
rect 1810 820 1870 860
rect 1910 820 1970 860
rect 2010 820 2070 860
rect 2110 820 2170 860
rect 2210 820 2270 860
rect 2310 820 2370 860
rect 2410 820 2470 860
rect 2510 820 2570 860
rect 2610 820 2670 860
rect 2710 820 2770 860
rect 2810 820 2870 860
rect 2910 820 2970 860
rect 3010 820 3070 860
rect 3110 820 3170 860
rect 3210 820 3270 860
rect 3310 820 3370 860
rect 3410 820 3470 860
rect 3510 820 3570 860
rect 3610 820 3670 860
rect 3710 820 3770 860
rect 3810 820 3870 860
rect 3910 820 3970 860
rect 4010 820 4070 860
rect 4110 820 4170 860
rect 4210 820 4270 860
rect 4310 820 4370 860
rect 4410 820 4470 860
rect 4510 820 4570 860
rect 4610 820 4670 860
rect 4710 820 4770 860
rect 4810 820 4870 860
rect 4910 820 4970 860
rect 5010 820 5070 860
rect 5110 820 5170 860
rect 5210 820 5270 860
rect 5310 820 5370 860
rect 5410 820 5470 860
rect 5510 820 5570 860
rect 5610 820 5670 860
rect 5710 820 5770 860
rect 5810 820 5870 860
rect 5910 820 5970 860
rect 6010 820 6070 860
rect 6110 820 6170 860
rect 6210 820 6270 860
rect 6310 820 6370 860
rect 6410 820 6470 860
rect 6510 820 6570 860
rect 6610 820 6670 860
rect 6710 820 6770 860
rect 6810 820 6870 860
rect 6910 820 6970 860
rect 7010 820 7070 860
rect 7110 820 7170 860
rect 7210 820 7270 860
rect 7310 820 7370 860
rect 7410 820 7470 860
rect 7510 820 7570 860
rect 7610 820 7670 860
rect 7710 820 7770 860
rect 7810 820 7870 860
rect 7910 820 7970 860
rect 8010 820 8070 860
rect 8110 820 8170 860
rect 8210 820 8270 860
rect 8310 820 8370 860
rect 8410 820 8470 860
rect 8510 820 8570 860
rect 8610 820 8670 860
rect 8710 820 8770 860
rect 8810 820 8870 860
rect 8910 820 8970 860
rect 9010 820 9070 860
rect 9110 820 9170 860
rect 9210 820 9270 860
rect 9310 820 9370 860
rect 9410 820 9470 860
rect 9510 820 9570 860
rect 9610 820 9670 860
rect 9710 820 9770 860
rect 9810 820 9870 860
rect 9910 820 9970 860
rect 10010 820 10070 860
rect 10110 820 10170 860
rect 10210 820 10270 860
rect 10310 820 10370 860
rect 10410 820 10470 860
rect 10510 820 10570 860
rect 10610 820 10670 860
rect 10710 820 10770 860
rect 10810 820 10870 860
rect 10910 820 10970 860
rect 11010 820 11070 860
rect 11110 820 11170 860
rect 11210 820 11270 860
rect 11310 820 11370 860
rect 11410 820 11470 860
rect 11510 820 11570 860
rect 11610 820 11670 860
rect 11710 820 11770 860
rect 11810 820 11870 860
rect 11910 820 11970 860
rect 12010 820 12070 860
rect 12110 820 12190 860
rect 1620 800 12190 820
rect 12250 800 12270 860
rect 12170 780 12270 800
rect 12590 850 12670 870
rect 12590 810 12610 850
rect 12650 810 12670 850
rect 12590 750 12670 810
rect 12590 710 12610 750
rect 12650 710 12670 750
rect 12590 690 12670 710
rect 13190 850 13270 870
rect 13190 810 13210 850
rect 13250 810 13270 850
rect 13190 750 13270 810
rect 13190 710 13210 750
rect 13250 710 13270 750
rect 13190 690 13270 710
rect 13790 850 13870 870
rect 13790 810 13810 850
rect 13850 810 13870 850
rect 13790 750 13870 810
rect 13790 710 13810 750
rect 13850 710 13870 750
rect 13790 690 13870 710
rect 12170 80 12270 100
rect 12170 20 12190 80
rect 12250 60 14640 80
rect 12250 20 12300 60
rect 12340 20 12400 60
rect 12440 20 12500 60
rect 12540 20 12600 60
rect 12640 20 12700 60
rect 12740 20 12800 60
rect 12840 20 12900 60
rect 12940 20 13000 60
rect 13040 20 13100 60
rect 13140 20 13200 60
rect 13240 20 13300 60
rect 13340 20 13400 60
rect 13440 20 13500 60
rect 13540 20 13600 60
rect 13640 20 13700 60
rect 13740 20 13800 60
rect 13840 20 13900 60
rect 13940 20 14000 60
rect 14040 20 14100 60
rect 14140 20 14200 60
rect 14240 20 14300 60
rect 14340 20 14400 60
rect 14440 20 14500 60
rect 14540 20 14640 60
rect 12170 0 14640 20
<< via1 >>
rect 120 15140 180 15200
rect 490 15030 550 15090
rect 490 14950 550 15010
rect 490 14870 550 14930
rect 920 15030 980 15090
rect 920 14950 980 15010
rect 920 14870 980 14930
rect 910 14548 980 14558
rect 910 14498 920 14548
rect 920 14498 970 14548
rect 970 14498 980 14548
rect 910 14488 980 14498
rect 480 14398 550 14408
rect 480 14348 490 14398
rect 490 14348 540 14398
rect 540 14348 550 14398
rect 480 14338 550 14348
rect 120 14188 190 14198
rect 120 14138 130 14188
rect 130 14138 180 14188
rect 180 14138 190 14188
rect 120 14128 190 14138
rect 120 12840 190 12850
rect 120 12790 130 12840
rect 130 12790 180 12840
rect 180 12790 190 12840
rect 120 12780 190 12790
rect 10 10160 70 10220
rect 10 7040 70 7100
rect 240 12790 310 12800
rect 240 12740 250 12790
rect 250 12740 300 12790
rect 300 12740 310 12790
rect 240 12730 310 12740
rect 120 7530 180 7590
rect 670 12410 740 12420
rect 670 12360 680 12410
rect 680 12360 730 12410
rect 730 12360 740 12410
rect 670 12350 740 12360
rect 670 10670 730 10730
rect 240 8470 300 8530
rect 240 7150 300 7210
rect 350 10440 410 10500
rect 350 8700 410 8760
rect 120 5710 180 5770
rect 620 10330 680 10390
rect 7290 15140 7350 15200
rect 3240 15080 3300 15090
rect 3240 15040 3250 15080
rect 3250 15040 3290 15080
rect 3290 15040 3300 15080
rect 3240 15030 3300 15040
rect 3240 15000 3300 15010
rect 3240 14960 3250 15000
rect 3250 14960 3290 15000
rect 3290 14960 3300 15000
rect 3240 14950 3300 14960
rect 3240 14920 3300 14930
rect 3240 14880 3250 14920
rect 3250 14880 3290 14920
rect 3290 14880 3300 14920
rect 3240 14870 3300 14880
rect 5440 15030 5500 15090
rect 5440 14950 5500 15010
rect 5440 14870 5500 14930
rect 5800 15030 5860 15090
rect 5800 14950 5860 15010
rect 5800 14870 5860 14930
rect 5440 14548 5510 14558
rect 5440 14498 5450 14548
rect 5450 14498 5500 14548
rect 5500 14498 5510 14548
rect 5440 14488 5510 14498
rect 5800 14398 5870 14408
rect 5800 14348 5810 14398
rect 5810 14348 5860 14398
rect 5860 14348 5870 14398
rect 5800 14338 5870 14348
rect 5940 15030 6000 15090
rect 6020 15030 6080 15090
rect 5940 14950 6000 15010
rect 6020 14950 6080 15010
rect 5940 14870 6000 14930
rect 6020 14870 6080 14930
rect 1140 12760 1200 12820
rect 1570 12760 1630 12820
rect 3240 12764 3300 12820
rect 3240 12760 3244 12764
rect 3244 12760 3300 12764
rect 5800 13260 5870 13270
rect 5800 13210 5810 13260
rect 5810 13210 5860 13260
rect 5860 13210 5870 13260
rect 5800 13200 5870 13210
rect 5340 12760 5400 12820
rect 5680 12410 5750 12420
rect 5680 12360 5690 12410
rect 5690 12360 5740 12410
rect 5740 12360 5750 12410
rect 5680 12350 5750 12360
rect 5340 10750 5400 10810
rect 5690 10750 5750 10810
rect 3950 10670 4010 10730
rect 1140 10560 1200 10620
rect 2542 10610 2612 10620
rect 2542 10560 2552 10610
rect 2552 10560 2602 10610
rect 2602 10560 2612 10610
rect 2542 10550 2612 10560
rect 3940 10610 4010 10620
rect 3940 10560 3950 10610
rect 3950 10560 4000 10610
rect 4000 10560 4010 10610
rect 3940 10550 4010 10560
rect 5810 10440 5870 10500
rect 1030 10330 1090 10390
rect 1080 10210 1140 10220
rect 1080 10170 1090 10210
rect 1090 10170 1130 10210
rect 1130 10170 1140 10210
rect 1080 10160 1140 10170
rect 5470 10250 5530 10260
rect 5470 10210 5480 10250
rect 5480 10210 5520 10250
rect 5520 10210 5530 10250
rect 5470 10200 5530 10210
rect 5470 10170 5530 10180
rect 5470 10130 5480 10170
rect 5480 10130 5520 10170
rect 5520 10130 5530 10170
rect 5470 10120 5530 10130
rect 7290 14800 7350 14860
rect 6460 14398 6530 14408
rect 6460 14348 6470 14398
rect 6470 14348 6520 14398
rect 6520 14348 6530 14398
rect 6460 14338 6530 14348
rect 6840 14340 6910 14410
rect 6460 13052 6530 13062
rect 6460 13002 6470 13052
rect 6470 13002 6520 13052
rect 6520 13002 6530 13052
rect 6460 12992 6530 13002
rect 6470 12700 6530 12760
rect 6240 10750 6300 10810
rect 6150 10550 6210 10610
rect 5940 10200 6000 10260
rect 6020 10200 6080 10260
rect 5940 10120 6000 10180
rect 6020 10120 6080 10180
rect 1160 10040 1220 10050
rect 1160 10000 1170 10040
rect 1170 10000 1210 10040
rect 1210 10000 1220 10040
rect 1160 9990 1220 10000
rect 1320 10040 1380 10050
rect 1320 10000 1330 10040
rect 1330 10000 1370 10040
rect 1370 10000 1380 10040
rect 1320 9990 1380 10000
rect 1480 10040 1540 10050
rect 1480 10000 1490 10040
rect 1490 10000 1530 10040
rect 1530 10000 1540 10040
rect 1480 9990 1540 10000
rect 1640 10040 1700 10050
rect 1640 10000 1650 10040
rect 1650 10000 1690 10040
rect 1690 10000 1700 10040
rect 1640 9990 1700 10000
rect 1800 10040 1860 10050
rect 1800 10000 1810 10040
rect 1810 10000 1850 10040
rect 1850 10000 1860 10040
rect 1800 9990 1860 10000
rect 1960 10040 2020 10050
rect 1960 10000 1970 10040
rect 1970 10000 2010 10040
rect 2010 10000 2020 10040
rect 1960 9990 2020 10000
rect 2120 10040 2180 10050
rect 2120 10000 2130 10040
rect 2130 10000 2170 10040
rect 2170 10000 2180 10040
rect 2120 9990 2180 10000
rect 2280 10040 2340 10050
rect 2280 10000 2290 10040
rect 2290 10000 2330 10040
rect 2330 10000 2340 10040
rect 2280 9990 2340 10000
rect 2440 10040 2500 10050
rect 2440 10000 2450 10040
rect 2450 10000 2490 10040
rect 2490 10000 2500 10040
rect 2440 9990 2500 10000
rect 2600 10040 2660 10050
rect 2600 10000 2610 10040
rect 2610 10000 2650 10040
rect 2650 10000 2660 10040
rect 2600 9990 2660 10000
rect 2760 10040 2820 10050
rect 2760 10000 2770 10040
rect 2770 10000 2810 10040
rect 2810 10000 2820 10040
rect 2760 9990 2820 10000
rect 2920 10040 2980 10050
rect 2920 10000 2930 10040
rect 2930 10000 2970 10040
rect 2970 10000 2980 10040
rect 2920 9990 2980 10000
rect 3080 10040 3140 10050
rect 3080 10000 3090 10040
rect 3090 10000 3130 10040
rect 3130 10000 3140 10040
rect 3080 9990 3140 10000
rect 3240 10040 3300 10050
rect 3240 10000 3250 10040
rect 3250 10000 3290 10040
rect 3290 10000 3300 10040
rect 3240 9990 3300 10000
rect 3400 10040 3460 10050
rect 3400 10000 3410 10040
rect 3410 10000 3450 10040
rect 3450 10000 3460 10040
rect 3400 9990 3460 10000
rect 3560 10040 3620 10050
rect 3560 10000 3570 10040
rect 3570 10000 3610 10040
rect 3610 10000 3620 10040
rect 3560 9990 3620 10000
rect 3720 10040 3780 10050
rect 3720 10000 3730 10040
rect 3730 10000 3770 10040
rect 3770 10000 3780 10040
rect 3720 9990 3780 10000
rect 3880 10040 3940 10050
rect 3880 10000 3890 10040
rect 3890 10000 3930 10040
rect 3930 10000 3940 10040
rect 3880 9990 3940 10000
rect 4040 10040 4100 10050
rect 4040 10000 4050 10040
rect 4050 10000 4090 10040
rect 4090 10000 4100 10040
rect 4040 9990 4100 10000
rect 4200 10040 4260 10050
rect 4200 10000 4210 10040
rect 4210 10000 4250 10040
rect 4250 10000 4260 10040
rect 4200 9990 4260 10000
rect 4360 10040 4420 10050
rect 4360 10000 4370 10040
rect 4370 10000 4410 10040
rect 4410 10000 4420 10040
rect 4360 9990 4420 10000
rect 4520 10040 4580 10050
rect 4520 10000 4530 10040
rect 4530 10000 4570 10040
rect 4570 10000 4580 10040
rect 4520 9990 4580 10000
rect 4680 10040 4740 10050
rect 4680 10000 4690 10040
rect 4690 10000 4730 10040
rect 4730 10000 4740 10040
rect 4680 9990 4740 10000
rect 4840 10040 4900 10050
rect 4840 10000 4850 10040
rect 4850 10000 4890 10040
rect 4890 10000 4900 10040
rect 4840 9990 4900 10000
rect 5000 10040 5060 10050
rect 5000 10000 5010 10040
rect 5010 10000 5050 10040
rect 5050 10000 5060 10040
rect 5000 9990 5060 10000
rect 5160 10040 5220 10050
rect 5160 10000 5170 10040
rect 5170 10000 5210 10040
rect 5210 10000 5220 10040
rect 5160 9990 5220 10000
rect 1900 9880 1960 9940
rect 1900 9800 1960 9860
rect 1900 9770 1960 9780
rect 1900 9730 1910 9770
rect 1910 9730 1950 9770
rect 1950 9730 1960 9770
rect 1900 9720 1960 9730
rect 3160 9880 3220 9940
rect 3240 9880 3300 9940
rect 3320 9880 3380 9940
rect 3160 9800 3220 9860
rect 3240 9800 3300 9860
rect 3320 9800 3380 9860
rect 3160 9720 3220 9780
rect 3240 9720 3300 9780
rect 3320 9720 3380 9780
rect 920 9130 980 9140
rect 920 9090 930 9130
rect 930 9090 970 9130
rect 970 9090 980 9130
rect 920 9080 980 9090
rect 920 9000 980 9060
rect 920 8920 980 8980
rect 1160 9130 1220 9140
rect 1160 9090 1170 9130
rect 1170 9090 1210 9130
rect 1210 9090 1220 9130
rect 1160 9080 1220 9090
rect 1160 9000 1220 9060
rect 1160 8920 1220 8980
rect 1400 9130 1460 9140
rect 1400 9090 1410 9130
rect 1410 9090 1450 9130
rect 1450 9090 1460 9130
rect 1400 9080 1460 9090
rect 1400 9000 1460 9060
rect 1400 8920 1460 8980
rect 1640 9130 1700 9140
rect 1640 9090 1650 9130
rect 1650 9090 1690 9130
rect 1690 9090 1700 9130
rect 1640 9080 1700 9090
rect 1640 9000 1700 9060
rect 1640 8920 1700 8980
rect 2280 9130 2340 9140
rect 2280 9090 2290 9130
rect 2290 9090 2330 9130
rect 2330 9090 2340 9130
rect 2280 9080 2340 9090
rect 2280 9000 2340 9060
rect 2280 8920 2340 8980
rect 2520 9130 2580 9140
rect 2520 9090 2530 9130
rect 2530 9090 2570 9130
rect 2570 9090 2580 9130
rect 2520 9080 2580 9090
rect 2520 9000 2580 9060
rect 2520 8920 2580 8980
rect 2760 9130 2820 9140
rect 2760 9090 2770 9130
rect 2770 9090 2810 9130
rect 2810 9090 2820 9130
rect 2760 9080 2820 9090
rect 2760 9000 2820 9060
rect 2760 8920 2820 8980
rect 740 8810 800 8870
rect 1490 8810 1550 8870
rect 1710 8810 1770 8870
rect 1970 8810 2030 8870
rect 2190 8810 2250 8870
rect 2450 8810 2510 8870
rect 1423 8752 1475 8760
rect 1423 8718 1433 8752
rect 1433 8718 1467 8752
rect 1467 8718 1475 8752
rect 1423 8708 1475 8718
rect 1783 8752 1835 8760
rect 1783 8718 1793 8752
rect 1793 8718 1827 8752
rect 1827 8718 1835 8752
rect 1783 8708 1835 8718
rect 1903 8752 1955 8760
rect 1903 8718 1913 8752
rect 1913 8718 1947 8752
rect 1947 8718 1955 8752
rect 1903 8708 1955 8718
rect 2263 8752 2315 8760
rect 2263 8718 2273 8752
rect 2273 8718 2307 8752
rect 2307 8718 2315 8752
rect 2263 8708 2315 8718
rect 2383 8752 2435 8760
rect 2383 8718 2393 8752
rect 2393 8718 2427 8752
rect 2427 8718 2435 8752
rect 2383 8708 2435 8718
rect 2800 8730 2860 8740
rect 2800 8690 2810 8730
rect 2810 8690 2850 8730
rect 2850 8690 2860 8730
rect 2800 8680 2860 8690
rect 2800 8650 2860 8660
rect 2800 8610 2810 8650
rect 2810 8610 2850 8650
rect 2850 8610 2860 8650
rect 2800 8600 2860 8610
rect 1526 8522 1578 8532
rect 1526 8488 1534 8522
rect 1534 8488 1568 8522
rect 1568 8488 1578 8522
rect 1526 8480 1578 8488
rect 1684 8522 1736 8532
rect 1684 8488 1692 8522
rect 1692 8488 1726 8522
rect 1726 8488 1736 8522
rect 1684 8480 1736 8488
rect 1600 8370 1660 8430
rect 1360 8260 1420 8320
rect 620 7990 680 8050
rect 700 7990 760 8050
rect 1120 7990 1180 8050
rect 1360 7990 1420 8050
rect 880 7920 940 7930
rect 880 7880 890 7920
rect 890 7880 930 7920
rect 930 7880 940 7920
rect 880 7870 940 7880
rect 640 7530 700 7590
rect 2008 8522 2060 8532
rect 2008 8488 2016 8522
rect 2016 8488 2050 8522
rect 2050 8488 2060 8522
rect 2008 8480 2060 8488
rect 2162 8522 2214 8532
rect 2162 8488 2170 8522
rect 2170 8488 2204 8522
rect 2204 8488 2214 8522
rect 2162 8480 2214 8488
rect 2080 8370 2140 8430
rect 2486 8522 2538 8532
rect 2486 8488 2494 8522
rect 2494 8488 2528 8522
rect 2528 8488 2538 8522
rect 2486 8480 2538 8488
rect 2800 8570 2860 8580
rect 2800 8530 2810 8570
rect 2810 8530 2850 8570
rect 2850 8530 2860 8570
rect 2800 8520 2860 8530
rect 2560 8370 2620 8430
rect 1840 8260 1900 8320
rect 2320 8260 2380 8320
rect 1840 7990 1900 8050
rect 2080 7990 2140 8050
rect 2560 7990 2620 8050
rect 2740 7990 2800 8050
rect 1600 7920 1660 7930
rect 1600 7880 1610 7920
rect 1610 7880 1650 7920
rect 1650 7880 1660 7920
rect 1600 7870 1660 7880
rect 1360 7530 1420 7590
rect 2320 7920 2380 7930
rect 2320 7880 2330 7920
rect 2330 7880 2370 7920
rect 2370 7880 2380 7920
rect 2320 7870 2380 7880
rect 2080 7530 2140 7590
rect 2800 7530 2860 7590
rect 4580 9880 4640 9940
rect 4580 9800 4640 9860
rect 4580 9770 4640 9780
rect 4580 9730 4590 9770
rect 4590 9730 4630 9770
rect 4630 9730 4640 9770
rect 4580 9720 4640 9730
rect 3160 8680 3220 8740
rect 3240 8680 3300 8740
rect 3320 8680 3380 8740
rect 3160 8600 3220 8660
rect 3240 8600 3300 8660
rect 3320 8600 3380 8660
rect 3160 8520 3220 8580
rect 3240 8520 3300 8580
rect 3320 8520 3380 8580
rect 3720 9130 3780 9140
rect 3720 9090 3730 9130
rect 3730 9090 3770 9130
rect 3770 9090 3780 9130
rect 3720 9080 3780 9090
rect 3720 9000 3780 9060
rect 3720 8920 3780 8980
rect 3960 9130 4020 9140
rect 3960 9090 3970 9130
rect 3970 9090 4010 9130
rect 4010 9090 4020 9130
rect 3960 9080 4020 9090
rect 3960 9000 4020 9060
rect 3960 8920 4020 8980
rect 4200 9130 4260 9140
rect 4200 9090 4210 9130
rect 4210 9090 4250 9130
rect 4250 9090 4260 9130
rect 4200 9080 4260 9090
rect 4200 9000 4260 9060
rect 4200 8920 4260 8980
rect 4840 9130 4900 9140
rect 4840 9090 4850 9130
rect 4850 9090 4890 9130
rect 4890 9090 4900 9130
rect 4840 9080 4900 9090
rect 4840 9000 4900 9060
rect 4840 8920 4900 8980
rect 5080 9130 5140 9140
rect 5080 9090 5090 9130
rect 5090 9090 5130 9130
rect 5130 9090 5140 9130
rect 5080 9080 5140 9090
rect 5080 9000 5140 9060
rect 5080 8920 5140 8980
rect 5320 9130 5380 9140
rect 5320 9090 5330 9130
rect 5330 9090 5370 9130
rect 5370 9090 5380 9130
rect 5320 9080 5380 9090
rect 5320 9000 5380 9060
rect 5320 8920 5380 8980
rect 5560 9130 5620 9140
rect 5560 9090 5570 9130
rect 5570 9090 5610 9130
rect 5610 9090 5620 9130
rect 5560 9080 5620 9090
rect 5560 9000 5620 9060
rect 5560 8920 5620 8980
rect 4030 8810 4090 8870
rect 4290 8810 4350 8870
rect 4510 8810 4570 8870
rect 4770 8810 4830 8870
rect 4990 8810 5050 8870
rect 5740 8810 5800 8870
rect 3680 8730 3740 8740
rect 3680 8690 3690 8730
rect 3690 8690 3730 8730
rect 3730 8690 3740 8730
rect 3680 8680 3740 8690
rect 4105 8752 4157 8760
rect 4105 8718 4113 8752
rect 4113 8718 4147 8752
rect 4147 8718 4157 8752
rect 4105 8708 4157 8718
rect 4225 8752 4277 8760
rect 4225 8718 4233 8752
rect 4233 8718 4267 8752
rect 4267 8718 4277 8752
rect 4225 8708 4277 8718
rect 4585 8752 4637 8760
rect 4585 8718 4593 8752
rect 4593 8718 4627 8752
rect 4627 8718 4637 8752
rect 4585 8708 4637 8718
rect 4705 8752 4757 8760
rect 4705 8718 4713 8752
rect 4713 8718 4747 8752
rect 4747 8718 4757 8752
rect 4705 8708 4757 8718
rect 5065 8752 5117 8760
rect 5065 8718 5073 8752
rect 5073 8718 5107 8752
rect 5107 8718 5117 8752
rect 5065 8708 5117 8718
rect 6150 8700 6210 8760
rect 3680 8650 3740 8660
rect 3680 8610 3690 8650
rect 3690 8610 3730 8650
rect 3730 8610 3740 8650
rect 3680 8600 3740 8610
rect 3680 8570 3740 8580
rect 3680 8530 3690 8570
rect 3690 8530 3730 8570
rect 3730 8530 3740 8570
rect 3680 8520 3740 8530
rect 4002 8522 4054 8532
rect 4002 8488 4012 8522
rect 4012 8488 4046 8522
rect 4046 8488 4054 8522
rect 4002 8480 4054 8488
rect 3920 8370 3980 8430
rect 4326 8522 4378 8532
rect 4326 8488 4336 8522
rect 4336 8488 4370 8522
rect 4370 8488 4378 8522
rect 4326 8480 4378 8488
rect 4480 8522 4532 8532
rect 4480 8488 4490 8522
rect 4490 8488 4524 8522
rect 4524 8488 4532 8522
rect 4480 8480 4532 8488
rect 4400 8370 4460 8430
rect 4804 8522 4856 8532
rect 4804 8488 4814 8522
rect 4814 8488 4848 8522
rect 4848 8488 4856 8522
rect 4804 8480 4856 8488
rect 4962 8522 5014 8532
rect 4962 8488 4972 8522
rect 4972 8488 5006 8522
rect 5006 8488 5014 8522
rect 4962 8480 5014 8488
rect 4880 8370 4940 8430
rect 4160 8260 4220 8320
rect 4640 8260 4700 8320
rect 3740 8150 3800 8210
rect 3740 8070 3800 8130
rect 3740 7990 3800 8050
rect 3920 8150 3980 8210
rect 3920 8070 3980 8130
rect 3920 7990 3980 8050
rect 4160 8150 4220 8210
rect 4160 8070 4220 8130
rect 4160 7990 4220 8050
rect 4400 8150 4460 8210
rect 4400 8070 4460 8130
rect 4400 7990 4460 8050
rect 4640 8150 4700 8210
rect 4640 8070 4700 8130
rect 4640 7990 4700 8050
rect 3060 7530 3120 7590
rect 3420 7530 3480 7590
rect 520 7420 580 7480
rect 520 7340 580 7400
rect 520 7260 580 7320
rect 760 7420 820 7480
rect 760 7340 820 7400
rect 760 7260 820 7320
rect 1000 7420 1060 7480
rect 1000 7340 1060 7400
rect 1000 7260 1060 7320
rect 1240 7420 1300 7480
rect 1240 7340 1300 7400
rect 1240 7260 1300 7320
rect 1480 7420 1540 7480
rect 1480 7340 1540 7400
rect 1480 7260 1540 7320
rect 1720 7420 1780 7480
rect 1720 7340 1780 7400
rect 1720 7260 1780 7320
rect 1960 7420 2020 7480
rect 1960 7340 2020 7400
rect 1960 7260 2020 7320
rect 2200 7420 2260 7480
rect 2200 7340 2260 7400
rect 2200 7260 2260 7320
rect 2440 7420 2500 7480
rect 2440 7340 2500 7400
rect 2440 7260 2500 7320
rect 2680 7420 2740 7480
rect 2680 7340 2740 7400
rect 2680 7260 2740 7320
rect 2920 7420 2980 7480
rect 2920 7340 2980 7400
rect 2920 7260 2980 7320
rect 1800 7150 1860 7210
rect 3240 7150 3300 7210
rect 2160 7040 2220 7100
rect 1890 6760 1950 6770
rect 1890 6720 1900 6760
rect 1900 6720 1940 6760
rect 1940 6720 1950 6760
rect 1890 6710 1950 6720
rect 2070 6760 2130 6770
rect 2070 6720 2080 6760
rect 2080 6720 2120 6760
rect 2120 6720 2130 6760
rect 2070 6710 2130 6720
rect 2520 6930 2580 6990
rect 2250 6760 2310 6770
rect 2250 6720 2260 6760
rect 2260 6720 2300 6760
rect 2300 6720 2310 6760
rect 2250 6710 2310 6720
rect 2430 6760 2490 6770
rect 2430 6720 2440 6760
rect 2440 6720 2480 6760
rect 2480 6720 2490 6760
rect 2430 6710 2490 6720
rect 2880 6820 2940 6880
rect 2610 6760 2670 6770
rect 2610 6720 2620 6760
rect 2620 6720 2660 6760
rect 2660 6720 2670 6760
rect 2610 6710 2670 6720
rect 2790 6760 2850 6770
rect 2790 6720 2800 6760
rect 2800 6720 2840 6760
rect 2840 6720 2850 6760
rect 2790 6710 2850 6720
rect 2970 6760 3030 6770
rect 2970 6720 2980 6760
rect 2980 6720 3020 6760
rect 3020 6720 3030 6760
rect 2970 6710 3030 6720
rect 3150 6760 3210 6770
rect 3150 6720 3160 6760
rect 3160 6720 3200 6760
rect 3200 6720 3210 6760
rect 3150 6710 3210 6720
rect 3680 7530 3740 7590
rect 4160 7920 4220 7930
rect 4160 7880 4170 7920
rect 4170 7880 4210 7920
rect 4210 7880 4220 7920
rect 4160 7870 4220 7880
rect 4400 7530 4460 7590
rect 5120 8260 5180 8320
rect 5120 8150 5180 8210
rect 5120 8070 5180 8130
rect 5120 7990 5180 8050
rect 5360 8150 5420 8210
rect 5360 8070 5420 8130
rect 5360 7990 5420 8050
rect 5780 8150 5840 8210
rect 5780 8070 5840 8130
rect 5780 7990 5840 8050
rect 4880 7920 4940 7930
rect 4880 7880 4890 7920
rect 4890 7880 4930 7920
rect 4930 7880 4940 7920
rect 4880 7870 4940 7880
rect 5120 7530 5180 7590
rect 5600 7920 5660 7930
rect 5600 7880 5610 7920
rect 5610 7880 5650 7920
rect 5650 7880 5660 7920
rect 5600 7870 5660 7880
rect 5840 7530 5900 7590
rect 3560 7420 3620 7480
rect 3560 7340 3620 7400
rect 3560 7260 3620 7320
rect 3800 7420 3860 7480
rect 3800 7340 3860 7400
rect 3800 7260 3860 7320
rect 4040 7420 4100 7480
rect 4040 7340 4100 7400
rect 4040 7260 4100 7320
rect 4280 7420 4340 7480
rect 4280 7340 4340 7400
rect 4280 7260 4340 7320
rect 4520 7420 4580 7480
rect 4520 7340 4580 7400
rect 4520 7260 4580 7320
rect 4760 7420 4820 7480
rect 4760 7340 4820 7400
rect 4760 7260 4820 7320
rect 5000 7420 5060 7480
rect 5000 7340 5060 7400
rect 5000 7260 5060 7320
rect 5240 7420 5300 7480
rect 5240 7340 5300 7400
rect 5240 7260 5300 7320
rect 5480 7420 5540 7480
rect 5480 7340 5540 7400
rect 5480 7260 5540 7320
rect 5720 7420 5780 7480
rect 5720 7340 5780 7400
rect 5720 7260 5780 7320
rect 4680 7150 4740 7210
rect 4320 7040 4380 7100
rect 3960 6930 4020 6990
rect 3600 6820 3660 6880
rect 3330 6760 3390 6770
rect 3330 6720 3340 6760
rect 3340 6720 3380 6760
rect 3380 6720 3390 6760
rect 3330 6710 3390 6720
rect 3420 6710 3480 6770
rect 3510 6760 3570 6770
rect 3510 6720 3520 6760
rect 3520 6720 3560 6760
rect 3560 6720 3570 6760
rect 3510 6710 3570 6720
rect 3690 6760 3750 6770
rect 3690 6720 3700 6760
rect 3700 6720 3740 6760
rect 3740 6720 3750 6760
rect 3690 6710 3750 6720
rect 3870 6760 3930 6770
rect 3870 6720 3880 6760
rect 3880 6720 3920 6760
rect 3920 6720 3930 6760
rect 3870 6710 3930 6720
rect 4050 6760 4110 6770
rect 4050 6720 4060 6760
rect 4060 6720 4100 6760
rect 4100 6720 4110 6760
rect 4050 6710 4110 6720
rect 4230 6760 4290 6770
rect 4230 6720 4240 6760
rect 4240 6720 4280 6760
rect 4280 6720 4290 6760
rect 4230 6710 4290 6720
rect 4410 6760 4470 6770
rect 4410 6720 4420 6760
rect 4420 6720 4460 6760
rect 4460 6720 4470 6760
rect 4410 6710 4470 6720
rect 4590 6760 4650 6770
rect 4590 6720 4600 6760
rect 4600 6720 4640 6760
rect 4640 6720 4650 6760
rect 4590 6710 4650 6720
rect 5710 7040 5770 7100
rect 5240 6930 5300 6990
rect 5590 6560 5650 6570
rect 5590 6520 5600 6560
rect 5600 6520 5640 6560
rect 5640 6520 5650 6560
rect 5590 6510 5650 6520
rect 5960 7420 6020 7480
rect 5960 7340 6020 7400
rect 5960 7260 6020 7320
rect 6240 8470 6300 8530
rect 6970 14100 7030 14160
rect 6850 12000 6910 12060
rect 6580 11300 6640 11360
rect 6660 11300 6720 11360
rect 6740 11300 6800 11360
rect 7220 13400 7280 13460
rect 7090 12700 7150 12760
rect 7090 11300 7150 11360
rect 6970 10330 7030 10390
rect 11770 9750 11830 9810
rect 7220 9050 7280 9110
rect 7220 8950 7280 9010
rect 6580 8150 6640 8210
rect 6660 8150 6720 8210
rect 6740 8150 6800 8210
rect 9800 8270 9860 8280
rect 9800 8230 9810 8270
rect 9810 8230 9850 8270
rect 9850 8230 9860 8270
rect 9800 8220 9860 8230
rect 6580 8070 6640 8130
rect 6660 8070 6720 8130
rect 6740 8070 6800 8130
rect 7850 8100 7910 8160
rect 6580 7990 6640 8050
rect 6660 7990 6720 8050
rect 6740 7990 6800 8050
rect 9800 8050 9860 8060
rect 9800 8010 9810 8050
rect 9810 8010 9850 8050
rect 9850 8010 9860 8050
rect 9800 8000 9860 8010
rect 11770 7810 11840 7880
rect 7560 7650 7620 7710
rect 8080 7640 8140 7700
rect 8900 7660 8960 7720
rect 9580 7770 9640 7780
rect 9580 7730 9590 7770
rect 9590 7730 9630 7770
rect 9630 7730 9640 7770
rect 9580 7720 9640 7730
rect 6470 7530 6530 7590
rect 7450 7480 7510 7540
rect 6240 6930 6300 6990
rect 6150 6820 6210 6880
rect 5830 6560 5890 6570
rect 5830 6520 5840 6560
rect 5840 6520 5880 6560
rect 5880 6520 5890 6560
rect 5830 6510 5890 6520
rect 5240 6170 5300 6230
rect 5710 6220 5770 6230
rect 5710 6180 5720 6220
rect 5720 6180 5760 6220
rect 5760 6180 5770 6220
rect 5710 6170 5770 6180
rect 1620 6020 1680 6030
rect 1620 5980 1630 6020
rect 1630 5980 1670 6020
rect 1670 5980 1680 6020
rect 1620 5970 1680 5980
rect 1620 5890 1680 5950
rect 1620 5810 1680 5870
rect 1980 6020 2040 6030
rect 1980 5980 1990 6020
rect 1990 5980 2030 6020
rect 2030 5980 2040 6020
rect 1980 5970 2040 5980
rect 1980 5890 2040 5950
rect 1980 5810 2040 5870
rect 2340 6020 2400 6030
rect 2340 5980 2350 6020
rect 2350 5980 2390 6020
rect 2390 5980 2400 6020
rect 2340 5970 2400 5980
rect 2340 5890 2400 5950
rect 2340 5810 2400 5870
rect 2700 6020 2760 6030
rect 2700 5980 2710 6020
rect 2710 5980 2750 6020
rect 2750 5980 2760 6020
rect 2700 5970 2760 5980
rect 2700 5890 2760 5950
rect 2700 5810 2760 5870
rect 3060 6020 3120 6030
rect 3060 5980 3070 6020
rect 3070 5980 3110 6020
rect 3110 5980 3120 6020
rect 3060 5970 3120 5980
rect 3060 5890 3120 5950
rect 3060 5810 3120 5870
rect 3420 6020 3480 6030
rect 3420 5980 3430 6020
rect 3430 5980 3470 6020
rect 3470 5980 3480 6020
rect 3420 5970 3480 5980
rect 3420 5890 3480 5950
rect 3420 5810 3480 5870
rect 3780 6020 3840 6030
rect 3780 5980 3790 6020
rect 3790 5980 3830 6020
rect 3830 5980 3840 6020
rect 3780 5970 3840 5980
rect 3780 5890 3840 5950
rect 3780 5810 3840 5870
rect 4140 6020 4200 6030
rect 4140 5980 4150 6020
rect 4150 5980 4190 6020
rect 4190 5980 4200 6020
rect 4140 5970 4200 5980
rect 4140 5890 4200 5950
rect 4140 5810 4200 5870
rect 4500 6020 4560 6030
rect 4500 5980 4510 6020
rect 4510 5980 4550 6020
rect 4550 5980 4560 6020
rect 4500 5970 4560 5980
rect 4500 5890 4560 5950
rect 4500 5810 4560 5870
rect 4860 6020 4920 6030
rect 4860 5980 4870 6020
rect 4870 5980 4910 6020
rect 4910 5980 4920 6020
rect 4860 5970 4920 5980
rect 4860 5890 4920 5950
rect 4860 5810 4920 5870
rect 5490 5970 5550 6030
rect 5490 5890 5550 5950
rect 5490 5810 5550 5870
rect 5930 5970 5990 6030
rect 5930 5890 5990 5950
rect 5930 5810 5990 5870
rect 1798 5752 1850 5760
rect 1798 5718 1808 5752
rect 1808 5718 1842 5752
rect 1842 5718 1850 5752
rect 1798 5708 1850 5718
rect 1908 5752 1960 5760
rect 1908 5718 1918 5752
rect 1918 5718 1952 5752
rect 1952 5718 1960 5752
rect 1908 5708 1960 5718
rect 2018 5752 2070 5760
rect 2018 5718 2028 5752
rect 2028 5718 2062 5752
rect 2062 5718 2070 5752
rect 2018 5708 2070 5718
rect 2128 5752 2180 5760
rect 2128 5718 2138 5752
rect 2138 5718 2172 5752
rect 2172 5718 2180 5752
rect 2128 5708 2180 5718
rect 2238 5752 2290 5760
rect 2238 5718 2248 5752
rect 2248 5718 2282 5752
rect 2282 5718 2290 5752
rect 2238 5708 2290 5718
rect 2348 5752 2400 5760
rect 2348 5718 2358 5752
rect 2358 5718 2392 5752
rect 2392 5718 2400 5752
rect 2348 5708 2400 5718
rect 2458 5752 2510 5760
rect 2458 5718 2468 5752
rect 2468 5718 2502 5752
rect 2502 5718 2510 5752
rect 2458 5708 2510 5718
rect 2568 5752 2620 5760
rect 2568 5718 2578 5752
rect 2578 5718 2612 5752
rect 2612 5718 2620 5752
rect 2568 5708 2620 5718
rect 2678 5752 2730 5760
rect 2678 5718 2688 5752
rect 2688 5718 2722 5752
rect 2722 5718 2730 5752
rect 2678 5708 2730 5718
rect 2788 5752 2840 5760
rect 2788 5718 2798 5752
rect 2798 5718 2832 5752
rect 2832 5718 2840 5752
rect 2788 5708 2840 5718
rect 3698 5752 3750 5760
rect 3698 5718 3708 5752
rect 3708 5718 3742 5752
rect 3742 5718 3750 5752
rect 3698 5708 3750 5718
rect 3808 5752 3860 5760
rect 3808 5718 3818 5752
rect 3818 5718 3852 5752
rect 3852 5718 3860 5752
rect 3808 5708 3860 5718
rect 3918 5752 3970 5760
rect 3918 5718 3928 5752
rect 3928 5718 3962 5752
rect 3962 5718 3970 5752
rect 3918 5708 3970 5718
rect 4028 5752 4080 5760
rect 4028 5718 4038 5752
rect 4038 5718 4072 5752
rect 4072 5718 4080 5752
rect 4028 5708 4080 5718
rect 4138 5752 4190 5760
rect 4138 5718 4148 5752
rect 4148 5718 4182 5752
rect 4182 5718 4190 5752
rect 4138 5708 4190 5718
rect 4248 5752 4300 5760
rect 4248 5718 4258 5752
rect 4258 5718 4292 5752
rect 4292 5718 4300 5752
rect 4248 5708 4300 5718
rect 4358 5752 4410 5760
rect 4358 5718 4368 5752
rect 4368 5718 4402 5752
rect 4402 5718 4410 5752
rect 4358 5708 4410 5718
rect 4468 5752 4520 5760
rect 4468 5718 4478 5752
rect 4478 5718 4512 5752
rect 4512 5718 4520 5752
rect 4468 5708 4520 5718
rect 4578 5752 4630 5760
rect 4578 5718 4588 5752
rect 4588 5718 4622 5752
rect 4622 5718 4630 5752
rect 4578 5708 4630 5718
rect 4688 5752 4740 5760
rect 4688 5718 4698 5752
rect 4698 5718 4732 5752
rect 4732 5718 4740 5752
rect 4688 5708 4740 5718
rect 1630 5420 1690 5430
rect 1630 5380 1640 5420
rect 1640 5380 1680 5420
rect 1680 5380 1690 5420
rect 1630 5370 1690 5380
rect 1850 5370 1910 5430
rect 2070 5370 2130 5430
rect 2290 5370 2350 5430
rect 2510 5370 2570 5430
rect 2730 5370 2790 5430
rect 2950 5420 3010 5430
rect 2950 5380 2960 5420
rect 2960 5380 3000 5420
rect 3000 5380 3010 5420
rect 2950 5370 3010 5380
rect 3530 5420 3590 5430
rect 3530 5380 3540 5420
rect 3540 5380 3580 5420
rect 3580 5380 3590 5420
rect 3530 5370 3590 5380
rect 3750 5370 3810 5430
rect 3970 5370 4030 5430
rect 4190 5370 4250 5430
rect 4410 5370 4470 5430
rect 4630 5370 4690 5430
rect 4850 5420 4910 5430
rect 4850 5380 4860 5420
rect 4860 5380 4900 5420
rect 4900 5380 4910 5420
rect 4850 5370 4910 5380
rect 350 5260 410 5320
rect 1740 5260 1800 5320
rect 1960 5260 2020 5320
rect 2180 5260 2240 5320
rect 2400 5260 2460 5320
rect 2620 5260 2680 5320
rect 2840 5260 2900 5320
rect 3640 5260 3700 5320
rect 1160 5150 1220 5210
rect 1240 5150 1300 5210
rect 1320 5150 1380 5210
rect 1160 5070 1220 5130
rect 1240 5070 1300 5130
rect 1320 5070 1380 5130
rect 1160 4990 1220 5050
rect 1240 4990 1300 5050
rect 1320 4990 1380 5050
rect 3640 5150 3700 5210
rect 3640 5070 3700 5130
rect 3640 4990 3700 5050
rect 3860 5260 3920 5320
rect 3860 5150 3920 5210
rect 3860 5070 3920 5130
rect 3860 4990 3920 5050
rect 4080 5260 4140 5320
rect 4080 5150 4140 5210
rect 4080 5070 4140 5130
rect 4080 4990 4140 5050
rect 4300 5260 4360 5320
rect 4300 5150 4360 5210
rect 4300 5070 4360 5130
rect 4300 4990 4360 5050
rect 4520 5260 4580 5320
rect 4520 5150 4580 5210
rect 4520 5070 4580 5130
rect 4520 4990 4580 5050
rect 4740 5260 4800 5320
rect 4740 5150 4800 5210
rect 4740 5070 4800 5130
rect 7450 5130 7510 5190
rect 4740 4990 4800 5050
rect 7360 5020 7420 5080
rect 1740 4920 1800 4930
rect 1740 4880 1750 4920
rect 1750 4880 1790 4920
rect 1790 4880 1800 4920
rect 7060 4880 7120 4940
rect 1740 4870 1800 4880
rect 6350 4820 6410 4830
rect 6350 4780 6360 4820
rect 6360 4780 6400 4820
rect 6400 4780 6410 4820
rect 6350 4770 6410 4780
rect 1940 4470 2000 4480
rect 1940 4430 1950 4470
rect 1950 4430 1990 4470
rect 1990 4430 2000 4470
rect 1940 4420 2000 4430
rect 3850 4470 3910 4480
rect 3850 4430 3860 4470
rect 3860 4430 3900 4470
rect 3900 4430 3910 4470
rect 3850 4420 3910 4430
rect 7450 4770 7510 4830
rect 6650 4640 6710 4700
rect 7360 4640 7420 4700
rect 5020 4430 5080 4440
rect 5020 4390 5030 4430
rect 5030 4390 5070 4430
rect 5070 4390 5080 4430
rect 5020 4380 5080 4390
rect 6650 4400 6710 4410
rect 6650 4360 6660 4400
rect 6660 4360 6700 4400
rect 6700 4360 6710 4400
rect 6650 4350 6710 4360
rect 6890 4400 6950 4410
rect 6890 4360 6900 4400
rect 6900 4360 6940 4400
rect 6940 4360 6950 4400
rect 6890 4350 6950 4360
rect 7360 4350 7420 4410
rect 4150 3860 4210 3870
rect 4150 3820 4160 3860
rect 4160 3820 4200 3860
rect 4200 3820 4210 3860
rect 4150 3810 4210 3820
rect 7220 3760 7280 3770
rect 1920 3700 1980 3760
rect 7220 3720 7230 3760
rect 7230 3720 7270 3760
rect 7270 3720 7280 3760
rect 7220 3710 7280 3720
rect 7450 3830 7510 3890
rect 8080 7480 8140 7540
rect 8440 7500 8500 7560
rect 9580 7490 9640 7550
rect 14240 7550 14300 7610
rect 8440 7440 8500 7450
rect 8440 7400 8450 7440
rect 8450 7400 8490 7440
rect 8490 7400 8500 7440
rect 8440 7390 8500 7400
rect 8880 7440 8940 7450
rect 8880 7400 8890 7440
rect 8890 7400 8930 7440
rect 8930 7400 8940 7440
rect 8880 7390 8940 7400
rect 11770 7310 11840 7380
rect 8760 7060 8820 7070
rect 8760 7020 8770 7060
rect 8770 7020 8810 7060
rect 8810 7020 8820 7060
rect 8760 7010 8820 7020
rect 7850 6910 7910 6970
rect 8760 6840 8820 6850
rect 8760 6800 8770 6840
rect 8770 6800 8810 6840
rect 8810 6800 8820 6840
rect 8760 6790 8820 6800
rect 11770 5380 11830 5440
rect 7670 5240 7730 5300
rect 14240 5230 14300 5290
rect 13190 5130 13250 5190
rect 11610 5020 11680 5090
rect 7770 4500 7830 4560
rect 7670 3830 7730 3890
rect 8470 3880 8530 3890
rect 8470 3840 8480 3880
rect 8480 3840 8520 3880
rect 8520 3840 8530 3880
rect 8470 3830 8530 3840
rect 7560 3740 7620 3800
rect 8600 3790 8660 3800
rect 8600 3750 8610 3790
rect 8610 3750 8650 3790
rect 8650 3750 8660 3790
rect 8600 3740 8660 3750
rect 7360 3670 7420 3730
rect 11370 3840 11440 3910
rect 4130 3590 4190 3650
rect 1620 2980 1680 3040
rect 3870 3070 3930 3080
rect 3870 3030 3880 3070
rect 3880 3030 3920 3070
rect 3920 3030 3930 3070
rect 3870 3020 3930 3030
rect 4950 3070 5010 3080
rect 4950 3030 4960 3070
rect 4960 3030 5000 3070
rect 5000 3030 5010 3070
rect 4950 3020 5010 3030
rect 5720 3640 5780 3650
rect 5720 3600 5730 3640
rect 5730 3600 5770 3640
rect 5770 3600 5780 3640
rect 5720 3590 5780 3600
rect 5840 3590 5900 3650
rect 9990 3650 10050 3710
rect 11190 3710 11250 3720
rect 11190 3670 11200 3710
rect 11200 3670 11240 3710
rect 11240 3670 11250 3710
rect 11190 3660 11250 3670
rect 13190 3660 13250 3720
rect 6650 3610 6710 3620
rect 6650 3570 6660 3610
rect 6660 3570 6700 3610
rect 6700 3570 6710 3610
rect 6650 3560 6710 3570
rect 7280 3560 7340 3620
rect 7360 3560 7420 3620
rect 7440 3560 7500 3620
rect 6900 3070 6960 3080
rect 6900 3030 6910 3070
rect 6910 3030 6950 3070
rect 6950 3030 6960 3070
rect 6900 3020 6960 3030
rect 1160 2400 1220 2460
rect 1240 2400 1300 2460
rect 1320 2400 1380 2460
rect 1160 2320 1220 2380
rect 1240 2320 1300 2380
rect 1320 2320 1380 2380
rect 1160 2240 1220 2300
rect 1240 2240 1300 2300
rect 1320 2240 1380 2300
rect 5680 2630 5740 2690
rect 5800 2680 5860 2690
rect 5800 2640 5810 2680
rect 5810 2640 5850 2680
rect 5850 2640 5860 2680
rect 5800 2630 5860 2640
rect 6440 2680 6500 2690
rect 6440 2640 6450 2680
rect 6450 2640 6490 2680
rect 6490 2640 6500 2680
rect 6440 2630 6500 2640
rect 1740 2580 1800 2590
rect 1740 2540 1750 2580
rect 1750 2540 1790 2580
rect 1790 2540 1800 2580
rect 1740 2530 1800 2540
rect 7060 2520 7120 2580
rect 8400 3610 8460 3620
rect 8400 3570 8410 3610
rect 8410 3570 8450 3610
rect 8450 3570 8460 3610
rect 8400 3560 8460 3570
rect 7760 3440 7820 3500
rect 10430 3500 10490 3510
rect 10430 3460 10440 3500
rect 10440 3460 10480 3500
rect 10480 3460 10490 3500
rect 10430 3450 10490 3460
rect 11370 3430 11440 3500
rect 7760 3020 7820 3080
rect 7770 2800 7830 2860
rect 11720 2640 11790 2710
rect 17110 2660 17180 2730
rect 17610 2660 17680 2730
rect 7280 2400 7340 2460
rect 7360 2400 7420 2460
rect 7440 2400 7500 2460
rect 13190 2450 13250 2510
rect 14310 2450 14370 2510
rect 14430 2460 14490 2520
rect 31500 2460 31560 2520
rect 7280 2320 7340 2380
rect 7360 2320 7420 2380
rect 7440 2320 7500 2380
rect 7280 2240 7340 2300
rect 7360 2240 7420 2300
rect 7440 2240 7500 2300
rect 7060 2120 7120 2180
rect 12190 2100 12250 2160
rect 12190 1600 12250 1660
rect 1620 1260 1680 1270
rect 1620 1220 1630 1260
rect 1630 1220 1670 1260
rect 1670 1220 1680 1260
rect 1620 1210 1680 1220
rect 1640 820 1700 880
rect 14310 1810 14370 1820
rect 14310 1770 14320 1810
rect 14320 1770 14360 1810
rect 14360 1770 14370 1810
rect 14310 1760 14370 1770
rect 12190 800 12250 860
rect 12190 20 12250 80
<< metal2 >>
rect 110 15200 7360 15210
rect 110 15140 120 15200
rect 180 15140 7290 15200
rect 7350 15140 7360 15200
rect 110 15130 7360 15140
rect 480 15090 6090 15100
rect 480 15030 490 15090
rect 550 15030 920 15090
rect 980 15030 3240 15090
rect 3300 15030 5440 15090
rect 5500 15030 5800 15090
rect 5860 15030 5940 15090
rect 6000 15030 6020 15090
rect 6080 15030 6090 15090
rect 480 15010 6090 15030
rect 480 14950 490 15010
rect 550 14950 920 15010
rect 980 14950 3240 15010
rect 3300 14950 5440 15010
rect 5500 14950 5800 15010
rect 5860 14950 5940 15010
rect 6000 14950 6020 15010
rect 6080 14950 6090 15010
rect 480 14930 6090 14950
rect 480 14870 490 14930
rect 550 14870 920 14930
rect 980 14870 3240 14930
rect 3300 14870 5440 14930
rect 5500 14870 5800 14930
rect 5860 14870 5940 14930
rect 6000 14870 6020 14930
rect 6080 14870 6090 14930
rect 480 14860 6090 14870
rect 7280 14860 7360 14870
rect 7280 14800 7290 14860
rect 7350 14800 7360 14860
rect 7280 14790 7360 14800
rect 930 14568 970 14570
rect 5450 14568 5490 14570
rect 910 14558 980 14568
rect 910 14478 980 14488
rect 5440 14558 5510 14568
rect 5440 14478 5510 14488
rect 500 14418 540 14420
rect 5810 14418 5850 14420
rect 480 14408 550 14418
rect 480 14328 550 14338
rect 5800 14408 5870 14418
rect 5800 14328 5870 14338
rect 6460 14410 6920 14420
rect 6460 14408 6840 14410
rect 6530 14340 6840 14408
rect 6910 14340 6920 14410
rect 6530 14338 6920 14340
rect 6460 14330 6920 14338
rect 6460 14328 6530 14330
rect 130 14208 170 14210
rect 120 14198 190 14208
rect 120 14118 190 14128
rect 6950 14160 7050 14180
rect 6950 14100 6970 14160
rect 7030 14100 7050 14160
rect 6950 14080 7050 14100
rect 7210 13460 7290 13470
rect 7210 13400 7220 13460
rect 7280 13400 7290 13460
rect 7210 13390 7290 13400
rect 5800 13270 5870 13280
rect 5800 13190 5870 13200
rect 6460 13062 6530 13072
rect 6460 12980 6530 12992
rect 120 12850 190 12870
rect 1130 12820 1640 12830
rect 120 12770 190 12780
rect 240 12800 310 12810
rect 1130 12760 1140 12820
rect 1200 12760 1570 12820
rect 1630 12760 1640 12820
rect 1130 12750 1640 12760
rect 3230 12820 5410 12830
rect 3230 12760 3240 12820
rect 3300 12760 5340 12820
rect 5400 12760 5410 12820
rect 3230 12750 5410 12760
rect 6460 12760 7170 12780
rect 240 12720 310 12730
rect 6460 12700 6470 12760
rect 6530 12700 7090 12760
rect 7150 12700 7170 12760
rect 6460 12680 7170 12700
rect 670 12420 740 12430
rect 670 12340 740 12350
rect 5680 12420 5750 12430
rect 5680 12340 5750 12350
rect 6840 12060 7360 12070
rect 6840 12000 6850 12060
rect 6910 12000 7290 12060
rect 7350 12000 7360 12060
rect 6840 11990 7360 12000
rect 6570 11360 7170 11380
rect 6570 11300 6580 11360
rect 6640 11300 6660 11360
rect 6720 11300 6740 11360
rect 6800 11300 7090 11360
rect 7150 11300 7170 11360
rect 6570 11280 7170 11300
rect 5330 10810 5410 10820
rect 5330 10750 5340 10810
rect 5400 10800 5410 10810
rect 5680 10810 5760 10820
rect 5680 10800 5690 10810
rect 5400 10760 5690 10800
rect 5400 10750 5410 10760
rect 5330 10740 5410 10750
rect 5680 10750 5690 10760
rect 5750 10800 5760 10810
rect 6230 10810 6310 10820
rect 6230 10800 6240 10810
rect 5750 10760 6240 10800
rect 5750 10750 5760 10760
rect 5680 10740 5760 10750
rect 6230 10750 6240 10760
rect 6300 10750 6310 10810
rect 6230 10740 6310 10750
rect 660 10730 4020 10740
rect 660 10670 670 10730
rect 730 10670 3950 10730
rect 4010 10670 4020 10730
rect 660 10660 4020 10670
rect 1130 10620 2540 10630
rect 1130 10560 1140 10620
rect 1200 10560 2542 10620
rect 1130 10550 2542 10560
rect 2612 10550 2622 10620
rect 3930 10550 3940 10620
rect 4010 10600 4020 10620
rect 6140 10610 6220 10620
rect 6140 10600 6150 10610
rect 4010 10560 6150 10600
rect 4010 10550 4020 10560
rect 6140 10550 6150 10560
rect 6210 10550 6220 10610
rect 6140 10540 6220 10550
rect 340 10500 5880 10510
rect 340 10440 350 10500
rect 410 10440 5810 10500
rect 5870 10440 5880 10500
rect 340 10430 5880 10440
rect 610 10390 7040 10400
rect 610 10330 620 10390
rect 680 10330 1030 10390
rect 1090 10330 6970 10390
rect 7030 10330 7040 10390
rect 610 10320 7040 10330
rect 5460 10260 7140 10270
rect 0 10220 1150 10230
rect 0 10160 10 10220
rect 70 10160 1080 10220
rect 1140 10160 1150 10220
rect 0 10150 1150 10160
rect 5460 10200 5470 10260
rect 5530 10200 5940 10260
rect 6000 10200 6020 10260
rect 6080 10220 7140 10260
rect 6080 10200 7060 10220
rect 5460 10180 7060 10200
rect 5460 10120 5470 10180
rect 5530 10120 5940 10180
rect 6000 10120 6020 10180
rect 6080 10160 7060 10180
rect 7120 10160 7140 10220
rect 6080 10120 7140 10160
rect 5460 10110 7140 10120
rect 1150 10050 1230 10060
rect 1150 9990 1160 10050
rect 1220 10040 1230 10050
rect 1310 10050 1390 10060
rect 1310 10040 1320 10050
rect 1220 10000 1320 10040
rect 1220 9990 1230 10000
rect 1150 9980 1230 9990
rect 1310 9990 1320 10000
rect 1380 10040 1390 10050
rect 1470 10050 1550 10060
rect 1470 10040 1480 10050
rect 1380 10000 1480 10040
rect 1380 9990 1390 10000
rect 1310 9980 1390 9990
rect 1470 9990 1480 10000
rect 1540 10040 1550 10050
rect 1630 10050 1710 10060
rect 1630 10040 1640 10050
rect 1540 10000 1640 10040
rect 1540 9990 1550 10000
rect 1470 9980 1550 9990
rect 1630 9990 1640 10000
rect 1700 10040 1710 10050
rect 1790 10050 1870 10060
rect 1790 10040 1800 10050
rect 1700 10000 1800 10040
rect 1700 9990 1710 10000
rect 1630 9980 1710 9990
rect 1790 9990 1800 10000
rect 1860 10040 1870 10050
rect 1950 10050 2030 10060
rect 1950 10040 1960 10050
rect 1860 10000 1960 10040
rect 1860 9990 1870 10000
rect 1790 9980 1870 9990
rect 1950 9990 1960 10000
rect 2020 10040 2030 10050
rect 2110 10050 2190 10060
rect 2110 10040 2120 10050
rect 2020 10000 2120 10040
rect 2020 9990 2030 10000
rect 1950 9980 2030 9990
rect 2110 9990 2120 10000
rect 2180 10040 2190 10050
rect 2270 10050 2350 10060
rect 2270 10040 2280 10050
rect 2180 10000 2280 10040
rect 2180 9990 2190 10000
rect 2110 9980 2190 9990
rect 2270 9990 2280 10000
rect 2340 10040 2350 10050
rect 2430 10050 2510 10060
rect 2430 10040 2440 10050
rect 2340 10000 2440 10040
rect 2340 9990 2350 10000
rect 2270 9980 2350 9990
rect 2430 9990 2440 10000
rect 2500 10040 2510 10050
rect 2590 10050 2670 10060
rect 2590 10040 2600 10050
rect 2500 10000 2600 10040
rect 2500 9990 2510 10000
rect 2430 9980 2510 9990
rect 2590 9990 2600 10000
rect 2660 10040 2670 10050
rect 2750 10050 2830 10060
rect 2750 10040 2760 10050
rect 2660 10000 2760 10040
rect 2660 9990 2670 10000
rect 2590 9980 2670 9990
rect 2750 9990 2760 10000
rect 2820 10040 2830 10050
rect 2910 10050 2990 10060
rect 2910 10040 2920 10050
rect 2820 10000 2920 10040
rect 2820 9990 2830 10000
rect 2750 9980 2830 9990
rect 2910 9990 2920 10000
rect 2980 10040 2990 10050
rect 3070 10050 3150 10060
rect 3070 10040 3080 10050
rect 2980 10000 3080 10040
rect 2980 9990 2990 10000
rect 2910 9980 2990 9990
rect 3070 9990 3080 10000
rect 3140 9990 3150 10050
rect 3070 9980 3150 9990
rect 3230 10050 3310 10060
rect 3230 9990 3240 10050
rect 3300 10040 3310 10050
rect 3390 10050 3470 10060
rect 3390 10040 3400 10050
rect 3300 10000 3400 10040
rect 3300 9990 3310 10000
rect 3230 9980 3310 9990
rect 3390 9990 3400 10000
rect 3460 10040 3470 10050
rect 3550 10050 3630 10060
rect 3550 10040 3560 10050
rect 3460 10000 3560 10040
rect 3460 9990 3470 10000
rect 3390 9980 3470 9990
rect 3550 9990 3560 10000
rect 3620 10040 3630 10050
rect 3710 10050 3790 10060
rect 3710 10040 3720 10050
rect 3620 10000 3720 10040
rect 3620 9990 3630 10000
rect 3550 9980 3630 9990
rect 3710 9990 3720 10000
rect 3780 10040 3790 10050
rect 3870 10050 3950 10060
rect 3870 10040 3880 10050
rect 3780 10000 3880 10040
rect 3780 9990 3790 10000
rect 3710 9980 3790 9990
rect 3870 9990 3880 10000
rect 3940 10040 3950 10050
rect 4030 10050 4110 10060
rect 4030 10040 4040 10050
rect 3940 10000 4040 10040
rect 3940 9990 3950 10000
rect 3870 9980 3950 9990
rect 4030 9990 4040 10000
rect 4100 10040 4110 10050
rect 4190 10050 4270 10060
rect 4190 10040 4200 10050
rect 4100 10000 4200 10040
rect 4100 9990 4110 10000
rect 4030 9980 4110 9990
rect 4190 9990 4200 10000
rect 4260 10040 4270 10050
rect 4350 10050 4430 10060
rect 4350 10040 4360 10050
rect 4260 10000 4360 10040
rect 4260 9990 4270 10000
rect 4190 9980 4270 9990
rect 4350 9990 4360 10000
rect 4420 10040 4430 10050
rect 4510 10050 4590 10060
rect 4510 10040 4520 10050
rect 4420 10000 4520 10040
rect 4420 9990 4430 10000
rect 4350 9980 4430 9990
rect 4510 9990 4520 10000
rect 4580 10040 4590 10050
rect 4670 10050 4750 10060
rect 4670 10040 4680 10050
rect 4580 10000 4680 10040
rect 4580 9990 4590 10000
rect 4510 9980 4590 9990
rect 4670 9990 4680 10000
rect 4740 10040 4750 10050
rect 4830 10050 4910 10060
rect 4830 10040 4840 10050
rect 4740 10000 4840 10040
rect 4740 9990 4750 10000
rect 4670 9980 4750 9990
rect 4830 9990 4840 10000
rect 4900 10040 4910 10050
rect 4990 10050 5070 10060
rect 4990 10040 5000 10050
rect 4900 10000 5000 10040
rect 4900 9990 4910 10000
rect 4830 9980 4910 9990
rect 4990 9990 5000 10000
rect 5060 10040 5070 10050
rect 5150 10050 5230 10060
rect 5150 10040 5160 10050
rect 5060 10000 5160 10040
rect 5060 9990 5070 10000
rect 4990 9980 5070 9990
rect 5150 9990 5160 10000
rect 5220 9990 5230 10050
rect 5150 9980 5230 9990
rect 1890 9940 7140 9950
rect 1890 9880 1900 9940
rect 1960 9880 3160 9940
rect 3220 9880 3240 9940
rect 3300 9880 3320 9940
rect 3380 9880 4580 9940
rect 4640 9910 7140 9940
rect 4640 9880 7060 9910
rect 1890 9860 7060 9880
rect 1890 9800 1900 9860
rect 1960 9800 3160 9860
rect 3220 9800 3240 9860
rect 3300 9800 3320 9860
rect 3380 9800 4580 9860
rect 4640 9850 7060 9860
rect 7120 9850 7140 9910
rect 4640 9810 7140 9850
rect 4640 9800 7060 9810
rect 1890 9780 7060 9800
rect 1890 9720 1900 9780
rect 1960 9720 3160 9780
rect 3220 9720 3240 9780
rect 3300 9720 3320 9780
rect 3380 9720 4580 9780
rect 4640 9750 7060 9780
rect 7120 9750 7140 9810
rect 4640 9720 7140 9750
rect 11750 9810 11850 9830
rect 11750 9750 11770 9810
rect 11830 9750 11850 9810
rect 11750 9730 11850 9750
rect 1890 9710 7140 9720
rect 910 9140 7300 9150
rect 910 9080 920 9140
rect 980 9080 1160 9140
rect 1220 9080 1400 9140
rect 1460 9080 1640 9140
rect 1700 9080 2280 9140
rect 2340 9080 2520 9140
rect 2580 9080 2760 9140
rect 2820 9080 3720 9140
rect 3780 9080 3960 9140
rect 4020 9080 4200 9140
rect 4260 9080 4840 9140
rect 4900 9080 5080 9140
rect 5140 9080 5320 9140
rect 5380 9080 5560 9140
rect 5620 9110 7300 9140
rect 5620 9080 7220 9110
rect 910 9060 7220 9080
rect 910 9000 920 9060
rect 980 9000 1160 9060
rect 1220 9000 1400 9060
rect 1460 9000 1640 9060
rect 1700 9000 2280 9060
rect 2340 9000 2520 9060
rect 2580 9000 2760 9060
rect 2820 9000 3720 9060
rect 3780 9000 3960 9060
rect 4020 9000 4200 9060
rect 4260 9000 4840 9060
rect 4900 9000 5080 9060
rect 5140 9000 5320 9060
rect 5380 9000 5560 9060
rect 5620 9050 7220 9060
rect 7280 9050 7300 9110
rect 5620 9010 7300 9050
rect 5620 9000 7220 9010
rect 910 8980 7220 9000
rect 910 8920 920 8980
rect 980 8920 1160 8980
rect 1220 8920 1400 8980
rect 1460 8920 1640 8980
rect 1700 8920 2280 8980
rect 2340 8920 2520 8980
rect 2580 8920 2760 8980
rect 2820 8920 3720 8980
rect 3780 8920 3960 8980
rect 4020 8920 4200 8980
rect 4260 8920 4840 8980
rect 4900 8920 5080 8980
rect 5140 8920 5320 8980
rect 5380 8920 5560 8980
rect 5620 8950 7220 8980
rect 7280 8950 7300 9010
rect 5620 8920 7300 8950
rect 910 8910 7300 8920
rect 730 8870 2520 8880
rect 730 8810 740 8870
rect 800 8810 1490 8870
rect 1550 8810 1710 8870
rect 1770 8810 1970 8870
rect 2030 8810 2190 8870
rect 2250 8810 2450 8870
rect 2510 8810 2520 8870
rect 730 8800 2520 8810
rect 4020 8870 5810 8880
rect 4020 8810 4030 8870
rect 4090 8810 4290 8870
rect 4350 8810 4510 8870
rect 4570 8810 4770 8870
rect 4830 8810 4990 8870
rect 5050 8810 5740 8870
rect 5800 8810 5810 8870
rect 4020 8800 5810 8810
rect 340 8760 2439 8770
rect 340 8700 350 8760
rect 410 8708 1423 8760
rect 1475 8708 1783 8760
rect 1835 8708 1903 8760
rect 1955 8708 2263 8760
rect 2315 8708 2383 8760
rect 2435 8708 2439 8760
rect 4101 8760 6220 8770
rect 410 8700 2439 8708
rect 2790 8740 3750 8750
rect 340 8690 420 8700
rect 2790 8680 2800 8740
rect 2860 8680 3160 8740
rect 3220 8680 3240 8740
rect 3300 8680 3320 8740
rect 3380 8680 3680 8740
rect 3740 8680 3750 8740
rect 4101 8708 4105 8760
rect 4157 8708 4225 8760
rect 4277 8708 4585 8760
rect 4637 8708 4705 8760
rect 4757 8708 5065 8760
rect 5117 8708 6150 8760
rect 4101 8700 6150 8708
rect 6210 8700 6220 8760
rect 6140 8690 6220 8700
rect 2790 8660 3750 8680
rect 2790 8600 2800 8660
rect 2860 8600 3160 8660
rect 3220 8600 3240 8660
rect 3300 8600 3320 8660
rect 3380 8600 3680 8660
rect 3740 8600 3750 8660
rect 2790 8580 3750 8600
rect 230 8532 2540 8540
rect 230 8530 1526 8532
rect 230 8470 240 8530
rect 300 8480 1526 8530
rect 1578 8480 1684 8532
rect 1736 8480 2008 8532
rect 2060 8480 2162 8532
rect 2214 8480 2486 8532
rect 2538 8480 2540 8532
rect 2790 8520 2800 8580
rect 2860 8520 3160 8580
rect 3220 8520 3240 8580
rect 3300 8520 3320 8580
rect 3380 8520 3680 8580
rect 3740 8520 3750 8580
rect 2790 8510 3750 8520
rect 4000 8532 6310 8540
rect 300 8470 2540 8480
rect 4000 8480 4002 8532
rect 4054 8480 4326 8532
rect 4378 8480 4480 8532
rect 4532 8480 4804 8532
rect 4856 8480 4962 8532
rect 5014 8530 6310 8532
rect 5014 8480 6240 8530
rect 4000 8470 6240 8480
rect 6300 8470 6310 8530
rect 230 8460 310 8470
rect 6230 8460 6310 8470
rect 1590 8430 2630 8440
rect 1590 8370 1600 8430
rect 1660 8370 2080 8430
rect 2140 8370 2560 8430
rect 2620 8370 2630 8430
rect 1590 8360 2630 8370
rect 3910 8430 4950 8440
rect 3910 8370 3920 8430
rect 3980 8370 4400 8430
rect 4460 8370 4880 8430
rect 4940 8370 4950 8430
rect 3910 8360 4950 8370
rect 1350 8320 2390 8330
rect 1350 8260 1360 8320
rect 1420 8260 1840 8320
rect 1900 8260 2320 8320
rect 2380 8260 2390 8320
rect 1350 8250 2390 8260
rect 4150 8320 5190 8330
rect 4150 8260 4160 8320
rect 4220 8260 4640 8320
rect 4700 8260 5120 8320
rect 5180 8260 5190 8320
rect 4150 8250 5190 8260
rect 9790 8280 9870 8290
rect 9790 8220 9800 8280
rect 9860 8220 9870 8280
rect 3730 8210 6810 8220
rect 9790 8210 9870 8220
rect 3730 8150 3740 8210
rect 3800 8150 3920 8210
rect 3980 8150 4160 8210
rect 4220 8150 4400 8210
rect 4460 8150 4640 8210
rect 4700 8150 5120 8210
rect 5180 8150 5360 8210
rect 5420 8150 5780 8210
rect 5840 8150 6580 8210
rect 6640 8150 6660 8210
rect 6720 8150 6740 8210
rect 6800 8150 6810 8210
rect 3730 8130 6810 8150
rect 3730 8070 3740 8130
rect 3800 8070 3920 8130
rect 3980 8070 4160 8130
rect 4220 8070 4400 8130
rect 4460 8070 4640 8130
rect 4700 8070 5120 8130
rect 5180 8070 5360 8130
rect 5420 8070 5780 8130
rect 5840 8070 6580 8130
rect 6640 8070 6660 8130
rect 6720 8070 6740 8130
rect 6800 8070 6810 8130
rect 7830 8160 7930 8180
rect 7830 8100 7850 8160
rect 7910 8100 7930 8160
rect 7830 8080 7930 8100
rect 9810 8070 9850 8210
rect 610 8050 2810 8060
rect 610 7990 620 8050
rect 680 7990 700 8050
rect 760 7990 1120 8050
rect 1180 7990 1360 8050
rect 1420 7990 1840 8050
rect 1900 7990 2080 8050
rect 2140 7990 2560 8050
rect 2620 7990 2740 8050
rect 2800 7990 2810 8050
rect 610 7980 2810 7990
rect 3730 8050 6810 8070
rect 3730 7990 3740 8050
rect 3800 7990 3920 8050
rect 3980 7990 4160 8050
rect 4220 7990 4400 8050
rect 4460 7990 4640 8050
rect 4700 7990 5120 8050
rect 5180 7990 5360 8050
rect 5420 7990 5780 8050
rect 5840 7990 6580 8050
rect 6640 7990 6660 8050
rect 6720 7990 6740 8050
rect 6800 7990 6810 8050
rect 9790 8060 9870 8070
rect 9790 8000 9800 8060
rect 9860 8000 9870 8060
rect 9790 7990 9870 8000
rect 3730 7980 6810 7990
rect 870 7930 950 7940
rect 870 7870 880 7930
rect 940 7920 950 7930
rect 1590 7930 1670 7940
rect 1590 7920 1600 7930
rect 940 7880 1600 7920
rect 940 7870 950 7880
rect 870 7860 950 7870
rect 1590 7870 1600 7880
rect 1660 7920 1670 7930
rect 2310 7930 2390 7940
rect 2310 7920 2320 7930
rect 1660 7880 2320 7920
rect 1660 7870 1670 7880
rect 1590 7860 1670 7870
rect 2310 7870 2320 7880
rect 2380 7870 2390 7930
rect 2310 7860 2390 7870
rect 4150 7930 4230 7940
rect 4150 7870 4160 7930
rect 4220 7920 4230 7930
rect 4870 7930 4950 7940
rect 4870 7920 4880 7930
rect 4220 7880 4880 7920
rect 4220 7870 4230 7880
rect 4150 7860 4230 7870
rect 4870 7870 4880 7880
rect 4940 7920 4950 7930
rect 5590 7930 5670 7940
rect 5590 7920 5600 7930
rect 4940 7880 5600 7920
rect 4940 7870 4950 7880
rect 4870 7860 4950 7870
rect 5590 7870 5600 7880
rect 5660 7870 5670 7930
rect 5590 7860 5670 7870
rect 11750 7880 11860 7900
rect 11750 7810 11770 7880
rect 11840 7810 11860 7880
rect 11750 7790 11860 7810
rect 9570 7780 9650 7790
rect 8890 7720 8970 7730
rect 7550 7710 7630 7720
rect 7550 7650 7560 7710
rect 7620 7680 7630 7710
rect 8070 7700 8150 7710
rect 8070 7680 8080 7700
rect 7620 7650 8080 7680
rect 7550 7640 7630 7650
rect 8070 7640 8080 7650
rect 8140 7640 8150 7700
rect 1360 7600 1420 7630
rect 5120 7600 5180 7640
rect 8070 7630 8150 7640
rect 8890 7660 8900 7720
rect 8960 7660 8970 7720
rect 9570 7720 9580 7780
rect 9640 7720 9650 7780
rect 9570 7710 9650 7720
rect 8890 7650 8970 7660
rect 110 7590 3130 7600
rect 110 7530 120 7590
rect 180 7530 640 7590
rect 700 7530 1360 7590
rect 1420 7530 2080 7590
rect 2140 7530 2800 7590
rect 2860 7530 3060 7590
rect 3120 7530 3130 7590
rect 110 7520 3130 7530
rect 3410 7590 6540 7600
rect 3410 7530 3420 7590
rect 3480 7530 3680 7590
rect 3740 7530 4400 7590
rect 4460 7530 5120 7590
rect 5180 7530 5840 7590
rect 5900 7530 6470 7590
rect 6530 7530 6540 7590
rect 8430 7560 8510 7570
rect 3410 7520 6540 7530
rect 7440 7540 7520 7550
rect 510 7480 7300 7490
rect 510 7420 520 7480
rect 580 7420 760 7480
rect 820 7420 1000 7480
rect 1060 7420 1240 7480
rect 1300 7420 1480 7480
rect 1540 7420 1720 7480
rect 1780 7420 1960 7480
rect 2020 7420 2200 7480
rect 2260 7420 2440 7480
rect 2500 7420 2680 7480
rect 2740 7420 2920 7480
rect 2980 7420 3560 7480
rect 3620 7420 3800 7480
rect 3860 7420 4040 7480
rect 4100 7420 4280 7480
rect 4340 7420 4520 7480
rect 4580 7420 4760 7480
rect 4820 7420 5000 7480
rect 5060 7420 5240 7480
rect 5300 7420 5480 7480
rect 5540 7420 5720 7480
rect 5780 7420 5960 7480
rect 6020 7450 7300 7480
rect 7440 7480 7450 7540
rect 7510 7520 7520 7540
rect 8070 7540 8150 7550
rect 8070 7520 8080 7540
rect 7510 7490 8080 7520
rect 7510 7480 7520 7490
rect 7440 7470 7520 7480
rect 8070 7480 8080 7490
rect 8140 7480 8150 7540
rect 8430 7500 8440 7560
rect 8500 7500 8510 7560
rect 8430 7490 8510 7500
rect 8070 7470 8150 7480
rect 8450 7460 8480 7490
rect 8890 7460 8920 7650
rect 9590 7560 9620 7710
rect 14230 7610 14310 7620
rect 9570 7550 9650 7560
rect 9570 7490 9580 7550
rect 9640 7490 9650 7550
rect 14230 7550 14240 7610
rect 14300 7550 14310 7610
rect 14230 7540 14310 7550
rect 9570 7480 9650 7490
rect 6020 7420 7220 7450
rect 510 7400 7220 7420
rect 510 7340 520 7400
rect 580 7340 760 7400
rect 820 7340 1000 7400
rect 1060 7340 1240 7400
rect 1300 7340 1480 7400
rect 1540 7340 1720 7400
rect 1780 7340 1960 7400
rect 2020 7340 2200 7400
rect 2260 7340 2440 7400
rect 2500 7340 2680 7400
rect 2740 7340 2920 7400
rect 2980 7340 3560 7400
rect 3620 7340 3800 7400
rect 3860 7340 4040 7400
rect 4100 7340 4280 7400
rect 4340 7340 4520 7400
rect 4580 7340 4760 7400
rect 4820 7340 5000 7400
rect 5060 7340 5240 7400
rect 5300 7340 5480 7400
rect 5540 7340 5720 7400
rect 5780 7340 5960 7400
rect 6020 7390 7220 7400
rect 7280 7390 7300 7450
rect 6020 7350 7300 7390
rect 8430 7450 8510 7460
rect 8430 7390 8440 7450
rect 8500 7390 8510 7450
rect 8430 7380 8510 7390
rect 8870 7450 8950 7460
rect 8870 7390 8880 7450
rect 8940 7390 8950 7450
rect 8870 7380 8950 7390
rect 11750 7380 11860 7400
rect 6020 7340 7220 7350
rect 510 7320 7220 7340
rect 510 7260 520 7320
rect 580 7260 760 7320
rect 820 7260 1000 7320
rect 1060 7260 1240 7320
rect 1300 7260 1480 7320
rect 1540 7260 1720 7320
rect 1780 7260 1960 7320
rect 2020 7260 2200 7320
rect 2260 7260 2440 7320
rect 2500 7260 2680 7320
rect 2740 7260 2920 7320
rect 2980 7260 3560 7320
rect 3620 7260 3800 7320
rect 3860 7260 4040 7320
rect 4100 7260 4280 7320
rect 4340 7260 4520 7320
rect 4580 7260 4760 7320
rect 4820 7260 5000 7320
rect 5060 7260 5240 7320
rect 5300 7260 5480 7320
rect 5540 7260 5720 7320
rect 5780 7260 5960 7320
rect 6020 7290 7220 7320
rect 7280 7290 7300 7350
rect 11750 7310 11770 7380
rect 11840 7310 11860 7380
rect 11750 7290 11860 7310
rect 6020 7260 7300 7290
rect 510 7250 7300 7260
rect 230 7210 4750 7220
rect 230 7150 240 7210
rect 300 7150 1800 7210
rect 1860 7150 3240 7210
rect 3300 7150 4680 7210
rect 4740 7150 4750 7210
rect 230 7140 4750 7150
rect 0 7100 5780 7110
rect 0 7040 10 7100
rect 70 7040 2160 7100
rect 2220 7040 4320 7100
rect 4380 7040 5710 7100
rect 5770 7040 5780 7100
rect 0 7030 5780 7040
rect 8750 7070 8830 7080
rect 8750 7010 8760 7070
rect 8820 7010 8830 7070
rect 8750 7000 8830 7010
rect 2510 6990 6310 7000
rect 2510 6930 2520 6990
rect 2580 6930 3960 6990
rect 4020 6930 5240 6990
rect 5300 6930 6240 6990
rect 6300 6930 6310 6990
rect 2510 6920 6310 6930
rect 7830 6970 7930 6990
rect 7830 6910 7850 6970
rect 7910 6910 7930 6970
rect 7830 6890 7930 6910
rect 2870 6880 6220 6890
rect 2870 6820 2880 6880
rect 2940 6820 3600 6880
rect 3660 6820 6150 6880
rect 6210 6820 6220 6880
rect 8770 6860 8810 7000
rect 2870 6810 6220 6820
rect 8750 6850 8830 6860
rect 8750 6790 8760 6850
rect 8820 6790 8830 6850
rect 8750 6780 8830 6790
rect 1890 6770 4650 6780
rect 1950 6710 2070 6770
rect 2130 6710 2250 6770
rect 2310 6710 2430 6770
rect 2490 6710 2610 6770
rect 2670 6710 2790 6770
rect 2850 6710 2970 6770
rect 3030 6710 3150 6770
rect 3210 6710 3330 6770
rect 3390 6710 3420 6770
rect 3480 6710 3510 6770
rect 3570 6710 3690 6770
rect 3750 6710 3870 6770
rect 3930 6710 4050 6770
rect 4110 6710 4230 6770
rect 4290 6710 4410 6770
rect 4470 6710 4590 6770
rect 1890 6700 4650 6710
rect 5580 6570 5900 6580
rect 5580 6510 5590 6570
rect 5650 6510 5830 6570
rect 5890 6510 5900 6570
rect 5580 6500 5900 6510
rect 5230 6230 5310 6240
rect 5230 6170 5240 6230
rect 5300 6220 5310 6230
rect 5700 6230 5780 6240
rect 5700 6220 5710 6230
rect 5300 6180 5710 6220
rect 5300 6170 5310 6180
rect 5230 6160 5310 6170
rect 5700 6170 5710 6180
rect 5770 6170 5780 6230
rect 5700 6160 5780 6170
rect 1610 6030 7300 6040
rect 1610 5970 1620 6030
rect 1680 5970 1980 6030
rect 2040 5970 2340 6030
rect 2400 5970 2700 6030
rect 2760 5970 3060 6030
rect 3120 5970 3420 6030
rect 3480 5970 3780 6030
rect 3840 5970 4140 6030
rect 4200 5970 4500 6030
rect 4560 5970 4860 6030
rect 4920 5970 5490 6030
rect 5550 5970 5930 6030
rect 5990 6000 7300 6030
rect 5990 5970 7220 6000
rect 1610 5950 7220 5970
rect 1610 5890 1620 5950
rect 1680 5890 1980 5950
rect 2040 5890 2340 5950
rect 2400 5890 2700 5950
rect 2760 5890 3060 5950
rect 3120 5890 3420 5950
rect 3480 5890 3780 5950
rect 3840 5890 4140 5950
rect 4200 5890 4500 5950
rect 4560 5890 4860 5950
rect 4920 5890 5490 5950
rect 5550 5890 5930 5950
rect 5990 5940 7220 5950
rect 7280 5940 7300 6000
rect 5990 5900 7300 5940
rect 5990 5890 7220 5900
rect 1610 5870 7220 5890
rect 1610 5810 1620 5870
rect 1680 5810 1980 5870
rect 2040 5810 2340 5870
rect 2400 5810 2700 5870
rect 2760 5810 3060 5870
rect 3120 5810 3420 5870
rect 3480 5810 3780 5870
rect 3840 5810 4140 5870
rect 4200 5810 4500 5870
rect 4560 5810 4860 5870
rect 4920 5810 5490 5870
rect 5550 5810 5930 5870
rect 5990 5840 7220 5870
rect 7280 5840 7300 5900
rect 5990 5810 7300 5840
rect 1610 5800 7300 5810
rect 110 5710 120 5770
rect 180 5760 4744 5770
rect 180 5710 1798 5760
rect 110 5708 1798 5710
rect 1850 5708 1908 5760
rect 1960 5708 2018 5760
rect 2070 5708 2128 5760
rect 2180 5708 2238 5760
rect 2290 5708 2348 5760
rect 2400 5708 2458 5760
rect 2510 5708 2568 5760
rect 2620 5708 2678 5760
rect 2730 5708 2788 5760
rect 2840 5708 3698 5760
rect 3750 5708 3808 5760
rect 3860 5708 3918 5760
rect 3970 5708 4028 5760
rect 4080 5708 4138 5760
rect 4190 5708 4248 5760
rect 4300 5708 4358 5760
rect 4410 5708 4468 5760
rect 4520 5708 4578 5760
rect 4630 5708 4688 5760
rect 4740 5708 4744 5760
rect 110 5700 4744 5708
rect 7200 5440 7300 5450
rect 1620 5430 7300 5440
rect 1620 5370 1630 5430
rect 1690 5370 1850 5430
rect 1910 5370 2070 5430
rect 2130 5370 2290 5430
rect 2350 5370 2510 5430
rect 2570 5370 2730 5430
rect 2790 5370 2950 5430
rect 3010 5370 3530 5430
rect 3590 5370 3750 5430
rect 3810 5370 3970 5430
rect 4030 5370 4190 5430
rect 4250 5370 4410 5430
rect 4470 5370 4630 5430
rect 4690 5370 4850 5430
rect 4910 5370 7220 5430
rect 7280 5370 7300 5430
rect 1620 5360 7300 5370
rect 11750 5440 11850 5460
rect 11750 5380 11770 5440
rect 11830 5380 11850 5440
rect 11750 5360 11850 5380
rect 7200 5350 7300 5360
rect 340 5320 2910 5330
rect 340 5260 350 5320
rect 410 5260 1740 5320
rect 1800 5260 1960 5320
rect 2020 5260 2180 5320
rect 2240 5260 2400 5320
rect 2460 5260 2620 5320
rect 2680 5260 2840 5320
rect 2900 5260 2910 5320
rect 340 5250 2910 5260
rect 3630 5320 4810 5330
rect 3630 5260 3640 5320
rect 3700 5260 3860 5320
rect 3920 5260 4080 5320
rect 4140 5260 4300 5320
rect 4360 5260 4520 5320
rect 4580 5260 4740 5320
rect 4800 5260 4810 5320
rect 3630 5250 4810 5260
rect 7660 5300 7740 5310
rect 14250 5300 14280 7540
rect 7660 5240 7670 5300
rect 7730 5280 7740 5300
rect 14230 5290 14310 5300
rect 14230 5280 14240 5290
rect 7730 5250 14240 5280
rect 7730 5240 7740 5250
rect 7660 5230 7740 5240
rect 14230 5230 14240 5250
rect 14300 5230 14310 5290
rect 14230 5220 14310 5230
rect 1150 5210 4810 5220
rect 1150 5150 1160 5210
rect 1220 5150 1240 5210
rect 1300 5150 1320 5210
rect 1380 5150 3640 5210
rect 3700 5150 3860 5210
rect 3920 5150 4080 5210
rect 4140 5150 4300 5210
rect 4360 5150 4520 5210
rect 4580 5150 4740 5210
rect 4800 5150 4810 5210
rect 1150 5130 4810 5150
rect 1150 5070 1160 5130
rect 1220 5070 1240 5130
rect 1300 5070 1320 5130
rect 1380 5070 3640 5130
rect 3700 5070 3860 5130
rect 3920 5070 4080 5130
rect 4140 5070 4300 5130
rect 4360 5070 4520 5130
rect 4580 5070 4740 5130
rect 4800 5070 4810 5130
rect 7440 5190 7520 5200
rect 7440 5130 7450 5190
rect 7510 5180 7520 5190
rect 13180 5190 13260 5200
rect 13180 5180 13190 5190
rect 7510 5140 13190 5180
rect 7510 5130 7520 5140
rect 7440 5120 7520 5130
rect 13180 5130 13190 5140
rect 13250 5130 13260 5190
rect 13180 5120 13260 5130
rect 11590 5090 11700 5110
rect 1150 5050 4810 5070
rect 1150 4990 1160 5050
rect 1220 4990 1240 5050
rect 1300 4990 1320 5050
rect 1380 4990 3640 5050
rect 3700 4990 3860 5050
rect 3920 4990 4080 5050
rect 4140 4990 4300 5050
rect 4360 4990 4520 5050
rect 4580 4990 4740 5050
rect 4800 4990 4810 5050
rect 7350 5080 7430 5090
rect 7350 5020 7360 5080
rect 7420 5070 7430 5080
rect 11590 5070 11610 5090
rect 7420 5040 11610 5070
rect 7420 5020 7430 5040
rect 7350 5010 7430 5020
rect 11590 5020 11610 5040
rect 11680 5020 11700 5090
rect 11590 5000 11700 5020
rect 1150 4980 4810 4990
rect 1720 4930 1820 4950
rect 1720 4870 1740 4930
rect 1800 4870 1820 4930
rect 1720 4850 1820 4870
rect 7040 4940 7140 4960
rect 7040 4880 7060 4940
rect 7120 4880 7140 4940
rect 7040 4860 7140 4880
rect 6340 4830 6420 4840
rect 6340 4770 6350 4830
rect 6410 4820 6420 4830
rect 7440 4830 7520 4840
rect 7440 4820 7450 4830
rect 6410 4780 7450 4820
rect 6410 4770 6420 4780
rect 6340 4760 6420 4770
rect 7440 4770 7450 4780
rect 7510 4770 7520 4830
rect 7440 4760 7520 4770
rect 6640 4700 6720 4710
rect 6640 4640 6650 4700
rect 6710 4690 6720 4700
rect 7350 4700 7430 4710
rect 7350 4690 7360 4700
rect 6710 4650 7360 4690
rect 6710 4640 6720 4650
rect 6640 4630 6720 4640
rect 7350 4640 7360 4650
rect 7420 4640 7430 4700
rect 7350 4630 7430 4640
rect 7750 4560 7850 4580
rect 7750 4500 7770 4560
rect 7830 4500 7850 4560
rect 550 4480 2010 4490
rect 550 4420 1940 4480
rect 2000 4420 2010 4480
rect 550 4410 2010 4420
rect 3840 4480 3920 4490
rect 7750 4480 7850 4500
rect 3840 4420 3850 4480
rect 3910 4420 3920 4480
rect 3840 4410 3920 4420
rect 1900 3760 2000 3780
rect 1900 3700 1920 3760
rect 1980 3700 2000 3760
rect 1900 3680 2000 3700
rect 3880 3090 3920 4410
rect 5010 4440 5090 4450
rect 5010 4380 5020 4440
rect 5080 4380 5090 4440
rect 5010 4370 5090 4380
rect 6640 4410 6720 4420
rect 4140 3870 4220 3880
rect 4140 3810 4150 3870
rect 4210 3810 4220 3870
rect 4140 3800 4220 3810
rect 4160 3660 4200 3800
rect 4120 3650 4200 3660
rect 4120 3590 4130 3650
rect 4190 3590 4200 3650
rect 4120 3580 4200 3590
rect 5020 3090 5060 4370
rect 6640 4350 6650 4410
rect 6710 4350 6720 4410
rect 6640 4340 6720 4350
rect 6880 4410 6960 4420
rect 6880 4350 6890 4410
rect 6950 4400 6960 4410
rect 7350 4410 7430 4420
rect 7350 4400 7360 4410
rect 6950 4360 7360 4400
rect 6950 4350 6960 4360
rect 6880 4340 6960 4350
rect 7350 4350 7360 4360
rect 7420 4350 7430 4410
rect 7350 4340 7430 4350
rect 11350 3910 11460 3930
rect 7440 3890 7520 3900
rect 7440 3830 7450 3890
rect 7510 3880 7520 3890
rect 7660 3890 7740 3900
rect 7660 3880 7670 3890
rect 7510 3840 7670 3880
rect 7510 3830 7520 3840
rect 7440 3820 7520 3830
rect 7660 3830 7670 3840
rect 7730 3880 7740 3890
rect 8460 3890 8540 3900
rect 8460 3880 8470 3890
rect 7730 3840 8470 3880
rect 7730 3830 7740 3840
rect 7660 3820 7740 3830
rect 8460 3830 8470 3840
rect 8530 3830 8540 3890
rect 8460 3820 8540 3830
rect 11350 3840 11370 3910
rect 11440 3840 11460 3910
rect 11350 3820 11460 3840
rect 7550 3800 7630 3810
rect 7200 3770 7300 3790
rect 7200 3710 7220 3770
rect 7280 3710 7300 3770
rect 7550 3740 7560 3800
rect 7620 3790 7630 3800
rect 8590 3800 8670 3810
rect 8590 3790 8600 3800
rect 7620 3750 8600 3790
rect 7620 3740 7630 3750
rect 7200 3690 7300 3710
rect 7350 3730 7430 3740
rect 7550 3730 7630 3740
rect 8590 3740 8600 3750
rect 8660 3740 8670 3800
rect 8590 3730 8670 3740
rect 7350 3670 7360 3730
rect 7420 3700 7430 3730
rect 11180 3720 11260 3730
rect 9980 3710 10060 3720
rect 9980 3700 9990 3710
rect 7420 3670 9990 3700
rect 7350 3660 9990 3670
rect 3860 3080 3940 3090
rect 1610 3040 1690 3050
rect 1610 2980 1620 3040
rect 1680 2980 1690 3040
rect 3860 3020 3870 3080
rect 3930 3020 3940 3080
rect 3860 3010 3940 3020
rect 4940 3080 5060 3090
rect 4940 3020 4950 3080
rect 5010 3020 5060 3080
rect 4940 3010 5060 3020
rect 5710 3650 5790 3660
rect 5710 3590 5720 3650
rect 5780 3590 5790 3650
rect 5710 3580 5790 3590
rect 5830 3650 5910 3660
rect 5830 3590 5840 3650
rect 5900 3590 5910 3650
rect 9980 3650 9990 3660
rect 10050 3650 10060 3710
rect 11180 3660 11190 3720
rect 11250 3710 11260 3720
rect 13180 3720 13260 3730
rect 13180 3710 13190 3720
rect 11250 3670 13190 3710
rect 11250 3660 11260 3670
rect 11180 3650 11260 3660
rect 13180 3660 13190 3670
rect 13250 3660 13260 3720
rect 13180 3650 13260 3660
rect 9980 3640 10060 3650
rect 5830 3580 5910 3590
rect 6640 3620 8470 3630
rect 1610 2970 1690 2980
rect 5710 2700 5750 3580
rect 5830 2700 5870 3580
rect 6640 3560 6650 3620
rect 6710 3560 7280 3620
rect 7340 3560 7360 3620
rect 7420 3560 7440 3620
rect 7500 3560 8400 3620
rect 8460 3560 8470 3620
rect 6640 3550 8470 3560
rect 10420 3510 10500 3520
rect 7750 3500 7830 3510
rect 10420 3500 10430 3510
rect 7750 3440 7760 3500
rect 7820 3460 10430 3500
rect 7820 3440 7830 3460
rect 10420 3450 10430 3460
rect 10490 3450 10500 3510
rect 10420 3440 10500 3450
rect 11350 3500 11460 3520
rect 7750 3430 7830 3440
rect 11350 3430 11370 3500
rect 11440 3430 11460 3500
rect 11350 3410 11460 3430
rect 6890 3080 6970 3090
rect 6890 3020 6900 3080
rect 6960 3070 6970 3080
rect 7750 3080 7830 3090
rect 7750 3070 7760 3080
rect 6960 3030 7760 3070
rect 6960 3020 6970 3030
rect 6890 3010 6970 3020
rect 7750 3020 7760 3030
rect 7820 3020 7830 3080
rect 7750 3010 7830 3020
rect 7750 2860 7850 2880
rect 7750 2800 7770 2860
rect 7830 2800 7850 2860
rect 7750 2780 7850 2800
rect 17090 2730 17200 2750
rect 11700 2710 11810 2730
rect 5670 2690 5750 2700
rect 5670 2630 5680 2690
rect 5740 2630 5750 2690
rect 5670 2620 5750 2630
rect 5790 2690 5870 2700
rect 5790 2630 5800 2690
rect 5860 2630 5870 2690
rect 5790 2620 5870 2630
rect 6430 2690 6510 2700
rect 11700 2690 11720 2710
rect 6430 2630 6440 2690
rect 6500 2660 11720 2690
rect 6500 2630 6510 2660
rect 6430 2620 6510 2630
rect 11700 2640 11720 2660
rect 11790 2640 11810 2710
rect 17090 2660 17110 2730
rect 17180 2660 17200 2730
rect 17090 2640 17200 2660
rect 17590 2730 17700 2750
rect 17590 2660 17610 2730
rect 17680 2660 17700 2730
rect 17590 2640 17700 2660
rect 11700 2620 11810 2640
rect 1720 2590 1820 2610
rect 1720 2530 1740 2590
rect 1800 2530 1820 2590
rect 1720 2510 1820 2530
rect 7040 2580 7140 2600
rect 7040 2520 7060 2580
rect 7120 2520 7140 2580
rect 14410 2520 14510 2540
rect 7040 2500 7140 2520
rect 13180 2510 13260 2520
rect 1150 2460 7510 2470
rect 1150 2400 1160 2460
rect 1220 2400 1240 2460
rect 1300 2400 1320 2460
rect 1380 2400 7280 2460
rect 7340 2400 7360 2460
rect 7420 2400 7440 2460
rect 7500 2400 7510 2460
rect 13180 2450 13190 2510
rect 13250 2500 13260 2510
rect 14300 2510 14430 2520
rect 14300 2500 14310 2510
rect 13250 2460 14310 2500
rect 13250 2450 13260 2460
rect 13180 2440 13260 2450
rect 14300 2450 14310 2460
rect 14370 2460 14430 2510
rect 14490 2460 14510 2520
rect 14370 2450 14510 2460
rect 14300 2440 14510 2450
rect 31480 2520 31580 2540
rect 31480 2460 31500 2520
rect 31560 2460 31580 2520
rect 31480 2440 31580 2460
rect 1150 2380 7510 2400
rect 1150 2320 1160 2380
rect 1220 2320 1240 2380
rect 1300 2320 1320 2380
rect 1380 2320 7280 2380
rect 7340 2320 7360 2380
rect 7420 2320 7440 2380
rect 7500 2320 7510 2380
rect 1150 2300 7510 2320
rect 1150 2240 1160 2300
rect 1220 2240 1240 2300
rect 1300 2240 1320 2300
rect 1380 2240 7280 2300
rect 7340 2240 7360 2300
rect 7420 2240 7440 2300
rect 7500 2240 7510 2300
rect 1150 2230 7510 2240
rect 7040 2180 7140 2200
rect 7040 2120 7060 2180
rect 7120 2120 7140 2180
rect 7040 2100 7140 2120
rect 12170 2160 12270 2180
rect 12170 2100 12190 2160
rect 12250 2100 12270 2160
rect 12170 2080 12270 2100
rect 14320 1830 14350 2440
rect 14300 1820 14380 1830
rect 14300 1760 14310 1820
rect 14370 1760 14380 1820
rect 14300 1750 14380 1760
rect 12170 1660 12270 1680
rect 12170 1600 12190 1660
rect 12250 1600 12270 1660
rect 12170 1580 12270 1600
rect 1610 1270 1690 1280
rect 1610 1210 1620 1270
rect 1680 1210 1690 1270
rect 1610 1200 1690 1210
rect 1620 880 1720 900
rect 1620 820 1640 880
rect 1700 820 1720 880
rect 1620 800 1720 820
rect 12170 860 12270 880
rect 12170 800 12190 860
rect 12250 800 12270 860
rect 12170 780 12270 800
rect 12170 80 12270 100
rect 12170 20 12190 80
rect 12250 20 12270 80
rect 12170 0 12270 20
<< via2 >>
rect 7290 14800 7350 14860
rect 6970 14100 7030 14160
rect 7220 13400 7280 13460
rect 7090 12700 7150 12760
rect 7290 12000 7350 12060
rect 7090 11300 7150 11360
rect 7060 10160 7120 10220
rect 7060 9850 7120 9910
rect 7060 9750 7120 9810
rect 11770 9750 11830 9810
rect 7220 9050 7280 9110
rect 7220 8950 7280 9010
rect 7850 8100 7910 8160
rect 11770 7810 11840 7880
rect 7220 7390 7280 7450
rect 7220 7290 7280 7350
rect 11770 7310 11840 7380
rect 7850 6910 7910 6970
rect 7220 5940 7280 6000
rect 7220 5840 7280 5900
rect 7220 5370 7280 5430
rect 11770 5380 11830 5440
rect 11610 5020 11680 5090
rect 1740 4870 1800 4930
rect 7060 4880 7120 4940
rect 7770 4500 7830 4560
rect 1920 3700 1980 3760
rect 11370 3840 11440 3910
rect 7220 3710 7280 3770
rect 11370 3430 11440 3500
rect 7770 2800 7830 2860
rect 11720 2640 11790 2710
rect 17110 2660 17180 2730
rect 17610 2660 17680 2730
rect 1740 2530 1800 2590
rect 7060 2520 7120 2580
rect 14430 2460 14490 2520
rect 31500 2460 31560 2520
rect 7060 2120 7120 2180
rect 12190 2100 12250 2160
rect 12190 1600 12250 1660
rect 1640 820 1700 880
rect 12190 800 12250 860
rect 12190 20 12250 80
<< metal3 >>
rect 7410 14880 7870 15050
rect 8110 14880 8570 15050
rect 8810 14880 9270 15050
rect 9510 14880 9970 15050
rect 10210 14880 10670 15050
rect 10910 14880 11370 15050
rect 11610 14880 12070 15050
rect 12310 14880 12770 15050
rect 13010 14880 13470 15050
rect 13710 14880 14170 15050
rect 7410 14870 14170 14880
rect 7280 14860 14170 14870
rect 7280 14800 7290 14860
rect 7350 14800 14170 14860
rect 7280 14790 14170 14800
rect 7410 14780 14170 14790
rect 7410 14590 7870 14780
rect 8110 14590 8570 14780
rect 8810 14590 9270 14780
rect 9510 14590 9970 14780
rect 10210 14590 10670 14780
rect 10910 14590 11370 14780
rect 11610 14590 12070 14780
rect 12310 14590 12770 14780
rect 13010 14590 13470 14780
rect 13710 14590 14170 14780
rect 13890 14350 13990 14590
rect 7410 14180 7870 14350
rect 8110 14180 8570 14350
rect 8810 14180 9270 14350
rect 9510 14180 9970 14350
rect 10210 14180 10670 14350
rect 10910 14180 11370 14350
rect 11610 14180 12070 14350
rect 12310 14180 12770 14350
rect 13010 14180 13470 14350
rect 13710 14180 14170 14350
rect 6950 14170 7050 14180
rect 6950 14090 6960 14170
rect 7040 14090 7050 14170
rect 6950 14080 7050 14090
rect 7410 14080 14170 14180
rect 7410 13890 7870 14080
rect 8110 13890 8570 14080
rect 8810 13890 9270 14080
rect 9510 13890 9970 14080
rect 10210 13890 10670 14080
rect 10910 13890 11370 14080
rect 11610 13890 12070 14080
rect 12310 13890 12770 14080
rect 13010 13890 13470 14080
rect 13710 13890 14170 14080
rect 7410 13480 7870 13650
rect 8110 13480 8570 13650
rect 8810 13480 9270 13650
rect 9510 13480 9970 13650
rect 10210 13480 10670 13650
rect 10910 13480 11370 13650
rect 11610 13480 12070 13650
rect 12310 13480 12770 13650
rect 13010 13480 13470 13650
rect 13710 13480 14170 13650
rect 7410 13470 14170 13480
rect 7210 13460 14170 13470
rect 7210 13400 7220 13460
rect 7280 13400 14170 13460
rect 7210 13390 14170 13400
rect 7410 13380 14170 13390
rect 7410 13190 7870 13380
rect 8110 13190 8570 13380
rect 8810 13190 9270 13380
rect 9510 13190 9970 13380
rect 10210 13190 10670 13380
rect 10910 13190 11370 13380
rect 11610 13190 12070 13380
rect 12310 13190 12770 13380
rect 13010 13190 13470 13380
rect 13710 13190 14170 13380
rect 13890 12950 13990 13190
rect 7410 12780 7870 12950
rect 8110 12780 8570 12950
rect 8810 12780 9270 12950
rect 9510 12780 9970 12950
rect 10210 12780 10670 12950
rect 10910 12780 11370 12950
rect 11610 12780 12070 12950
rect 12310 12780 12770 12950
rect 13010 12780 13470 12950
rect 13710 12780 14170 12950
rect 7070 12770 7170 12780
rect 7070 12690 7080 12770
rect 7160 12690 7170 12770
rect 7070 12680 7170 12690
rect 7410 12680 14170 12780
rect 7410 12490 7870 12680
rect 8110 12490 8570 12680
rect 8810 12490 9270 12680
rect 9510 12490 9970 12680
rect 10210 12490 10670 12680
rect 10910 12490 11370 12680
rect 11610 12490 12070 12680
rect 12310 12490 12770 12680
rect 13010 12490 13470 12680
rect 13710 12490 14170 12680
rect 7410 12080 7870 12250
rect 8110 12080 8570 12250
rect 8810 12080 9270 12250
rect 9510 12080 9970 12250
rect 10210 12080 10670 12250
rect 10910 12080 11370 12250
rect 11610 12080 12070 12250
rect 12310 12080 12770 12250
rect 13010 12080 13470 12250
rect 13710 12080 14170 12250
rect 7410 12070 14170 12080
rect 7280 12060 14170 12070
rect 7280 12000 7290 12060
rect 7350 12000 14170 12060
rect 7280 11990 14170 12000
rect 7410 11980 14170 11990
rect 7410 11790 7870 11980
rect 8110 11790 8570 11980
rect 8810 11790 9270 11980
rect 9510 11790 9970 11980
rect 10210 11790 10670 11980
rect 10910 11790 11370 11980
rect 11610 11790 12070 11980
rect 12310 11790 12770 11980
rect 13010 11790 13470 11980
rect 13710 11790 14170 11980
rect 13890 11550 13990 11790
rect 7410 11380 7870 11550
rect 8110 11380 8570 11550
rect 8810 11380 9270 11550
rect 9510 11380 9970 11550
rect 10210 11380 10670 11550
rect 10910 11380 11370 11550
rect 11610 11380 12070 11550
rect 12310 11380 12770 11550
rect 13010 11380 13470 11550
rect 13710 11380 14170 11550
rect 7070 11370 7170 11380
rect 7070 11290 7080 11370
rect 7160 11290 7170 11370
rect 7070 11280 7170 11290
rect 7410 11280 14170 11380
rect 7410 11090 7870 11280
rect 8110 11090 8570 11280
rect 8810 11090 9270 11280
rect 9510 11090 9970 11280
rect 10210 11090 10670 11280
rect 10910 11090 11370 11280
rect 11610 11090 12070 11280
rect 12310 11090 12770 11280
rect 13010 11090 13470 11280
rect 13710 11090 14170 11280
rect 7040 10220 7140 10270
rect 7040 10160 7060 10220
rect 7120 10160 7140 10220
rect 7040 9910 7140 10160
rect 7040 9850 7060 9910
rect 7120 9850 7140 9910
rect 7040 9810 7140 9850
rect 7040 9750 7060 9810
rect 7120 9750 7140 9810
rect 7040 8170 7140 9750
rect 11750 9820 11850 9830
rect 11750 9810 14160 9820
rect 11750 9750 11770 9810
rect 11830 9750 14160 9810
rect 11750 9730 14160 9750
rect 7040 8090 7050 8170
rect 7130 8090 7140 8170
rect 1720 4940 1820 4950
rect 1720 4860 1730 4940
rect 1810 4860 1820 4940
rect 1720 4850 1820 4860
rect 7040 4940 7140 8090
rect 7040 4880 7060 4940
rect 7120 4880 7140 4940
rect 1420 3770 2000 3780
rect 1420 3690 1430 3770
rect 1510 3760 2000 3770
rect 1510 3700 1920 3760
rect 1980 3700 2000 3760
rect 1510 3690 2000 3700
rect 1420 3680 2000 3690
rect 7040 2870 7140 4880
rect 7200 9110 7300 9150
rect 7200 9050 7220 9110
rect 7280 9050 7300 9110
rect 7200 9010 7300 9050
rect 7200 8950 7220 9010
rect 7280 8950 7300 9010
rect 7200 7450 7300 8950
rect 7830 8170 7930 8180
rect 7830 8090 7840 8170
rect 7920 8090 7930 8170
rect 7830 8080 7930 8090
rect 11750 7880 11860 7900
rect 11750 7810 11770 7880
rect 11840 7810 11860 7880
rect 11750 7790 11860 7810
rect 12100 7760 14160 9730
rect 7200 7390 7220 7450
rect 7280 7390 7300 7450
rect 7200 7350 7300 7390
rect 7200 7290 7220 7350
rect 7280 7290 7300 7350
rect 11750 7380 11860 7400
rect 11750 7310 11770 7380
rect 11840 7310 11860 7380
rect 11750 7290 11860 7310
rect 7200 6980 7300 7290
rect 7200 6900 7210 6980
rect 7290 6900 7300 6980
rect 7200 6000 7300 6900
rect 7830 6980 7930 6990
rect 7830 6900 7840 6980
rect 7920 6900 7930 6980
rect 7830 6890 7930 6900
rect 7200 5940 7220 6000
rect 7280 5940 7300 6000
rect 7200 5900 7300 5940
rect 7200 5840 7220 5900
rect 7280 5840 7300 5900
rect 7200 5430 7300 5840
rect 12100 5460 14160 7430
rect 7200 5370 7220 5430
rect 7280 5370 7300 5430
rect 7200 4570 7300 5370
rect 11750 5440 14160 5460
rect 11750 5380 11770 5440
rect 11830 5380 14160 5440
rect 11750 5370 14160 5380
rect 11750 5360 11850 5370
rect 11590 5090 12800 5110
rect 11590 5020 11610 5090
rect 11680 5020 12800 5090
rect 11590 5000 12800 5020
rect 7200 4490 7210 4570
rect 7290 4490 7300 4570
rect 7200 3770 7300 4490
rect 7750 4570 7850 4580
rect 7750 4490 7760 4570
rect 7840 4490 7850 4570
rect 7750 4480 7850 4490
rect 11350 3910 11460 3930
rect 11350 3840 11370 3910
rect 11440 3840 11460 3910
rect 11350 3820 11460 3840
rect 11700 3790 12800 5000
rect 7200 3710 7220 3770
rect 7280 3710 7300 3770
rect 7200 3690 7300 3710
rect 11350 3500 11460 3520
rect 11350 3430 11370 3500
rect 11440 3430 11460 3500
rect 11350 3410 11460 3430
rect 7040 2790 7050 2870
rect 7130 2790 7140 2870
rect 1720 2600 1820 2610
rect 1720 2520 1730 2600
rect 1810 2520 1820 2600
rect 1720 2510 1820 2520
rect 7040 2580 7140 2790
rect 7750 2870 7850 2880
rect 7750 2790 7760 2870
rect 7840 2790 7850 2870
rect 7750 2780 7850 2790
rect 11700 2730 12300 3550
rect 14410 2990 17230 15050
rect 17560 2990 31580 15050
rect 11700 2710 11810 2730
rect 11700 2640 11720 2710
rect 11790 2640 11810 2710
rect 11700 2620 11810 2640
rect 7040 2520 7060 2580
rect 7120 2520 7140 2580
rect 7040 2180 7140 2520
rect 14410 2520 14510 2990
rect 17090 2730 17200 2750
rect 17090 2660 17110 2730
rect 17180 2660 17200 2730
rect 17090 2640 17200 2660
rect 17590 2730 17700 2750
rect 17590 2660 17610 2730
rect 17680 2660 17700 2730
rect 17590 2640 17700 2660
rect 14410 2460 14430 2520
rect 14490 2460 14510 2520
rect 14410 2440 14510 2460
rect 31480 2520 31580 2990
rect 31480 2460 31500 2520
rect 31560 2460 31580 2520
rect 31480 2440 31580 2460
rect 7040 2120 7060 2180
rect 7120 2120 7140 2180
rect 7040 2100 7140 2120
rect 12170 2170 12270 2180
rect 12170 2090 12180 2170
rect 12260 2090 12270 2170
rect 12170 2080 12270 2090
rect 12170 1670 12270 1680
rect 12170 1590 12180 1670
rect 12260 1590 12270 1670
rect 12170 1580 12270 1590
rect 1420 890 1720 900
rect 1420 810 1430 890
rect 1510 880 1720 890
rect 1510 820 1640 880
rect 1700 820 1720 880
rect 1510 810 1720 820
rect 1420 800 1720 810
rect 12170 870 12270 880
rect 12170 790 12180 870
rect 12260 790 12270 870
rect 12170 780 12270 790
rect 12170 90 12270 100
rect 12170 10 12180 90
rect 12260 10 12270 90
rect 12170 0 12270 10
<< via3 >>
rect 6960 14160 7040 14170
rect 6960 14100 6970 14160
rect 6970 14100 7030 14160
rect 7030 14100 7040 14160
rect 6960 14090 7040 14100
rect 7080 12760 7160 12770
rect 7080 12700 7090 12760
rect 7090 12700 7150 12760
rect 7150 12700 7160 12760
rect 7080 12690 7160 12700
rect 7080 11360 7160 11370
rect 7080 11300 7090 11360
rect 7090 11300 7150 11360
rect 7150 11300 7160 11360
rect 7080 11290 7160 11300
rect 7050 8090 7130 8170
rect 1730 4930 1810 4940
rect 1730 4870 1740 4930
rect 1740 4870 1800 4930
rect 1800 4870 1810 4930
rect 1730 4860 1810 4870
rect 1430 3690 1510 3770
rect 7840 8160 7920 8170
rect 7840 8100 7850 8160
rect 7850 8100 7910 8160
rect 7910 8100 7920 8160
rect 7840 8090 7920 8100
rect 11770 7810 11840 7880
rect 11770 7310 11840 7380
rect 7210 6900 7290 6980
rect 7840 6970 7920 6980
rect 7840 6910 7850 6970
rect 7850 6910 7910 6970
rect 7910 6910 7920 6970
rect 7840 6900 7920 6910
rect 7210 4490 7290 4570
rect 7760 4560 7840 4570
rect 7760 4500 7770 4560
rect 7770 4500 7830 4560
rect 7830 4500 7840 4560
rect 7760 4490 7840 4500
rect 11370 3840 11440 3910
rect 11370 3430 11440 3500
rect 7050 2790 7130 2870
rect 1730 2590 1810 2600
rect 1730 2530 1740 2590
rect 1740 2530 1800 2590
rect 1800 2530 1810 2590
rect 1730 2520 1810 2530
rect 7760 2860 7840 2870
rect 7760 2800 7770 2860
rect 7770 2800 7830 2860
rect 7830 2800 7840 2860
rect 7760 2790 7840 2800
rect 17110 2660 17180 2730
rect 17610 2660 17680 2730
rect 12180 2160 12260 2170
rect 12180 2100 12190 2160
rect 12190 2100 12250 2160
rect 12250 2100 12260 2160
rect 12180 2090 12260 2100
rect 12180 1660 12260 1670
rect 12180 1600 12190 1660
rect 12190 1600 12250 1660
rect 12250 1600 12260 1660
rect 12180 1590 12260 1600
rect 1430 810 1510 890
rect 12180 860 12260 870
rect 12180 800 12190 860
rect 12190 800 12250 860
rect 12250 800 12260 860
rect 12180 790 12260 800
rect 12180 80 12260 90
rect 12180 20 12190 80
rect 12190 20 12250 80
rect 12250 20 12260 80
rect 12180 10 12260 20
<< mimcap >>
rect 7440 14870 7840 15020
rect 7440 14790 7610 14870
rect 7690 14790 7840 14870
rect 7440 14620 7840 14790
rect 8140 14870 8540 15020
rect 8140 14790 8300 14870
rect 8380 14790 8540 14870
rect 8140 14620 8540 14790
rect 8840 14870 9240 15020
rect 8840 14790 9000 14870
rect 9080 14790 9240 14870
rect 8840 14620 9240 14790
rect 9540 14870 9940 15020
rect 9540 14790 9700 14870
rect 9780 14790 9940 14870
rect 9540 14620 9940 14790
rect 10240 14870 10640 15020
rect 10240 14790 10400 14870
rect 10480 14790 10640 14870
rect 10240 14620 10640 14790
rect 10940 14870 11340 15020
rect 10940 14790 11100 14870
rect 11180 14790 11340 14870
rect 10940 14620 11340 14790
rect 11640 14870 12040 15020
rect 11640 14790 11800 14870
rect 11880 14790 12040 14870
rect 11640 14620 12040 14790
rect 12340 14870 12740 15020
rect 12340 14790 12500 14870
rect 12580 14790 12740 14870
rect 12340 14620 12740 14790
rect 13040 14870 13440 15020
rect 13040 14790 13200 14870
rect 13280 14790 13440 14870
rect 13040 14620 13440 14790
rect 13740 14870 14140 15020
rect 13740 14790 13900 14870
rect 13980 14790 14140 14870
rect 13740 14620 14140 14790
rect 7440 14170 7840 14320
rect 7440 14090 7610 14170
rect 7690 14090 7840 14170
rect 7440 13920 7840 14090
rect 8140 14170 8540 14320
rect 8140 14090 8300 14170
rect 8380 14090 8540 14170
rect 8140 13920 8540 14090
rect 8840 14170 9240 14320
rect 8840 14090 9000 14170
rect 9080 14090 9240 14170
rect 8840 13920 9240 14090
rect 9540 14170 9940 14320
rect 9540 14090 9700 14170
rect 9780 14090 9940 14170
rect 9540 13920 9940 14090
rect 10240 14170 10640 14320
rect 10240 14090 10400 14170
rect 10480 14090 10640 14170
rect 10240 13920 10640 14090
rect 10940 14170 11340 14320
rect 10940 14090 11100 14170
rect 11180 14090 11340 14170
rect 10940 13920 11340 14090
rect 11640 14170 12040 14320
rect 11640 14090 11800 14170
rect 11880 14090 12040 14170
rect 11640 13920 12040 14090
rect 12340 14170 12740 14320
rect 12340 14090 12500 14170
rect 12580 14090 12740 14170
rect 12340 13920 12740 14090
rect 13040 14170 13440 14320
rect 13040 14090 13200 14170
rect 13280 14090 13440 14170
rect 13040 13920 13440 14090
rect 13740 14170 14140 14320
rect 13740 14090 13900 14170
rect 13980 14090 14140 14170
rect 13740 13920 14140 14090
rect 7440 13470 7840 13620
rect 7440 13390 7610 13470
rect 7690 13390 7840 13470
rect 7440 13220 7840 13390
rect 8140 13470 8540 13620
rect 8140 13390 8300 13470
rect 8380 13390 8540 13470
rect 8140 13220 8540 13390
rect 8840 13470 9240 13620
rect 8840 13390 9000 13470
rect 9080 13390 9240 13470
rect 8840 13220 9240 13390
rect 9540 13470 9940 13620
rect 9540 13390 9700 13470
rect 9780 13390 9940 13470
rect 9540 13220 9940 13390
rect 10240 13470 10640 13620
rect 10240 13390 10400 13470
rect 10480 13390 10640 13470
rect 10240 13220 10640 13390
rect 10940 13470 11340 13620
rect 10940 13390 11100 13470
rect 11180 13390 11340 13470
rect 10940 13220 11340 13390
rect 11640 13470 12040 13620
rect 11640 13390 11800 13470
rect 11880 13390 12040 13470
rect 11640 13220 12040 13390
rect 12340 13470 12740 13620
rect 12340 13390 12500 13470
rect 12580 13390 12740 13470
rect 12340 13220 12740 13390
rect 13040 13470 13440 13620
rect 13040 13390 13200 13470
rect 13280 13390 13440 13470
rect 13040 13220 13440 13390
rect 13740 13470 14140 13620
rect 13740 13390 13900 13470
rect 13980 13390 14140 13470
rect 13740 13220 14140 13390
rect 7440 12770 7840 12920
rect 7440 12690 7610 12770
rect 7690 12690 7840 12770
rect 7440 12520 7840 12690
rect 8140 12770 8540 12920
rect 8140 12690 8300 12770
rect 8380 12690 8540 12770
rect 8140 12520 8540 12690
rect 8840 12770 9240 12920
rect 8840 12690 9000 12770
rect 9080 12690 9240 12770
rect 8840 12520 9240 12690
rect 9540 12770 9940 12920
rect 9540 12690 9700 12770
rect 9780 12690 9940 12770
rect 9540 12520 9940 12690
rect 10240 12770 10640 12920
rect 10240 12690 10400 12770
rect 10480 12690 10640 12770
rect 10240 12520 10640 12690
rect 10940 12770 11340 12920
rect 10940 12690 11100 12770
rect 11180 12690 11340 12770
rect 10940 12520 11340 12690
rect 11640 12770 12040 12920
rect 11640 12690 11800 12770
rect 11880 12690 12040 12770
rect 11640 12520 12040 12690
rect 12340 12770 12740 12920
rect 12340 12690 12500 12770
rect 12580 12690 12740 12770
rect 12340 12520 12740 12690
rect 13040 12770 13440 12920
rect 13040 12690 13200 12770
rect 13280 12690 13440 12770
rect 13040 12520 13440 12690
rect 13740 12770 14140 12920
rect 13740 12690 13900 12770
rect 13980 12690 14140 12770
rect 13740 12520 14140 12690
rect 7440 12070 7840 12220
rect 7440 11990 7610 12070
rect 7690 11990 7840 12070
rect 7440 11820 7840 11990
rect 8140 12070 8540 12220
rect 8140 11990 8300 12070
rect 8380 11990 8540 12070
rect 8140 11820 8540 11990
rect 8840 12070 9240 12220
rect 8840 11990 9000 12070
rect 9080 11990 9240 12070
rect 8840 11820 9240 11990
rect 9540 12070 9940 12220
rect 9540 11990 9700 12070
rect 9780 11990 9940 12070
rect 9540 11820 9940 11990
rect 10240 12070 10640 12220
rect 10240 11990 10400 12070
rect 10480 11990 10640 12070
rect 10240 11820 10640 11990
rect 10940 12070 11340 12220
rect 10940 11990 11100 12070
rect 11180 11990 11340 12070
rect 10940 11820 11340 11990
rect 11640 12070 12040 12220
rect 11640 11990 11800 12070
rect 11880 11990 12040 12070
rect 11640 11820 12040 11990
rect 12340 12070 12740 12220
rect 12340 11990 12500 12070
rect 12580 11990 12740 12070
rect 12340 11820 12740 11990
rect 13040 12070 13440 12220
rect 13040 11990 13200 12070
rect 13280 11990 13440 12070
rect 13040 11820 13440 11990
rect 13740 12070 14140 12220
rect 13740 11990 13900 12070
rect 13980 11990 14140 12070
rect 13740 11820 14140 11990
rect 7440 11370 7840 11520
rect 7440 11290 7610 11370
rect 7690 11290 7840 11370
rect 7440 11120 7840 11290
rect 8140 11370 8540 11520
rect 8140 11290 8300 11370
rect 8380 11290 8540 11370
rect 8140 11120 8540 11290
rect 8840 11370 9240 11520
rect 8840 11290 9000 11370
rect 9080 11290 9240 11370
rect 8840 11120 9240 11290
rect 9540 11370 9940 11520
rect 9540 11290 9700 11370
rect 9780 11290 9940 11370
rect 9540 11120 9940 11290
rect 10240 11370 10640 11520
rect 10240 11290 10400 11370
rect 10480 11290 10640 11370
rect 10240 11120 10640 11290
rect 10940 11370 11340 11520
rect 10940 11290 11100 11370
rect 11180 11290 11340 11370
rect 10940 11120 11340 11290
rect 11640 11370 12040 11520
rect 11640 11290 11800 11370
rect 11880 11290 12040 11370
rect 11640 11120 12040 11290
rect 12340 11370 12740 11520
rect 12340 11290 12500 11370
rect 12580 11290 12740 11370
rect 12340 11120 12740 11290
rect 13040 11370 13440 11520
rect 13040 11290 13200 11370
rect 13280 11290 13440 11370
rect 13040 11120 13440 11290
rect 13740 11370 14140 11520
rect 13740 11290 13900 11370
rect 13980 11290 14140 11370
rect 13740 11120 14140 11290
rect 12130 7880 14130 9790
rect 12130 7810 12150 7880
rect 12220 7810 14130 7880
rect 12130 7790 14130 7810
rect 12130 7380 14130 7400
rect 12130 7310 12150 7380
rect 12220 7310 14130 7380
rect 12130 5400 14130 7310
rect 11730 3910 12770 5080
rect 11730 3840 11750 3910
rect 11820 3840 12770 3910
rect 11730 3820 12770 3840
rect 11730 3500 12270 3520
rect 11730 3430 11750 3500
rect 11820 3430 12270 3500
rect 11730 2760 12270 3430
rect 14440 3110 17200 15020
rect 14440 3040 17110 3110
rect 17180 3040 17200 3110
rect 14440 3020 17200 3040
rect 17590 3110 31550 15020
rect 17590 3040 17610 3110
rect 17680 3040 31550 3110
rect 17590 3020 31550 3040
<< mimcapcontact >>
rect 7610 14790 7690 14870
rect 8300 14790 8380 14870
rect 9000 14790 9080 14870
rect 9700 14790 9780 14870
rect 10400 14790 10480 14870
rect 11100 14790 11180 14870
rect 11800 14790 11880 14870
rect 12500 14790 12580 14870
rect 13200 14790 13280 14870
rect 13900 14790 13980 14870
rect 7610 14090 7690 14170
rect 8300 14090 8380 14170
rect 9000 14090 9080 14170
rect 9700 14090 9780 14170
rect 10400 14090 10480 14170
rect 11100 14090 11180 14170
rect 11800 14090 11880 14170
rect 12500 14090 12580 14170
rect 13200 14090 13280 14170
rect 13900 14090 13980 14170
rect 7610 13390 7690 13470
rect 8300 13390 8380 13470
rect 9000 13390 9080 13470
rect 9700 13390 9780 13470
rect 10400 13390 10480 13470
rect 11100 13390 11180 13470
rect 11800 13390 11880 13470
rect 12500 13390 12580 13470
rect 13200 13390 13280 13470
rect 13900 13390 13980 13470
rect 7610 12690 7690 12770
rect 8300 12690 8380 12770
rect 9000 12690 9080 12770
rect 9700 12690 9780 12770
rect 10400 12690 10480 12770
rect 11100 12690 11180 12770
rect 11800 12690 11880 12770
rect 12500 12690 12580 12770
rect 13200 12690 13280 12770
rect 13900 12690 13980 12770
rect 7610 11990 7690 12070
rect 8300 11990 8380 12070
rect 9000 11990 9080 12070
rect 9700 11990 9780 12070
rect 10400 11990 10480 12070
rect 11100 11990 11180 12070
rect 11800 11990 11880 12070
rect 12500 11990 12580 12070
rect 13200 11990 13280 12070
rect 13900 11990 13980 12070
rect 7610 11290 7690 11370
rect 8300 11290 8380 11370
rect 9000 11290 9080 11370
rect 9700 11290 9780 11370
rect 10400 11290 10480 11370
rect 11100 11290 11180 11370
rect 11800 11290 11880 11370
rect 12500 11290 12580 11370
rect 13200 11290 13280 11370
rect 13900 11290 13980 11370
rect 12150 7810 12220 7880
rect 12150 7310 12220 7380
rect 11750 3840 11820 3910
rect 11750 3430 11820 3500
rect 17110 3040 17180 3110
rect 17610 3040 17680 3110
<< metal4 >>
rect 7600 14870 13990 14880
rect 7600 14790 7610 14870
rect 7690 14790 8300 14870
rect 8380 14790 9000 14870
rect 9080 14790 9700 14870
rect 9780 14790 10400 14870
rect 10480 14790 11100 14870
rect 11180 14790 11800 14870
rect 11880 14790 12500 14870
rect 12580 14790 13200 14870
rect 13280 14790 13900 14870
rect 13980 14790 13990 14870
rect 7600 14780 13990 14790
rect 13890 14180 13990 14780
rect 6950 14170 13990 14180
rect 6950 14090 6960 14170
rect 7040 14090 7610 14170
rect 7690 14090 8300 14170
rect 8380 14090 9000 14170
rect 9080 14090 9700 14170
rect 9780 14090 10400 14170
rect 10480 14090 11100 14170
rect 11180 14090 11800 14170
rect 11880 14090 12500 14170
rect 12580 14090 13200 14170
rect 13280 14090 13900 14170
rect 13980 14090 13990 14170
rect 6950 14080 13990 14090
rect 7600 13470 13990 13480
rect 7600 13390 7610 13470
rect 7690 13390 8300 13470
rect 8380 13390 9000 13470
rect 9080 13390 9700 13470
rect 9780 13390 10400 13470
rect 10480 13390 11100 13470
rect 11180 13390 11800 13470
rect 11880 13390 12500 13470
rect 12580 13390 13200 13470
rect 13280 13390 13900 13470
rect 13980 13390 13990 13470
rect 7600 13380 13990 13390
rect 13890 12780 13990 13380
rect 7070 12770 13990 12780
rect 7070 12690 7080 12770
rect 7160 12690 7610 12770
rect 7690 12690 8300 12770
rect 8380 12690 9000 12770
rect 9080 12690 9700 12770
rect 9780 12690 10400 12770
rect 10480 12690 11100 12770
rect 11180 12690 11800 12770
rect 11880 12690 12500 12770
rect 12580 12690 13200 12770
rect 13280 12690 13900 12770
rect 13980 12690 13990 12770
rect 7070 12680 13990 12690
rect 7600 12070 13990 12080
rect 7600 11990 7610 12070
rect 7690 11990 8300 12070
rect 8380 11990 9000 12070
rect 9080 11990 9700 12070
rect 9780 11990 10400 12070
rect 10480 11990 11100 12070
rect 11180 11990 11800 12070
rect 11880 11990 12500 12070
rect 12580 11990 13200 12070
rect 13280 11990 13900 12070
rect 13980 11990 13990 12070
rect 7600 11980 13990 11990
rect 13890 11380 13990 11980
rect 7070 11370 13990 11380
rect 7070 11290 7080 11370
rect 7160 11290 7610 11370
rect 7690 11290 8300 11370
rect 8380 11290 9000 11370
rect 9080 11290 9700 11370
rect 9780 11290 10400 11370
rect 10480 11290 11100 11370
rect 11180 11290 11800 11370
rect 11880 11290 12500 11370
rect 12580 11290 13200 11370
rect 13280 11290 13900 11370
rect 13980 11290 13990 11370
rect 7070 11280 13990 11290
rect 7040 8170 7930 8180
rect 7040 8090 7050 8170
rect 7130 8090 7840 8170
rect 7920 8090 7930 8170
rect 7040 8080 7930 8090
rect 11750 7880 12230 7900
rect 11750 7810 11770 7880
rect 11840 7810 12150 7880
rect 12220 7810 12230 7880
rect 11750 7790 12230 7810
rect 11750 7380 12230 7400
rect 11750 7310 11770 7380
rect 11840 7310 12150 7380
rect 12220 7310 12230 7380
rect 11750 7290 12230 7310
rect 7200 6980 7930 6990
rect 7200 6900 7210 6980
rect 7290 6900 7840 6980
rect 7920 6900 7930 6980
rect 7200 6890 7930 6900
rect 1720 4940 1820 4950
rect 1720 4860 1730 4940
rect 1810 4860 1820 4940
rect 1420 3770 1520 3780
rect 1420 3690 1430 3770
rect 1510 3690 1520 3770
rect 1420 890 1520 3690
rect 1720 2600 1820 4860
rect 7200 4570 7850 4580
rect 7200 4490 7210 4570
rect 7290 4490 7760 4570
rect 7840 4490 7850 4570
rect 7200 4480 7850 4490
rect 11350 3910 11840 3930
rect 11350 3840 11370 3910
rect 11440 3840 11750 3910
rect 11820 3840 11840 3910
rect 11350 3820 11840 3840
rect 11350 3500 11840 3520
rect 11350 3430 11370 3500
rect 11440 3430 11750 3500
rect 11820 3430 11840 3500
rect 11350 3410 11840 3430
rect 17090 3110 17200 3120
rect 17090 3040 17110 3110
rect 17180 3040 17200 3110
rect 7040 2870 7850 2880
rect 7040 2790 7050 2870
rect 7130 2790 7760 2870
rect 7840 2790 7850 2870
rect 7040 2780 7850 2790
rect 17090 2730 17200 3040
rect 17090 2660 17110 2730
rect 17180 2660 17200 2730
rect 17090 2640 17200 2660
rect 17590 3110 17700 3120
rect 17590 3040 17610 3110
rect 17680 3040 17700 3110
rect 17590 2730 17700 3040
rect 17590 2660 17610 2730
rect 17680 2660 17700 2730
rect 17590 2640 17700 2660
rect 1720 2520 1730 2600
rect 1810 2520 1820 2600
rect 1720 2510 1820 2520
rect 12170 2170 12270 2180
rect 12170 2090 12180 2170
rect 12260 2090 12270 2170
rect 12170 1670 12270 2090
rect 12170 1590 12180 1670
rect 12260 1590 12270 1670
rect 12170 1580 12270 1590
rect 1420 810 1430 890
rect 1510 810 1520 890
rect 1420 800 1520 810
rect 12170 870 12270 880
rect 12170 790 12180 870
rect 12260 790 12270 870
rect 12170 90 12270 790
rect 12170 10 12180 90
rect 12260 10 12270 90
rect 12170 0 12270 10
<< end >>
