* NGSPICE file created from pll_bgr_magic_3_flat.ext - technology: sky130A

.subckt pll_bgr_magic_3_flat
X0 a_2030_8210# a_1850_9420# w_n760_8620# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X1 w_n2590_4470# a_n2150_4460# a_n2150_4460# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X2 a_n1559_3570# a_n2860_n962# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X3 a_n10_8660# a_n530_8240# a_n450_8210# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X4 w_n760_8620# a_970_8210# a_890_9420# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X5 a_n1110_5640# w_n2590_4470# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6 a_990_12440# a_n220_12480# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X7 a_6200_5810# a_6200_5810# a_6200_5810# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=2.5 ps=17 w=0.5 l=0.15
X8 w_n1587_n2327# a_6080_5220# a_6080_5220# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X9 a_70_8210# a_450_8210# a_370_8660# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X10 w_n1587_n2327# a_990_12440# a_410_12110# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X11 a_760_4400# a_3480_n1988# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X12 a_3400_8240# a_3010_8240# w_n760_8620# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X13 a_250_12540# a_410_12110# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X14 w_n1587_n2327# w_n1587_n2327# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=100.167 ps=594.6 w=2 l=0.6
X15 a_2620_8240# a_n450_8210# w_n760_8620# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X16 w_n1550_12150# a_5660_12350# a_5250_12520# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X17 a_2760_12400# a_2870_12480# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X18 w_n2590_4470# a_890_4460# a_890_4460# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X19 w_n2590_4470# w_n2590_4470# a_n2740_n910# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X20 a_3560_12540# a_3530_12190# a_3450_12540# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X21 w_n2590_4470# a_n2860_n962# a_650_6670# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X22 a_5850_4590# a_6080_9390# a_6370_4590# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X23 a_0_12190# a_n1250_12490# w_n1550_12150# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X24 w_n760_8620# a_2030_8210# a_1700_8210# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X25 a_3560_9420# a_9240_3474# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X26 a_n1110_5640# w_n2590_4470# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X27 a_n2250_2660# a_n2740_n910# a_n2150_4460# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X28 w_n760_8620# a_70_8210# a_n10_8660# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X29 a_n450_8210# a_n530_8240# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X30 w_n1587_n2327# a_450_8210# a_70_8210# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X31 w_n1587_n2327# a_6100_5780# a_6200_5810# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X32 a_n2280_4390# a_n2150_4460# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X33 a_3400_8240# a_3010_8240# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X34 a_3690_9420# a_3010_9420# w_n760_8620# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X35 w_n1587_n2327# w_n1587_n2327# a_n1410_n2150# sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X36 a_n2280_4390# a_n2860_n1778# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X37 a_2620_8240# a_n450_8210# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X38 a_760_4400# a_3480_n1988# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 w_n1587_n2327# a_2030_8210# a_1700_8210# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X40 a_n2280_4390# a_n2860_n1778# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X41 a_4890_n2980# a_3690_9420# w_5500_9250# w_5500_9250# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X42 w_n1587_n2327# a_6100_5780# a_6100_5780# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X43 a_n1110_5640# w_n2590_4470# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X44 a_3010_9420# a_2620_9420# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X45 a_8640_12170# a_9930_11970# a_10340_10900# w_5500_9250# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X46 a_3560_9420# a_6370_4590# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X47 a_n1559_3570# a_n2860_n962# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X48 w_n1587_n2327# a_70_8210# a_n450_8210# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X49 a_8640_12170# a_9930_11970# a_10340_12730# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X50 a_n1830_2050# a_n1110_5640# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X51 a_9380_10870# a_4890_n2980# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X52 a_650_6670# a_n2860_n962# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X53 a_1050_3670# a_n2310_n530# a_760_4400# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X54 w_n1587_n2327# w_n1587_n2327# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X55 w_n2590_4470# a_n1110_5640# a_n2310_n530# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X56 w_n2590_4470# w_n2590_4470# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=41 ps=246.5 w=1 l=0.15
X57 m2_n4270_n3380# a_2978_n2980# sky130_fd_pr__cap_mim_m3_1 l=60 w=69.8
X58 a_760_4400# a_3480_n1988# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X59 a_n1110_5640# a_3480_n1988# w_n1587_n2327# sky130_fd_pr__res_high_po_0p35 l=2.05
X60 a_n2150_4460# a_n2150_4460# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X61 w_n2590_4470# a_n1110_5640# a_n2310_n530# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X62 w_5500_9250# a_9380_10870# a_9820_10900# w_5500_9250# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X63 a_2460_n530# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__res_xhigh_po_0p35 l=6
X64 w_n2590_4470# a_760_4400# a_n1110_5640# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X65 a_n2280_4390# a_n1559_3570# a_n2250_2660# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X66 w_n1587_n2327# a_2760_12400# a_2400_12190# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X67 w_n2590_4470# a_n2150_4460# a_n2280_4390# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X68 a_n2310_n530# a_n2310_n2138# w_n1587_n2327# sky130_fd_pr__res_xhigh_po_0p35 l=6
X69 a_3010_9420# a_2620_9420# w_n760_8620# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X70 a_n2150_4460# a_n2150_4460# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X71 w_5500_9250# w_5500_9250# w_5500_9250# w_5500_9250# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=14.4 ps=77.6 w=2 l=0.6
X72 w_n760_8620# a_n450_9390# a_1410_9420# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X73 w_5500_9250# w_n1587_n2327# a_9300_10900# w_5500_9250# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X74 a_n1110_5640# a_n1830_2050# a_n470_5670# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X75 w_n1587_n2327# a_4740_12170# a_5960_12630# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X76 a_6370_4590# a_6080_9390# a_5850_4590# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X77 a_5404_6290# a_6100_5780# sky130_fd_pr__res_generic_po w=0.33 l=2.4
X78 a_n530_9420# a_n760_9890# w_n760_8620# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X79 w_n2590_4470# a_5404_6290# a_5404_6290# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X80 a_n1110_5640# a_760_4400# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X81 a_5340_12190# a_6040_12170# w_n1550_12150# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X82 a_650_6670# w_n2590_4470# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X83 w_n1587_n2327# a_650_6670# a_6080_9390# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X84 a_4890_n2980# a_3690_8240# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X85 w_n760_8620# a_1370_8210# a_970_8210# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X86 w_n760_8620# a_970_8210# a_890_8660# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X87 a_n1110_5640# w_n2590_4470# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X88 a_n1110_5640# w_n2590_4470# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X89 w_n1587_n2327# w_n1587_n2327# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X90 a_n2150_4460# a_n2740_n910# a_n2250_2660# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X91 a_2620_9420# a_n450_9390# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X92 a_7260_12630# a_6640_12190# a_6960_12350# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X93 w_n2590_4470# a_5404_6290# a_5850_4590# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X94 w_n1587_n2327# a_4890_n2980# a_9300_12730# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X95 a_n220_12480# a_2400_12190# w_n1550_12150# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X96 a_n1110_5640# w_n2590_4470# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X97 w_n1550_12150# a_7340_12170# a_6640_12190# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X98 a_n1110_5640# a_760_4400# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X99 a_760_4400# a_3480_n1988# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X100 a_n330_12400# a_n220_12480# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X101 w_n1587_n2327# w_n1587_n2327# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X102 a_1050_3670# w_n2590_4470# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1.01 ps=6.15 w=2.5 l=5
X103 w_n1587_n2327# a_n1380_12430# a_n1510_12230# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X104 w_n1587_n2327# w_n1587_n2327# a_n1410_n2150# sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X105 a_n1380_12430# a_n1250_12490# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X106 a_n2280_4390# a_n2860_n1778# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X107 w_n1587_n2327# a_1370_8210# a_970_8210# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X108 w_n1587_n2327# a_970_8210# a_450_8210# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X109 a_n470_5670# a_n1110_5640# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X110 a_3950_12440# a_2870_12480# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X111 a_2870_12480# a_4740_12170# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X112 a_7940_12190# a_8640_12170# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X113 w_n2590_4470# a_7220_4560# a_7510_4590# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X114 a_760_4400# a_890_4460# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X115 w_n2590_4470# a_7510_4590# a_3560_9420# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X116 a_2978_n2980# a_4890_n2980# w_n1587_n2327# sky130_fd_pr__res_xhigh_po_0p35 l=7.52
X117 m2_n4270_n3380# a_4890_n2980# sky130_fd_pr__cap_mim_m3_1 l=60 w=13.8
X118 a_760_4400# a_3480_n1988# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X119 a_890_4460# a_n470_5670# a_1050_3670# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X120 w_n2590_4470# a_n1110_5640# a_n2740_n910# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X121 w_n1550_12150# a_5340_12190# a_4740_12170# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X122 w_5500_9250# a_9380_10870# a_10340_10900# w_5500_9250# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X123 a_5850_4590# a_5404_6290# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X124 a_1700_12190# a_n1250_12490# w_n1550_12150# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X125 w_n1587_n2327# w_n1587_n2327# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X126 a_6960_12350# a_6040_12170# w_n1550_12150# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X127 w_n1587_n2327# a_5250_12520# a_4740_12170# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X128 w_n1587_n2327# w_n1587_n2327# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X129 w_n2590_4470# a_n2280_4390# a_n2860_n962# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X130 w_n1587_n2327# w_5500_9250# a_9300_12730# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X131 a_1850_9420# a_1410_9420# w_n760_8620# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X132 a_760_4400# a_3480_n1988# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X133 a_760_4400# a_890_4460# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X134 a_3690_8240# a_3010_8240# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X135 a_n2280_4390# a_n2860_n1778# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X136 a_n2280_4390# a_n2150_4460# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X137 a_5404_6290# a_5404_6290# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X138 a_760_4400# a_n2310_n530# a_1050_3670# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X139 a_n2280_4390# a_n2860_n1778# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X140 a_5850_4590# a_4890_n2980# a_6080_5220# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X141 a_760_4400# a_3480_n1988# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X142 w_n2590_4470# w_n2590_4470# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X143 a_n750_12540# a_n1250_12490# a_n860_12540# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X144 a_n470_5670# a_2580_n2138# w_n1587_n2327# sky130_fd_pr__res_xhigh_po_0p35 l=6
X145 a_n1110_5640# w_n2590_4470# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X146 w_n1550_12150# a_4360_12350# a_3950_12440# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X147 w_n1587_n2327# a_6640_12190# a_6550_12520# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X148 a_1410_9420# a_n450_9390# a_1410_10040# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X149 w_n1550_12150# a_8260_12350# a_7850_12520# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X150 w_n760_8620# a_1700_8210# a_1370_8210# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X151 a_6550_12520# a_6640_12190# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X152 w_n2590_4470# a_n2280_4390# a_n2860_n962# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X153 a_760_4400# a_3480_n1988# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X154 w_n2590_4470# a_n1110_5640# a_n470_5670# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X155 a_760_4400# a_n2310_n530# a_1050_3670# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X156 w_5500_9250# a_9380_10870# a_9380_10870# w_5500_9250# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X157 a_n1110_5640# w_n2590_4470# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 a_n2280_4390# a_n2860_n1778# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X159 w_n1587_n2327# w_n1587_n2327# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X160 a_7510_4590# a_6080_9390# a_6200_5810# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X161 w_n2590_4470# a_760_4400# a_n1110_5640# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X162 w_n1587_n2327# a_n220_12480# a_990_12440# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X163 a_0_12190# a_n220_12480# a_580_12540# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X164 a_n2280_4390# a_n2860_n1778# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X165 a_3010_8240# w_n1587_n2327# a_2620_8240# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X166 w_n1587_n2327# a_n1510_12230# a_250_12540# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X167 a_7850_12520# a_7940_12190# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X168 a_3450_12540# a_2400_12190# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X169 w_n1587_n2327# a_1700_8210# a_1370_8210# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X170 a_370_9420# a_n530_10040# w_n760_8620# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X171 w_n1550_12150# a_410_12110# a_360_12220# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X172 a_n2250_2660# a_n1559_3570# a_n2280_4390# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X173 w_n2590_4470# a_n2860_n962# a_650_6670# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X174 a_n2150_4460# a_n2150_4460# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X175 w_n1587_n2327# a_8360_8230# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X176 a_2760_12400# a_3090_12190# w_n1550_12150# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X177 w_n1587_n2327# w_n2590_4470# a_n1110_5640# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=1.01 pd=6.15 as=1 ps=5.8 w=2.5 l=5
X178 a_n530_8660# a_n1510_12230# w_n760_8620# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X179 a_3090_12190# a_3530_12190# w_n1550_12150# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X180 a_250_2050# a_n1830_2050# a_n1830_2050# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X181 a_n2150_4460# a_n2740_n910# a_n2250_2660# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X182 a_n2190_n530# a_n2310_n2138# w_n1587_n2327# sky130_fd_pr__res_xhigh_po_0p35 l=6
X183 a_n330_12400# a_n220_12480# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X184 w_n1587_n2327# a_450_9390# a_70_9390# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X185 a_3560_9420# a_7510_4590# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X186 a_3010_8240# w_n760_8620# a_2620_8240# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X187 w_5500_9250# w_5500_9250# w_5500_9250# w_5500_9250# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X188 a_3690_9420# a_3400_9420# a_3560_9420# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X189 a_n2310_n530# a_n1110_5640# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X190 a_6080_5220# a_6080_5220# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X191 w_n2590_4470# a_890_4460# a_760_4400# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X192 w_n1587_n2327# w_n1587_n2327# a_n1410_n2150# sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X193 a_n2280_4390# a_n2860_n1778# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X194 a_n530_8240# a_n1510_12230# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X195 w_n1587_n2327# a_250_2050# a_250_2050# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X196 w_n1587_n2327# a_6370_4590# a_3560_9420# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X197 a_1050_3670# a_n470_5670# a_890_4460# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X198 a_n1559_3570# a_n2860_n962# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X199 w_n1587_n2327# w_n1587_n2327# a_n470_5670# sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X200 w_n2590_4470# a_n2860_n962# a_n1559_3570# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X201 a_n1830_2050# a_n1110_5640# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X202 a_n2860_n962# a_n2280_4390# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X203 a_n2280_4390# a_n1559_3570# a_n2250_2660# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X204 w_n2590_4470# a_890_4460# a_760_4400# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X205 w_n2590_4470# a_n2860_n962# a_650_6670# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X206 w_n1587_n2327# a_6100_5780# a_6100_5780# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X207 w_n1587_n2327# a_970_8210# a_450_9390# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X208 w_n1587_n2327# a_3690_8240# a_4890_n2980# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X209 a_n1410_n2150# a_n2310_n530# w_n1587_n2327# sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X210 w_n2590_4470# a_n2150_4460# a_n2150_4460# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X211 w_n2590_4470# a_n2860_n962# a_n1559_3570# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X212 a_n2280_4390# a_n2860_n1778# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X213 a_n2620_n910# a_n2740_n1988# w_n1587_n2327# sky130_fd_pr__res_xhigh_po_0p35 l=3.35
X214 w_n1587_n2327# a_2870_12480# a_2760_12400# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X215 a_n1110_5640# w_n2590_4470# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X216 a_760_4400# a_3480_n1988# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X217 a_6200_5810# a_4890_n2980# a_7220_4560# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X218 w_n1587_n2327# a_6100_5780# a_6200_5810# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X219 w_5500_9250# a_3560_9420# a_6080_9390# w_5500_9250# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X220 a_n2860_n962# w_n2590_4470# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X221 a_1050_3670# a_n2310_n530# a_760_4400# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X222 a_650_6670# a_n2860_n962# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X223 a_5850_4590# a_5850_4590# a_5850_4590# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=5 ps=27 w=1 l=0.15
X224 a_n1110_5640# w_n2590_4470# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.45 ps=2.9 w=1 l=0.15
X225 a_n2280_4390# a_n2150_4460# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X226 a_n1559_3570# a_n2860_n962# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X227 a_n1110_5640# w_n2590_4470# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X228 w_n1550_12150# a_6040_12170# a_5340_12190# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X229 w_n2590_4470# a_n2280_4390# a_n2860_n962# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X230 w_n2590_4470# w_n2590_4470# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X231 w_n1587_n2327# a_2400_12190# a_n220_12480# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X232 w_n1587_n2327# w_n1587_n2327# a_n1410_n2150# sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X233 a_760_4400# a_3480_n1988# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X234 a_n2250_2660# a_n1559_3570# a_n2280_4390# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X235 a_n2740_n910# a_n1110_5640# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X236 a_6640_12190# a_7340_12170# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X237 a_6200_5810# a_6100_5780# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X238 a_2030_8210# a_1850_9420# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X239 a_n1110_5640# w_n2590_4470# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X240 w_n2590_4470# a_n2860_n962# a_n1559_3570# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X241 a_890_9420# a_70_9390# a_450_9390# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X242 a_9410_11970# a_8640_12170# a_9300_10900# w_5500_9250# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X243 w_n2590_4470# a_n1110_5640# a_n1830_2050# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X244 a_9410_11970# a_8640_12170# a_9300_12730# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X245 a_2460_n530# a_2580_n2138# w_n1587_n2327# sky130_fd_pr__res_xhigh_po_0p35 l=6
X246 a_370_8660# a_n530_8240# w_n760_8620# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X247 a_n1110_5640# w_n2590_4470# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X248 a_3560_9420# a_6370_4590# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X249 w_n2590_4470# a_n2860_n962# a_650_6670# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X250 w_n1587_n2327# a_n220_12480# a_n330_12400# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X251 a_760_4400# a_3480_n1988# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X252 a_6080_9390# a_3560_9420# w_5500_9250# w_5500_9250# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X253 w_n1550_12150# a_2870_12480# a_3530_12190# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X254 w_5500_9250# w_n1587_n2327# a_9820_10900# w_5500_9250# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X255 a_n1380_12430# a_n1250_12490# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X256 a_n2280_4390# a_n2860_n1778# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X257 a_890_4460# a_890_4460# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X258 a_6100_5780# a_6100_5780# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X259 a_650_6670# a_n2860_n962# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X260 w_n2590_4470# w_n2590_4470# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X261 w_n1587_n2327# a_n220_12480# a_4660_12540# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X262 w_n1587_n2327# a_7340_12170# a_8560_12630# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X263 a_n1559_3570# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__res_xhigh_po_0p35 l=1
X264 a_n2280_4390# a_n2860_n1778# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X265 a_n1110_5640# w_n2590_4470# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X266 w_n1587_n2327# a_650_6670# a_650_6670# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X267 a_3690_8240# a_3010_8240# a_650_6670# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X268 a_760_4400# a_3480_n1988# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X269 w_n1587_n2327# w_n1587_n2327# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X270 a_7940_12190# a_8640_12170# w_n1550_12150# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X271 a_2870_12480# a_4740_12170# w_n1550_12150# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X272 a_n2280_4390# a_n2860_n1778# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X273 a_70_8210# a_n530_8240# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X274 a_n530_10040# a_n760_9890# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X275 a_6100_5780# a_6100_5780# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X276 w_n2590_4470# a_n2150_4460# a_n2280_4390# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X277 a_n2250_2660# a_n2740_n910# a_n2150_4460# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X278 a_890_4460# a_890_4460# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X279 w_n1550_12150# a_n1250_12490# a_1700_12190# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X280 a_760_4400# a_3480_n1988# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X281 w_n1587_n2327# a_4890_n2980# a_9820_12730# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X282 a_1620_12540# a_n220_12480# a_1510_12540# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X283 w_n1587_n2327# a_5340_12190# a_5250_12520# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X284 a_5960_12630# a_5340_12190# a_5660_12350# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X285 w_n1587_n2327# a_1700_12190# a_1620_12540# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X286 a_5250_12520# a_5340_12190# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X287 a_7220_4560# a_4890_n2980# a_6200_5810# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X288 a_n2280_4390# a_n2860_n1778# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X289 w_n2590_4470# w_n2590_4470# a_n1110_5640# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X290 a_3690_8240# a_3400_8240# a_650_6670# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X291 a_n2740_n910# w_n2590_4470# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X292 w_n2590_4470# a_n2860_n962# a_n1559_3570# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X293 w_n1587_n2327# a_70_9390# a_n450_9390# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X294 a_5850_4590# a_5850_4590# a_5850_4590# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X295 a_7510_4590# a_7220_4560# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X296 w_n2590_4470# a_n2860_n962# a_650_6670# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X297 a_3690_9420# a_3400_9420# sky130_fd_pr__cap_mim_m3_1 l=6.3 w=5.2
X298 a_n1110_5640# w_n2590_4470# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X299 a_6080_9390# a_3560_9420# w_5500_9250# w_5500_9250# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X300 a_890_4460# a_n470_5670# a_1050_3670# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X301 w_n1587_n2327# a_n1510_12230# a_n750_12540# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X302 a_760_4400# a_3480_n1988# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X303 w_n2590_4470# a_n1110_5640# a_n2740_n910# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X304 a_6550_12520# a_6640_12190# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X305 a_1410_10040# a_n450_8210# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X306 a_1850_9420# a_1410_9420# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X307 a_n1110_5640# w_n2590_4470# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X308 a_4890_n2980# a_3690_9420# w_5500_9250# w_5500_9250# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X309 w_n1550_12150# a_n860_12540# a_n1380_12430# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X310 a_9240_6410# a_6370_4590# w_n1587_n2327# sky130_fd_pr__res_xhigh_po_0p35 l=0.86
X311 a_5404_6290# a_5404_6290# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X312 w_n2590_4470# a_760_4400# a_n1110_5640# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X313 a_650_6670# a_650_6670# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X314 a_n1110_5640# a_760_4400# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X315 w_n1550_12150# a_7940_12190# a_7340_12170# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X316 a_990_12440# a_n220_12480# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X317 a_n2280_4390# a_n2860_n1778# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X318 a_580_12540# a_n1250_12490# a_250_12540# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X319 a_n2860_n962# a_n2280_4390# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X320 w_n1587_n2327# w_5500_9250# a_9820_12730# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X321 w_n1587_n2327# w_n1587_n2327# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.625 pd=3.5 as=0 ps=0 w=1.25 l=0.5
X322 a_5660_12350# a_4740_12170# w_n1550_12150# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X323 w_n1587_n2327# a_3950_12440# a_3530_12190# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X324 w_n1587_n2327# a_7850_12520# a_7340_12170# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X325 a_3090_12190# a_2870_12480# a_3560_12540# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X326 a_5850_4590# a_5404_6290# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X327 a_n2280_4390# a_n2860_n1778# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 a_360_12220# a_n1510_12230# a_0_12190# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X329 a_n1110_5640# w_n2590_4470# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X330 a_n2860_n962# w_n2590_4470# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X331 a_6080_5220# a_4890_n2980# a_5850_4590# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X332 a_n2620_n910# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__res_xhigh_po_0p35 l=3.35
X333 w_n2590_4470# a_890_4460# a_760_4400# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X334 a_1410_9420# a_n450_8210# w_n760_8620# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.805 ps=5 w=2 l=0.15
X335 w_5500_9250# w_n1587_n2327# a_10340_10900# w_5500_9250# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X336 w_n1550_12150# a_2400_12190# a_3090_12190# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X337 a_760_4400# a_3480_n1988# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X338 a_n1110_5640# w_n2590_4470# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X339 w_n2590_4470# a_7510_4590# a_3560_9420# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X340 a_n530_10040# a_n450_9390# a_n530_9420# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X341 a_70_9390# a_n530_10040# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X342 w_n2590_4470# w_n2590_4470# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0 ps=0 w=2.5 l=0.5
X343 w_n2590_4470# a_890_4460# a_890_4460# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X344 w_n1550_12150# a_6960_12350# a_6550_12520# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X345 a_n330_12400# a_0_12190# w_n1550_12150# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X346 w_n1587_n2327# a_6080_5220# a_6370_4590# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X347 w_5500_9250# a_5650_9820# w_5500_9250# w_5500_9250# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X348 w_5500_9250# a_9380_10870# a_9300_10900# w_5500_9250# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X349 w_n1587_n2327# w_n1587_n2327# a_n1410_n2150# sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X350 a_890_8660# a_70_8210# a_450_8210# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X351 w_5500_9250# a_3690_9420# a_4890_n2980# w_5500_9250# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X352 w_n1587_n2327# w_n1587_n2327# a_n1410_n2150# sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X353 a_n2280_4390# a_n2860_n1778# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X354 w_n1587_n2327# a_5450_8180# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X355 w_n1587_n2327# a_4890_n2980# a_10340_12730# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X356 w_n2590_4470# w_n2590_4470# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=1.25 pd=6 as=0 ps=0 w=2.5 l=0.5
X357 w_n2590_4470# a_n1110_5640# a_n470_5670# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X358 a_n2150_4460# a_n2740_n910# a_n2250_2660# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X359 w_n2590_4470# a_890_4460# a_890_4460# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X360 a_n2310_n530# a_n1110_5640# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X361 w_n1587_n2327# w_n1587_n2327# a_n1410_n2150# sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X362 w_n2590_4470# a_7220_4560# a_7220_4560# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X363 w_n1587_n2327# w_n1587_n2327# a_n1410_n2150# sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X364 a_450_8210# a_70_8210# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X365 a_450_9390# a_70_9390# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X366 a_3560_9420# a_9240_6410# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X367 w_n1550_12150# a_n1250_12490# a_n1510_12230# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X368 w_n2590_4470# a_5404_6290# a_5850_4590# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X369 a_1050_3670# a_n470_5670# a_890_4460# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X370 a_n2280_4390# a_n2860_n1778# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X371 a_2760_12400# a_2870_12480# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X372 a_1050_3670# a_n470_5670# a_890_4460# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X373 a_6200_5810# a_6200_5810# a_6200_5810# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X374 w_n1550_12150# a_n220_12480# a_410_12110# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X375 a_7510_4590# a_9240_3474# w_n1587_n2327# sky130_fd_pr__res_xhigh_po_0p35 l=1.14
X376 w_n2590_4470# a_5404_6290# a_5404_6290# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X377 a_n1110_5640# w_n2590_4470# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X378 a_n10_9420# a_n530_10040# a_n450_9390# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X379 w_n1550_12150# a_2870_12480# a_2400_12190# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X380 a_70_9390# a_450_9390# a_370_9420# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X381 a_n450_9390# a_n530_10040# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X382 a_3690_9420# a_3010_9420# a_3560_9420# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X383 w_n2590_4470# w_n2590_4470# a_n2860_n962# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X384 a_3400_9420# a_3010_9420# w_n760_8620# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X385 a_760_4400# a_890_4460# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X386 w_n1587_n2327# w_5500_9250# a_10340_12730# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X387 w_n2590_4470# w_n2590_4470# a_n1110_5640# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X388 w_5500_9250# a_8360_9360# w_5500_9250# w_5500_9250# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X389 a_2620_9420# a_n450_9390# w_n760_8620# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X390 a_n1110_5640# w_n2590_4470# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X391 a_5340_12190# a_6040_12170# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X392 a_760_4400# a_3480_n1988# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X393 a_n2280_4390# a_n2860_n1778# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X394 a_3400_9420# a_3010_9420# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X395 w_n760_8620# a_70_9390# a_n10_9420# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X396 a_3560_9420# a_7510_4590# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X397 a_760_4400# a_3480_n1988# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X398 a_760_4400# a_3480_n1988# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X399 a_890_4460# a_890_4460# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X400 a_6370_4590# a_6080_5220# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X401 a_n470_5670# a_n1110_5640# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X402 w_n2590_4470# w_n2590_4470# a_n1559_3570# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X403 w_n1587_n2327# a_6040_12170# a_7260_12630# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X404 w_n1550_12150# a_2400_12190# a_n220_12480# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X405 a_6640_12190# a_7340_12170# w_n1550_12150# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X406 a_n2860_n962# a_n2860_n1778# w_n1587_n2327# sky130_fd_pr__res_high_po_0p35 l=2.05
X407 w_n1587_n2327# a_n330_12400# a_n1250_12490# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X408 a_n2740_n910# a_n2740_n1988# w_n1587_n2327# sky130_fd_pr__res_xhigh_po_0p35 l=3.35
X409 a_n1559_3570# w_n2590_4470# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X410 a_760_4400# a_3480_n1988# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X411 w_n2590_4470# a_n2150_4460# a_n2280_4390# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X412 w_5500_9250# a_3560_9420# a_6080_9390# w_5500_9250# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X413 w_n1587_n2327# a_n1250_12490# a_n1380_12430# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X414 w_n1550_12150# a_n220_12480# a_n1250_12490# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X415 a_650_6670# a_n2860_n962# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X416 w_n1587_n2327# a_2870_12480# a_3950_12440# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X417 w_n1587_n2327# a_7940_12190# a_7850_12520# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X418 a_8560_12630# a_7940_12190# a_8260_12350# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X419 a_n2740_n910# a_n1110_5640# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X420 a_n530_8240# a_n450_8210# a_n530_8660# w_n760_8620# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X421 a_4660_12540# a_2870_12480# a_4360_12350# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X422 a_7850_12520# a_7940_12190# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X423 w_5500_9250# a_3690_9420# a_4890_n2980# w_5500_9250# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X424 a_3950_12440# a_2870_12480# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X425 a_3690_8240# a_3400_8240# sky130_fd_pr__cap_mim_m3_1 l=3.8 w=2.7
X426 a_7220_4560# a_7220_4560# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X427 w_n1550_12150# a_8640_12170# a_7940_12190# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X428 w_n1550_12150# a_4740_12170# a_2870_12480# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X429 w_n1587_n2327# a_n1250_12490# a_1700_12190# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X430 a_n1110_5640# w_n2590_4470# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X431 w_n1587_n2327# a_n450_9390# a_n530_10040# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X432 a_6080_9390# a_650_6670# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X433 w_n2590_4470# w_n2590_4470# a_650_6670# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X434 a_9930_11970# a_9410_11970# a_9820_10900# w_5500_9250# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X435 a_760_4400# a_n2310_n530# a_1050_3670# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X436 a_6200_5810# a_6080_9390# a_7510_4590# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X437 a_5250_12520# a_5340_12190# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X438 w_n1587_n2327# a_6370_4590# a_3560_9420# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X439 a_9930_11970# a_9410_11970# a_9820_12730# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X440 a_n1110_5640# w_n2590_4470# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X441 a_n2280_4390# a_n2860_n1778# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X442 w_n1587_n2327# a_n450_8210# a_n530_8240# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X443 a_n2190_n530# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__res_xhigh_po_0p35 l=6
X444 w_n1550_12150# a_1510_12540# a_990_12440# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X445 a_n470_5670# a_n1830_2050# a_n1110_5640# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X446 a_760_4400# a_3480_n1988# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X447 a_6200_5810# a_6100_5780# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X448 a_n2280_4390# a_n2860_n1778# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X449 w_n2590_4470# a_n2150_4460# a_n2150_4460# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X450 a_1510_12540# a_1700_12190# w_n1550_12150# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X451 w_n2590_4470# a_n2860_n962# a_n1559_3570# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X452 w_n1550_12150# a_6640_12190# a_6040_12170# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X453 a_n1559_3570# a_n2860_n962# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X454 a_n2250_2660# a_n1559_3570# a_n2280_4390# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X455 a_n2860_n962# a_n2280_4390# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X456 a_4360_12350# a_n220_12480# w_n1550_12150# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X457 w_n2590_4470# a_n1110_5640# a_n1830_2050# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X458 a_8260_12350# a_7340_12170# w_n1550_12150# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X459 w_n1587_n2327# a_6550_12520# a_6040_12170# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X460 w_n1587_n2327# w_n2590_4470# a_n2250_2660# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X461 a_650_6670# a_n2860_n962# w_n2590_4470# w_n2590_4470# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X462 w_n1587_n2327# w_n1587_n2327# w_n1587_n2327# w_n1587_n2327# sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0 ps=0 w=1.25 l=0.5
X463 a_n860_12540# a_n1510_12230# w_n1550_12150# w_n1550_12150# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
.ends

