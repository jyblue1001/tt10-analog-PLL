magic
tech sky130A
timestamp 1756780914
<< metal1 >>
rect 12150 9350 12350 9355
rect 12150 9320 12155 9350
rect 12185 9320 12195 9350
rect 12225 9320 12235 9350
rect 12265 9320 12275 9350
rect 12305 9320 12315 9350
rect 12345 9320 12350 9350
rect 12150 4085 12350 9320
rect 12150 4055 12155 4085
rect 12185 4055 12195 4085
rect 12225 4055 12235 4085
rect 12265 4055 12275 4085
rect 12305 4055 12315 4085
rect 12345 4055 12350 4085
rect 12150 4045 12350 4055
rect 12150 4015 12155 4045
rect 12185 4015 12195 4045
rect 12225 4015 12235 4045
rect 12265 4015 12275 4045
rect 12305 4015 12315 4045
rect 12345 4015 12350 4045
rect 12150 4005 12350 4015
rect 12150 3975 12155 4005
rect 12185 3975 12195 4005
rect 12225 3975 12235 4005
rect 12265 3975 12275 4005
rect 12305 3975 12315 4005
rect 12345 3975 12350 4005
rect 12150 3360 12350 3975
rect 12150 3330 12155 3360
rect 12185 3330 12195 3360
rect 12225 3330 12235 3360
rect 12265 3330 12275 3360
rect 12305 3330 12315 3360
rect 12345 3330 12350 3360
rect 5210 2915 5250 2920
rect 5210 2885 5215 2915
rect 5245 2885 5250 2915
rect 5210 665 5250 2885
rect 12150 1195 12350 3330
rect 12110 1155 12350 1195
rect 12150 1120 12350 1155
rect 12150 1090 12155 1120
rect 12185 1090 12195 1120
rect 12225 1090 12235 1120
rect 12265 1090 12275 1120
rect 12305 1090 12315 1120
rect 12345 1090 12350 1120
rect 12150 1085 12350 1090
rect 5210 635 5215 665
rect 5245 635 5250 665
rect 5210 630 5250 635
<< via1 >>
rect 12155 9320 12185 9350
rect 12195 9320 12225 9350
rect 12235 9320 12265 9350
rect 12275 9320 12305 9350
rect 12315 9320 12345 9350
rect 12155 4055 12185 4085
rect 12195 4055 12225 4085
rect 12235 4055 12265 4085
rect 12275 4055 12305 4085
rect 12315 4055 12345 4085
rect 12155 4015 12185 4045
rect 12195 4015 12225 4045
rect 12235 4015 12265 4045
rect 12275 4015 12305 4045
rect 12315 4015 12345 4045
rect 12155 3975 12185 4005
rect 12195 3975 12225 4005
rect 12235 3975 12265 4005
rect 12275 3975 12305 4005
rect 12315 3975 12345 4005
rect 12155 3330 12185 3360
rect 12195 3330 12225 3360
rect 12235 3330 12265 3360
rect 12275 3330 12305 3360
rect 12315 3330 12345 3360
rect 5215 2885 5245 2915
rect 12155 1090 12185 1120
rect 12195 1090 12225 1120
rect 12235 1090 12265 1120
rect 12275 1090 12305 1120
rect 12315 1090 12345 1120
rect 5215 635 5245 665
<< metal2 >>
rect 3890 9590 4020 9595
rect 3890 9560 3895 9590
rect 3925 9560 3940 9590
rect 3970 9560 3985 9590
rect 4015 9560 4020 9590
rect 3890 9545 4020 9560
rect 3890 9515 3895 9545
rect 3925 9515 3940 9545
rect 3970 9515 3985 9545
rect 4015 9515 4020 9545
rect 3890 9500 4020 9515
rect 3890 9470 3895 9500
rect 3925 9470 3940 9500
rect 3970 9470 3985 9500
rect 4015 9470 4020 9500
rect 3890 9465 4020 9470
rect 12150 9350 12350 9355
rect 12150 9320 12155 9350
rect 12185 9320 12195 9350
rect 12225 9320 12235 9350
rect 12265 9320 12275 9350
rect 12305 9320 12315 9350
rect 12345 9320 12350 9350
rect 12150 9315 12350 9320
rect 3890 9225 4905 9245
rect 3890 9195 3895 9225
rect 3925 9195 3940 9225
rect 3970 9195 3985 9225
rect 4015 9195 4905 9225
rect 3890 9175 4905 9195
rect 3890 9145 3895 9175
rect 3925 9145 3940 9175
rect 3970 9145 3985 9175
rect 4015 9145 4905 9175
rect 3890 9125 4905 9145
rect 12150 4085 12350 4090
rect 12150 4055 12155 4085
rect 12185 4055 12195 4085
rect 12225 4055 12235 4085
rect 12265 4055 12275 4085
rect 12305 4055 12315 4085
rect 12345 4055 12350 4085
rect 12150 4045 12350 4055
rect 12150 4015 12155 4045
rect 12185 4015 12195 4045
rect 12225 4015 12235 4045
rect 12265 4015 12275 4045
rect 12305 4015 12315 4045
rect 12345 4015 12350 4045
rect 12150 4005 12350 4015
rect 12150 3975 12155 4005
rect 12185 3975 12195 4005
rect 12225 3975 12235 4005
rect 12265 3975 12275 4005
rect 12305 3975 12315 4005
rect 12345 3975 12350 4005
rect 12150 3970 12350 3975
rect 12150 3360 12350 3365
rect 12150 3330 12155 3360
rect 12185 3330 12195 3360
rect 12225 3330 12235 3360
rect 12265 3330 12275 3360
rect 12305 3330 12315 3360
rect 12345 3330 12350 3360
rect 12150 3325 12350 3330
rect 11910 1480 12410 1600
rect 12150 1090 12155 1120
rect 12185 1090 12195 1120
rect 12225 1090 12235 1120
rect 12265 1090 12275 1120
rect 12305 1090 12315 1120
rect 12345 1090 12350 1120
rect 12150 1085 12350 1090
rect 15185 670 15265 690
rect 5210 665 15205 670
rect 5210 635 5215 665
rect 5245 635 15205 665
rect 5210 630 15205 635
rect 15245 630 15265 670
rect 15185 610 15265 630
<< via2 >>
rect 3895 9560 3925 9590
rect 3940 9560 3970 9590
rect 3985 9560 4015 9590
rect 3895 9515 3925 9545
rect 3940 9515 3970 9545
rect 3985 9515 4015 9545
rect 3895 9470 3925 9500
rect 3940 9470 3970 9500
rect 3985 9470 4015 9500
rect 3895 9195 3925 9225
rect 3940 9195 3970 9225
rect 3985 9195 4015 9225
rect 3895 9145 3925 9175
rect 3940 9145 3970 9175
rect 3985 9145 4015 9175
rect 15205 630 15245 670
<< metal3 >>
rect 400 9590 4020 9595
rect 400 9580 3895 9590
rect 400 9540 405 9580
rect 445 9540 455 9580
rect 495 9540 505 9580
rect 545 9540 555 9580
rect 595 9560 3895 9580
rect 3925 9560 3940 9590
rect 3970 9560 3985 9590
rect 4015 9560 4020 9590
rect 595 9545 4020 9560
rect 595 9540 3895 9545
rect 400 9520 3895 9540
rect 400 9480 405 9520
rect 445 9480 455 9520
rect 495 9480 505 9520
rect 545 9480 555 9520
rect 595 9515 3895 9520
rect 3925 9515 3940 9545
rect 3970 9515 3985 9545
rect 4015 9515 4020 9545
rect 595 9500 4020 9515
rect 595 9480 3895 9500
rect 400 9470 3895 9480
rect 3925 9470 3940 9500
rect 3970 9470 3985 9500
rect 4015 9470 4020 9500
rect 400 9465 4020 9470
rect 400 9230 4020 9245
rect 400 9190 405 9230
rect 445 9190 455 9230
rect 495 9190 505 9230
rect 545 9190 555 9230
rect 595 9225 4020 9230
rect 595 9195 3895 9225
rect 3925 9195 3940 9225
rect 3970 9195 3985 9225
rect 4015 9195 4020 9225
rect 595 9190 4020 9195
rect 400 9180 4020 9190
rect 400 9140 405 9180
rect 445 9140 455 9180
rect 495 9140 505 9180
rect 545 9140 555 9180
rect 595 9175 4020 9180
rect 595 9145 3895 9175
rect 3925 9145 3940 9175
rect 3970 9145 3985 9175
rect 4015 9145 4020 9175
rect 595 9140 4020 9145
rect 400 9125 4020 9140
rect 100 4205 4020 4220
rect 100 4165 105 4205
rect 145 4165 155 4205
rect 195 4165 205 4205
rect 245 4165 255 4205
rect 295 4165 4020 4205
rect 100 4155 4020 4165
rect 100 4115 105 4155
rect 145 4115 155 4155
rect 195 4115 205 4155
rect 245 4115 255 4155
rect 295 4115 4020 4155
rect 100 4100 4020 4115
rect 400 4055 4020 4070
rect 400 4015 405 4055
rect 445 4015 455 4055
rect 495 4015 505 4055
rect 545 4015 555 4055
rect 595 4015 4020 4055
rect 400 4005 4020 4015
rect 400 3965 405 4005
rect 445 3965 455 4005
rect 495 3965 505 4005
rect 545 3965 555 4005
rect 595 3965 4020 4005
rect 400 3950 4020 3965
rect 400 3880 4020 3895
rect 400 3840 405 3880
rect 445 3840 455 3880
rect 495 3840 505 3880
rect 545 3840 555 3880
rect 595 3840 4020 3880
rect 400 3830 4020 3840
rect 400 3790 405 3830
rect 445 3790 455 3830
rect 495 3790 505 3830
rect 545 3790 555 3830
rect 595 3790 4020 3830
rect 400 3775 4020 3790
rect 100 3290 4020 3305
rect 100 3250 105 3290
rect 145 3250 155 3290
rect 195 3250 205 3290
rect 245 3250 255 3290
rect 295 3250 4020 3290
rect 100 3240 4020 3250
rect 100 3200 105 3240
rect 145 3200 155 3240
rect 195 3200 205 3240
rect 245 3200 255 3240
rect 295 3200 4020 3240
rect 100 3185 4020 3200
rect 400 2700 4020 2715
rect 400 2660 405 2700
rect 445 2660 455 2700
rect 495 2660 505 2700
rect 545 2660 555 2700
rect 595 2660 4020 2700
rect 400 2650 4020 2660
rect 400 2610 405 2650
rect 445 2610 455 2650
rect 495 2610 505 2650
rect 545 2610 555 2650
rect 595 2610 4020 2650
rect 400 2595 4020 2610
rect 100 2550 4020 2565
rect 100 2510 105 2550
rect 145 2510 155 2550
rect 195 2510 205 2550
rect 245 2510 255 2550
rect 295 2510 4020 2550
rect 100 2500 4020 2510
rect 100 2460 105 2500
rect 145 2460 155 2500
rect 195 2460 205 2500
rect 245 2460 255 2500
rect 295 2460 4020 2500
rect 100 2445 4020 2460
rect 100 1790 4020 1805
rect 100 1750 105 1790
rect 145 1750 155 1790
rect 195 1750 205 1790
rect 245 1750 255 1790
rect 295 1750 4020 1790
rect 100 1740 4020 1750
rect 100 1700 105 1740
rect 145 1700 155 1740
rect 195 1700 205 1740
rect 245 1700 255 1740
rect 295 1700 4020 1740
rect 100 1685 4020 1700
rect 400 1400 4020 1415
rect 400 1360 405 1400
rect 445 1360 455 1400
rect 495 1360 505 1400
rect 545 1360 555 1400
rect 595 1360 4020 1400
rect 400 1350 4020 1360
rect 400 1310 405 1350
rect 445 1310 455 1350
rect 495 1310 505 1350
rect 545 1310 555 1350
rect 595 1310 4020 1350
rect 400 1295 4020 1310
rect 400 790 4020 805
rect 400 750 405 790
rect 445 750 455 790
rect 495 750 505 790
rect 545 750 555 790
rect 595 750 4020 790
rect 400 740 4020 750
rect 400 700 405 740
rect 445 700 455 740
rect 495 700 505 740
rect 545 700 555 740
rect 595 700 4020 740
rect 400 685 4020 700
rect 15185 670 15265 690
rect 15185 630 15205 670
rect 15245 630 15265 670
rect 15185 610 15265 630
<< via3 >>
rect 405 9540 445 9580
rect 455 9540 495 9580
rect 505 9540 545 9580
rect 555 9540 595 9580
rect 405 9480 445 9520
rect 455 9480 495 9520
rect 505 9480 545 9520
rect 555 9480 595 9520
rect 405 9190 445 9230
rect 455 9190 495 9230
rect 505 9190 545 9230
rect 555 9190 595 9230
rect 405 9140 445 9180
rect 455 9140 495 9180
rect 505 9140 545 9180
rect 555 9140 595 9180
rect 105 4165 145 4205
rect 155 4165 195 4205
rect 205 4165 245 4205
rect 255 4165 295 4205
rect 105 4115 145 4155
rect 155 4115 195 4155
rect 205 4115 245 4155
rect 255 4115 295 4155
rect 405 4015 445 4055
rect 455 4015 495 4055
rect 505 4015 545 4055
rect 555 4015 595 4055
rect 405 3965 445 4005
rect 455 3965 495 4005
rect 505 3965 545 4005
rect 555 3965 595 4005
rect 405 3840 445 3880
rect 455 3840 495 3880
rect 505 3840 545 3880
rect 555 3840 595 3880
rect 405 3790 445 3830
rect 455 3790 495 3830
rect 505 3790 545 3830
rect 555 3790 595 3830
rect 105 3250 145 3290
rect 155 3250 195 3290
rect 205 3250 245 3290
rect 255 3250 295 3290
rect 105 3200 145 3240
rect 155 3200 195 3240
rect 205 3200 245 3240
rect 255 3200 295 3240
rect 405 2660 445 2700
rect 455 2660 495 2700
rect 505 2660 545 2700
rect 555 2660 595 2700
rect 405 2610 445 2650
rect 455 2610 495 2650
rect 505 2610 545 2650
rect 555 2610 595 2650
rect 105 2510 145 2550
rect 155 2510 195 2550
rect 205 2510 245 2550
rect 255 2510 295 2550
rect 105 2460 145 2500
rect 155 2460 195 2500
rect 205 2460 245 2500
rect 255 2460 295 2500
rect 105 1750 145 1790
rect 155 1750 195 1790
rect 205 1750 245 1790
rect 255 1750 295 1790
rect 105 1700 145 1740
rect 155 1700 195 1740
rect 205 1700 245 1740
rect 255 1700 295 1740
rect 405 1360 445 1400
rect 455 1360 495 1400
rect 505 1360 545 1400
rect 555 1360 595 1400
rect 405 1310 445 1350
rect 455 1310 495 1350
rect 505 1310 545 1350
rect 555 1310 595 1350
rect 405 750 445 790
rect 455 750 495 790
rect 505 750 545 790
rect 555 750 595 790
rect 405 700 445 740
rect 455 700 495 740
rect 505 700 545 740
rect 555 700 595 740
rect 15205 630 15245 670
<< metal4 >>
rect 100 4205 300 22076
rect 100 4165 105 4205
rect 145 4165 155 4205
rect 195 4165 205 4205
rect 245 4165 255 4205
rect 295 4165 300 4205
rect 100 4155 300 4165
rect 100 4115 105 4155
rect 145 4115 155 4155
rect 195 4115 205 4155
rect 245 4115 255 4155
rect 295 4115 300 4155
rect 100 3290 300 4115
rect 100 3250 105 3290
rect 145 3250 155 3290
rect 195 3250 205 3290
rect 245 3250 255 3290
rect 295 3250 300 3290
rect 100 3240 300 3250
rect 100 3200 105 3240
rect 145 3200 155 3240
rect 195 3200 205 3240
rect 245 3200 255 3240
rect 295 3200 300 3240
rect 100 2550 300 3200
rect 100 2510 105 2550
rect 145 2510 155 2550
rect 195 2510 205 2550
rect 245 2510 255 2550
rect 295 2510 300 2550
rect 100 2500 300 2510
rect 100 2460 105 2500
rect 145 2460 155 2500
rect 195 2460 205 2500
rect 245 2460 255 2500
rect 295 2460 300 2500
rect 100 1790 300 2460
rect 100 1750 105 1790
rect 145 1750 155 1790
rect 195 1750 205 1790
rect 245 1750 255 1790
rect 295 1750 300 1790
rect 100 1740 300 1750
rect 100 1700 105 1740
rect 145 1700 155 1740
rect 195 1700 205 1740
rect 245 1700 255 1740
rect 295 1700 300 1740
rect 100 500 300 1700
rect 400 9580 600 22076
rect 400 9540 405 9580
rect 445 9540 455 9580
rect 495 9540 505 9580
rect 545 9540 555 9580
rect 595 9540 600 9580
rect 400 9520 600 9540
rect 400 9480 405 9520
rect 445 9480 455 9520
rect 495 9480 505 9520
rect 545 9480 555 9520
rect 595 9480 600 9520
rect 400 9230 600 9480
rect 400 9190 405 9230
rect 445 9190 455 9230
rect 495 9190 505 9230
rect 545 9190 555 9230
rect 595 9190 600 9230
rect 400 9180 600 9190
rect 400 9140 405 9180
rect 445 9140 455 9180
rect 495 9140 505 9180
rect 545 9140 555 9180
rect 595 9140 600 9180
rect 400 4055 600 9140
rect 400 4015 405 4055
rect 445 4015 455 4055
rect 495 4015 505 4055
rect 545 4015 555 4055
rect 595 4015 600 4055
rect 400 4005 600 4015
rect 400 3965 405 4005
rect 445 3965 455 4005
rect 495 3965 505 4005
rect 545 3965 555 4005
rect 595 3965 600 4005
rect 400 3880 600 3965
rect 400 3840 405 3880
rect 445 3840 455 3880
rect 495 3840 505 3880
rect 545 3840 555 3880
rect 595 3840 600 3880
rect 400 3830 600 3840
rect 400 3790 405 3830
rect 445 3790 455 3830
rect 495 3790 505 3830
rect 545 3790 555 3830
rect 595 3790 600 3830
rect 400 2700 600 3790
rect 400 2660 405 2700
rect 445 2660 455 2700
rect 495 2660 505 2700
rect 545 2660 555 2700
rect 595 2660 600 2700
rect 400 2650 600 2660
rect 400 2610 405 2650
rect 445 2610 455 2650
rect 495 2610 505 2650
rect 545 2610 555 2650
rect 595 2610 600 2650
rect 400 1400 600 2610
rect 400 1360 405 1400
rect 445 1360 455 1400
rect 495 1360 505 1400
rect 545 1360 555 1400
rect 595 1360 600 1400
rect 400 1350 600 1360
rect 400 1310 405 1350
rect 445 1310 455 1350
rect 495 1310 505 1350
rect 545 1310 555 1350
rect 595 1310 600 1350
rect 400 790 600 1310
rect 400 750 405 790
rect 445 750 455 790
rect 495 750 505 790
rect 545 750 555 790
rect 595 750 600 790
rect 400 740 600 750
rect 400 700 405 740
rect 445 700 455 740
rect 495 700 505 740
rect 545 700 555 740
rect 595 700 600 740
rect 400 500 600 700
rect 15185 670 15265 690
rect 15185 630 15205 670
rect 15245 630 15265 670
rect 15185 100 15265 630
rect 15181 0 15271 100
use pll_bgr_magic_3_flat  pll_bgr_magic_3_flat_0
timestamp 1756773826
transform 1 0 6155 0 -1 7865
box -2135 -7840 7050 7180
<< labels >>
flabel metal4 s 15181 0 15271 100 0 FreeSans 480 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 100 500 300 22076 1 FreeSans 200 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 400 500 600 22076 1 FreeSans 200 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal1 12150 1175 12150 1175 3 FreeSans 800 0 400 0 V_CONT
flabel metal2 12410 1540 12410 1540 3 FreeSans 800 0 400 0 ua1
<< properties >>
string FIXED_BBOX 0 0 16100 22576
<< end >>
