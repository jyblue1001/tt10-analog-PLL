magic
tech sky130A
magscale 1 2
timestamp 1756784274
<< nwell >>
rect -1570 12350 8880 12560
rect 9160 10760 11460 12610
rect -760 8620 4220 9860
rect 5500 9250 8720 9830
rect -1480 6630 160 6910
rect 420 6630 2060 6910
rect -1490 5630 2070 6310
rect 2370 5830 3140 6110
rect -2590 4470 140 4750
rect 440 4470 3170 4750
rect 5410 3530 8850 4840
<< pwell >>
rect 9160 12690 11270 13930
rect -1740 1427 -400 1580
rect -1740 393 -1587 1427
rect -553 393 -400 1427
rect -1740 240 -400 393
rect -380 1427 960 1580
rect -380 393 -227 1427
rect 807 393 960 1427
rect -380 240 960 393
rect 980 1427 2320 1580
rect 980 393 1133 1427
rect 2167 393 2320 1427
rect 980 240 2320 393
rect -1740 67 -400 220
rect -1740 -967 -1587 67
rect -553 -967 -400 67
rect -1740 -1120 -400 -967
rect -380 67 960 220
rect -380 -967 -227 67
rect 807 -967 960 67
rect -380 -1120 960 -967
rect 980 67 2320 220
rect 980 -967 1133 67
rect 2167 -967 2320 67
rect 980 -1120 2320 -967
rect -1740 -1293 -400 -1140
rect -1740 -2327 -1587 -1293
rect -553 -2327 -400 -1293
rect -1740 -2480 -400 -2327
rect -380 -1293 960 -1140
rect -380 -2327 -227 -1293
rect 807 -2327 960 -1293
rect -380 -2480 960 -2327
rect 980 -1293 2320 -1140
rect 980 -2327 1133 -1293
rect 2167 -2327 2320 -1293
rect 980 -2480 2320 -2327
rect 250 -2760 330 -2480
<< nbase >>
rect -1587 393 -553 1427
rect -227 393 807 1427
rect 1133 393 2167 1427
rect -1587 -967 -553 67
rect -227 -967 807 67
rect 1133 -967 2167 67
rect -1587 -2327 -553 -1293
rect -227 -2327 807 -1293
rect 1133 -2327 2167 -1293
<< nmos >>
rect 9380 13590 9410 13790
rect 9900 13590 9930 13790
rect 10420 13590 10450 13790
rect 11020 13590 11050 13790
rect 9380 13210 9410 13410
rect 9900 13210 9930 13410
rect 10420 13210 10450 13410
rect -1380 12740 -1350 12840
rect -1270 12740 -1240 12840
rect -1160 12740 -1130 12840
rect -1050 12740 -1020 12840
rect -800 12740 -770 12840
rect -690 12740 -660 12840
rect -350 12740 -320 12840
rect -240 12740 -210 12840
rect -130 12740 -100 12840
rect -20 12740 10 12840
rect 310 12740 340 12840
rect 420 12740 450 12840
rect 530 12740 560 12840
rect 640 12740 670 12840
rect 990 12740 1020 12840
rect 1100 12740 1130 12840
rect 1210 12740 1240 12840
rect 1320 12740 1350 12840
rect 1570 12740 1600 12840
rect 1680 12740 1710 12840
rect 2130 12740 2160 12840
rect 2490 12740 2520 12840
rect 2740 12740 2770 12840
rect 2850 12740 2880 12840
rect 2960 12740 2990 12840
rect 3070 12740 3100 12840
rect 3400 12740 3430 12840
rect 3510 12740 3540 12840
rect 3620 12740 3650 12840
rect 3950 12740 3980 12840
rect 4060 12740 4090 12840
rect 4170 12740 4200 12840
rect 4280 12740 4310 12840
rect 4610 12740 4640 12840
rect 4720 12740 4750 12840
rect 4830 12740 4860 12840
rect 5250 12830 5280 12930
rect 5360 12830 5390 12930
rect 5470 12830 5500 12930
rect 5580 12830 5610 12930
rect 5910 12830 5940 12930
rect 6020 12830 6050 12930
rect 6130 12830 6160 12930
rect 6550 12830 6580 12930
rect 6660 12830 6690 12930
rect 6770 12830 6800 12930
rect 6880 12830 6910 12930
rect 7210 12830 7240 12930
rect 7320 12830 7350 12930
rect 7430 12830 7460 12930
rect 7850 12830 7880 12930
rect 7960 12830 7990 12930
rect 8070 12830 8100 12930
rect 8180 12830 8210 12930
rect 8510 12830 8540 12930
rect 8620 12830 8650 12930
rect 8730 12830 8760 12930
rect 9380 12930 9410 13030
rect 9900 12930 9930 13030
rect 10420 12930 10450 13030
rect -560 10040 -530 10240
rect -450 10040 -420 10240
rect -40 10040 -10 10240
rect 70 10040 100 10240
rect 340 10040 370 10240
rect 450 10040 480 10240
rect 860 10040 890 10240
rect 970 10040 1000 10240
rect 1380 10040 1410 10240
rect 1490 10040 1520 10240
rect 1820 10040 1850 10240
rect 2150 10040 2180 10240
rect 2590 10040 2620 10240
rect 2980 10040 3010 10240
rect 3370 10040 3400 10240
rect 3660 10040 3690 10240
rect -560 8240 -530 8440
rect -450 8240 -420 8440
rect -40 8240 -10 8440
rect 70 8240 100 8440
rect 340 8240 370 8440
rect 450 8240 480 8440
rect 860 8240 890 8440
rect 970 8240 1000 8440
rect 1370 8240 1400 8440
rect 1700 8240 1730 8440
rect 2030 8240 2060 8440
rect 2590 8240 2620 8440
rect 2980 8240 3010 8440
rect 3370 8240 3400 8440
rect 3660 8240 3690 8440
rect 4050 8240 4080 8440
rect 5540 8290 5660 8690
rect 5760 8290 5880 8690
rect 5980 8290 6100 8690
rect 6200 8290 6320 8690
rect 6620 8290 6740 8690
rect 6840 8290 6960 8690
rect 7060 8290 7180 8690
rect 7280 8290 7400 8690
rect 7700 8290 7820 8690
rect 7920 8290 8040 8690
rect 8140 8290 8260 8690
rect 8360 8290 8480 8690
rect 5600 5810 5700 6060
rect 5800 5810 5900 6060
rect 6000 5810 6100 6060
rect 6200 5810 6300 6060
rect 6400 5810 6500 6060
rect 6600 5810 6700 6060
rect 6800 5810 6900 6060
rect 7000 5810 7100 6060
rect 7200 5810 7300 6060
rect 7400 5810 7500 6060
rect 5650 5270 5680 5370
rect 5780 5270 5810 5370
rect 5910 5270 5940 5370
rect 6040 5270 6070 5370
rect 6170 5270 6200 5370
rect 6300 5270 6330 5370
rect 6790 5270 6820 5370
rect 6920 5270 6950 5370
rect 7050 5270 7080 5370
rect 7180 5270 7210 5370
rect 7310 5270 7340 5370
rect 7440 5270 7470 5370
rect 7930 5270 7960 5370
rect 8060 5270 8090 5370
rect 8190 5270 8220 5370
rect 8320 5270 8350 5370
rect 8450 5270 8480 5370
rect 8580 5270 8610 5370
rect -1550 3670 -1510 3770
rect -1430 3670 -1390 3770
rect -1310 3670 -1270 3770
rect -1190 3670 -1150 3770
rect -1070 3670 -1030 3770
rect -950 3670 -910 3770
rect -830 3670 -790 3770
rect -710 3670 -670 3770
rect -590 3670 -550 3770
rect -470 3670 -430 3770
rect 1010 3670 1050 3770
rect 1130 3670 1170 3770
rect 1250 3670 1290 3770
rect 1370 3670 1410 3770
rect 1490 3670 1530 3770
rect 1610 3670 1650 3770
rect 1730 3670 1770 3770
rect 1850 3670 1890 3770
rect 1970 3670 2010 3770
rect 2090 3670 2130 3770
rect -2170 2660 -1170 3160
rect -930 2660 70 3160
rect 510 2660 1510 3160
rect 1750 2660 2750 3160
rect -1750 2050 250 2250
rect 330 2050 2330 2250
<< pmos >>
rect -1220 12420 -1190 12520
rect -800 12420 -770 12520
rect -690 12420 -660 12520
rect -130 12420 -100 12520
rect -20 12420 10 12520
rect 310 12420 340 12520
rect 420 12420 450 12520
rect 530 12420 560 12520
rect 1150 12420 1180 12520
rect 1570 12420 1600 12520
rect 1680 12420 1710 12520
rect 2020 12420 2050 12520
rect 2130 12420 2160 12520
rect 2380 12420 2410 12520
rect 2490 12420 2520 12520
rect 2960 12420 2990 12520
rect 3070 12420 3100 12520
rect 3400 12420 3430 12520
rect 3510 12420 3540 12520
rect 4020 12420 4050 12520
rect 4360 12420 4390 12520
rect 4470 12420 4500 12520
rect 4720 12420 4750 12520
rect 4830 12420 4860 12520
rect 5320 12420 5350 12520
rect 5660 12420 5690 12520
rect 5770 12420 5800 12520
rect 6020 12420 6050 12520
rect 6130 12420 6160 12520
rect 6620 12420 6650 12520
rect 6960 12420 6990 12520
rect 7070 12420 7100 12520
rect 7320 12420 7350 12520
rect 7430 12420 7460 12520
rect 7920 12420 7950 12520
rect 8260 12420 8290 12520
rect 8370 12420 8400 12520
rect 8620 12420 8650 12520
rect 8730 12420 8760 12520
rect 9380 12170 9410 12370
rect 9900 12170 9930 12370
rect 10420 12170 10450 12370
rect 9380 11590 9410 11990
rect 9900 11590 9930 11990
rect 10420 11590 10450 11990
rect 9380 10900 9680 11300
rect 9900 10900 10200 11300
rect 10420 10900 10720 11300
rect 10940 10900 11240 11300
rect -560 9420 -530 9820
rect -450 9420 -420 9820
rect -40 9420 -10 9820
rect 70 9420 100 9820
rect 340 9420 370 9820
rect 450 9420 480 9820
rect 860 9420 890 9820
rect 970 9420 1000 9820
rect 1380 9420 1410 9820
rect 1490 9420 1520 9820
rect 1820 9420 1850 9820
rect 2150 9420 2180 9820
rect 2590 9420 2620 9820
rect 2980 9420 3010 9820
rect 3370 9420 3400 9820
rect 3660 9420 3690 9820
rect 4050 9420 4080 9820
rect 5740 9390 5860 9790
rect 5960 9390 6080 9790
rect 6180 9390 6300 9790
rect 6400 9390 6520 9790
rect 6620 9390 6740 9790
rect 6840 9390 6960 9790
rect 7260 9390 7380 9790
rect 7480 9390 7600 9790
rect 7700 9390 7820 9790
rect 7920 9390 8040 9790
rect 8140 9390 8260 9790
rect 8360 9390 8480 9790
rect -560 8660 -530 9060
rect -450 8660 -420 9060
rect -40 8660 -10 9060
rect 70 8660 100 9060
rect 340 8660 370 9060
rect 450 8660 480 9060
rect 860 8660 890 9060
rect 970 8660 1000 9060
rect 1370 8660 1400 9060
rect 1700 8660 1730 9060
rect 2030 8660 2060 9060
rect 2590 8660 2620 9060
rect 2980 8660 3010 9060
rect 3370 8660 3400 9060
rect 3660 8660 3690 9060
rect -1280 6670 -1250 6870
rect -1170 6670 -1140 6870
rect -1060 6670 -1030 6870
rect -950 6670 -920 6870
rect -840 6670 -810 6870
rect -730 6670 -700 6870
rect -620 6670 -590 6870
rect -510 6670 -480 6870
rect -400 6670 -370 6870
rect -290 6670 -260 6870
rect -180 6670 -150 6870
rect -70 6670 -40 6870
rect 620 6670 650 6870
rect 730 6670 760 6870
rect 840 6670 870 6870
rect 950 6670 980 6870
rect 1060 6670 1090 6870
rect 1170 6670 1200 6870
rect 1280 6670 1310 6870
rect 1390 6670 1420 6870
rect 1500 6670 1530 6870
rect 1610 6670 1640 6870
rect 1720 6670 1750 6870
rect 1830 6670 1860 6870
rect -1290 5670 -1190 6270
rect -1110 5670 -1010 6270
rect -930 5670 -830 6270
rect -750 5670 -650 6270
rect -570 5670 -470 6270
rect -390 5670 -290 6270
rect -210 5670 -110 6270
rect -30 5670 70 6270
rect 150 5670 250 6270
rect 330 5670 430 6270
rect 510 5670 610 6270
rect 690 5670 790 6270
rect 870 5670 970 6270
rect 1050 5670 1150 6270
rect 1230 5670 1330 6270
rect 1410 5670 1510 6270
rect 1590 5670 1690 6270
rect 1770 5670 1870 6270
rect 2580 5870 2610 6070
rect 2690 5870 2720 6070
rect 2800 5870 2830 6070
rect 2910 5870 2940 6070
rect -2390 4510 -2350 4710
rect -2270 4510 -2230 4710
rect -2150 4510 -2110 4710
rect -2030 4510 -1990 4710
rect -1910 4510 -1870 4710
rect -1790 4510 -1750 4710
rect -1670 4510 -1630 4710
rect -1550 4510 -1510 4710
rect -1430 4510 -1390 4710
rect -1310 4510 -1270 4710
rect -1190 4510 -1150 4710
rect -1070 4510 -1030 4710
rect -950 4510 -910 4710
rect -830 4510 -790 4710
rect -710 4510 -670 4710
rect -590 4510 -550 4710
rect -470 4510 -430 4710
rect -350 4510 -310 4710
rect -230 4510 -190 4710
rect -110 4510 -70 4710
rect 650 4510 690 4710
rect 770 4510 810 4710
rect 890 4510 930 4710
rect 1010 4510 1050 4710
rect 1130 4510 1170 4710
rect 1250 4510 1290 4710
rect 1370 4510 1410 4710
rect 1490 4510 1530 4710
rect 1610 4510 1650 4710
rect 1730 4510 1770 4710
rect 1850 4510 1890 4710
rect 1970 4510 2010 4710
rect 2090 4510 2130 4710
rect 2210 4510 2250 4710
rect 2330 4510 2370 4710
rect 2450 4510 2490 4710
rect 2570 4510 2610 4710
rect 2690 4510 2730 4710
rect 2810 4510 2850 4710
rect 2930 4510 2970 4710
rect 5650 4590 5680 4790
rect 5780 4590 5810 4790
rect 5910 4590 5940 4790
rect 6040 4590 6070 4790
rect 6170 4590 6200 4790
rect 6300 4590 6330 4790
rect 6790 4590 6820 4790
rect 6920 4590 6950 4790
rect 7050 4590 7080 4790
rect 7180 4590 7210 4790
rect 7310 4590 7340 4790
rect 7440 4590 7470 4790
rect 7930 4590 7960 4790
rect 8060 4590 8090 4790
rect 8190 4590 8220 4790
rect 8320 4590 8350 4790
rect 8450 4590 8480 4790
rect 8580 4590 8610 4790
rect 5720 3640 5820 4140
rect 5920 3640 6020 4140
rect 6120 3640 6220 4140
rect 6320 3640 6420 4140
rect 6520 3640 6620 4140
rect 6720 3640 6820 4140
rect 6920 3640 7020 4140
rect 7120 3640 7220 4140
rect 7320 3640 7420 4140
rect 7520 3640 7620 4140
<< ndiff >>
rect 9300 13760 9380 13790
rect 9300 13720 9320 13760
rect 9360 13720 9380 13760
rect 9300 13660 9380 13720
rect 9300 13620 9320 13660
rect 9360 13620 9380 13660
rect 9300 13590 9380 13620
rect 9410 13760 9490 13790
rect 9410 13720 9430 13760
rect 9470 13720 9490 13760
rect 9410 13660 9490 13720
rect 9410 13620 9430 13660
rect 9470 13620 9490 13660
rect 9410 13590 9490 13620
rect 9820 13760 9900 13790
rect 9820 13720 9840 13760
rect 9880 13720 9900 13760
rect 9820 13660 9900 13720
rect 9820 13620 9840 13660
rect 9880 13620 9900 13660
rect 9820 13590 9900 13620
rect 9930 13760 10010 13790
rect 9930 13720 9950 13760
rect 9990 13720 10010 13760
rect 9930 13660 10010 13720
rect 9930 13620 9950 13660
rect 9990 13620 10010 13660
rect 9930 13590 10010 13620
rect 10340 13760 10420 13790
rect 10340 13720 10360 13760
rect 10400 13720 10420 13760
rect 10340 13660 10420 13720
rect 10340 13620 10360 13660
rect 10400 13620 10420 13660
rect 10340 13590 10420 13620
rect 10450 13760 10530 13790
rect 10450 13720 10470 13760
rect 10510 13720 10530 13760
rect 10450 13660 10530 13720
rect 10450 13620 10470 13660
rect 10510 13620 10530 13660
rect 10450 13590 10530 13620
rect 10940 13760 11020 13790
rect 10940 13720 10960 13760
rect 11000 13720 11020 13760
rect 10940 13660 11020 13720
rect 10940 13620 10960 13660
rect 11000 13620 11020 13660
rect 10940 13590 11020 13620
rect 11050 13760 11130 13790
rect 11050 13720 11070 13760
rect 11110 13720 11130 13760
rect 11050 13660 11130 13720
rect 11050 13620 11070 13660
rect 11110 13620 11130 13660
rect 11050 13590 11130 13620
rect 9300 13380 9380 13410
rect 9300 13340 9320 13380
rect 9360 13340 9380 13380
rect 9300 13280 9380 13340
rect 9300 13240 9320 13280
rect 9360 13240 9380 13280
rect 9300 13210 9380 13240
rect 9410 13380 9490 13410
rect 9410 13340 9430 13380
rect 9470 13340 9490 13380
rect 9410 13280 9490 13340
rect 9410 13240 9430 13280
rect 9470 13240 9490 13280
rect 9410 13210 9490 13240
rect 9820 13380 9900 13410
rect 9820 13340 9840 13380
rect 9880 13340 9900 13380
rect 9820 13280 9900 13340
rect 9820 13240 9840 13280
rect 9880 13240 9900 13280
rect 9820 13210 9900 13240
rect 9930 13380 10010 13410
rect 9930 13340 9950 13380
rect 9990 13340 10010 13380
rect 9930 13280 10010 13340
rect 9930 13240 9950 13280
rect 9990 13240 10010 13280
rect 9930 13210 10010 13240
rect 10340 13380 10420 13410
rect 10340 13340 10360 13380
rect 10400 13340 10420 13380
rect 10340 13280 10420 13340
rect 10340 13240 10360 13280
rect 10400 13240 10420 13280
rect 10340 13210 10420 13240
rect 10450 13380 10530 13410
rect 10450 13340 10470 13380
rect 10510 13340 10530 13380
rect 10450 13280 10530 13340
rect 10450 13240 10470 13280
rect 10510 13240 10530 13280
rect 10450 13210 10530 13240
rect -1460 12810 -1380 12840
rect -1460 12770 -1440 12810
rect -1400 12770 -1380 12810
rect -1460 12740 -1380 12770
rect -1350 12810 -1270 12840
rect -1350 12770 -1330 12810
rect -1290 12770 -1270 12810
rect -1350 12740 -1270 12770
rect -1240 12810 -1160 12840
rect -1240 12770 -1220 12810
rect -1180 12770 -1160 12810
rect -1240 12740 -1160 12770
rect -1130 12810 -1050 12840
rect -1130 12770 -1110 12810
rect -1070 12770 -1050 12810
rect -1130 12740 -1050 12770
rect -1020 12810 -940 12840
rect -1020 12770 -1000 12810
rect -960 12770 -940 12810
rect -1020 12740 -940 12770
rect -880 12810 -800 12840
rect -880 12770 -860 12810
rect -820 12770 -800 12810
rect -880 12740 -800 12770
rect -770 12810 -690 12840
rect -770 12770 -750 12810
rect -710 12770 -690 12810
rect -770 12740 -690 12770
rect -660 12810 -580 12840
rect -660 12770 -640 12810
rect -600 12770 -580 12810
rect -660 12740 -580 12770
rect -430 12810 -350 12840
rect -430 12770 -410 12810
rect -370 12770 -350 12810
rect -430 12740 -350 12770
rect -320 12810 -240 12840
rect -320 12770 -300 12810
rect -260 12770 -240 12810
rect -320 12740 -240 12770
rect -210 12810 -130 12840
rect -210 12770 -190 12810
rect -150 12770 -130 12810
rect -210 12740 -130 12770
rect -100 12810 -20 12840
rect -100 12770 -80 12810
rect -40 12770 -20 12810
rect -100 12740 -20 12770
rect 10 12810 90 12840
rect 10 12770 30 12810
rect 70 12770 90 12810
rect 10 12740 90 12770
rect 230 12810 310 12840
rect 230 12770 250 12810
rect 290 12770 310 12810
rect 230 12740 310 12770
rect 340 12810 420 12840
rect 340 12770 360 12810
rect 400 12770 420 12810
rect 340 12740 420 12770
rect 450 12810 530 12840
rect 450 12770 470 12810
rect 510 12770 530 12810
rect 450 12740 530 12770
rect 560 12810 640 12840
rect 560 12770 580 12810
rect 620 12770 640 12810
rect 560 12740 640 12770
rect 670 12810 750 12840
rect 670 12770 690 12810
rect 730 12770 750 12810
rect 670 12740 750 12770
rect 910 12810 990 12840
rect 910 12770 930 12810
rect 970 12770 990 12810
rect 910 12740 990 12770
rect 1020 12810 1100 12840
rect 1020 12770 1040 12810
rect 1080 12770 1100 12810
rect 1020 12740 1100 12770
rect 1130 12810 1210 12840
rect 1130 12770 1150 12810
rect 1190 12770 1210 12810
rect 1130 12740 1210 12770
rect 1240 12810 1320 12840
rect 1240 12770 1260 12810
rect 1300 12770 1320 12810
rect 1240 12740 1320 12770
rect 1350 12810 1430 12840
rect 1350 12770 1370 12810
rect 1410 12770 1430 12810
rect 1350 12740 1430 12770
rect 1490 12810 1570 12840
rect 1490 12770 1510 12810
rect 1550 12770 1570 12810
rect 1490 12740 1570 12770
rect 1600 12810 1680 12840
rect 1600 12770 1620 12810
rect 1660 12770 1680 12810
rect 1600 12740 1680 12770
rect 1710 12810 1790 12840
rect 1710 12770 1730 12810
rect 1770 12770 1790 12810
rect 1710 12740 1790 12770
rect 2050 12810 2130 12840
rect 2050 12770 2070 12810
rect 2110 12770 2130 12810
rect 2050 12740 2130 12770
rect 2160 12810 2240 12840
rect 2160 12770 2180 12810
rect 2220 12770 2240 12810
rect 2160 12740 2240 12770
rect 2410 12810 2490 12840
rect 2410 12770 2430 12810
rect 2470 12770 2490 12810
rect 2410 12740 2490 12770
rect 2520 12810 2600 12840
rect 2520 12770 2540 12810
rect 2580 12770 2600 12810
rect 2520 12740 2600 12770
rect 2660 12810 2740 12840
rect 2660 12770 2680 12810
rect 2720 12770 2740 12810
rect 2660 12740 2740 12770
rect 2770 12810 2850 12840
rect 2770 12770 2790 12810
rect 2830 12770 2850 12810
rect 2770 12740 2850 12770
rect 2880 12810 2960 12840
rect 2880 12770 2900 12810
rect 2940 12770 2960 12810
rect 2880 12740 2960 12770
rect 2990 12810 3070 12840
rect 2990 12770 3010 12810
rect 3050 12770 3070 12810
rect 2990 12740 3070 12770
rect 3100 12810 3180 12840
rect 3100 12770 3120 12810
rect 3160 12770 3180 12810
rect 3100 12740 3180 12770
rect 3320 12810 3400 12840
rect 3320 12770 3340 12810
rect 3380 12770 3400 12810
rect 3320 12740 3400 12770
rect 3430 12810 3510 12840
rect 3430 12770 3450 12810
rect 3490 12770 3510 12810
rect 3430 12740 3510 12770
rect 3540 12810 3620 12840
rect 3540 12770 3560 12810
rect 3600 12770 3620 12810
rect 3540 12740 3620 12770
rect 3650 12810 3730 12840
rect 3650 12770 3670 12810
rect 3710 12770 3730 12810
rect 3650 12740 3730 12770
rect 3870 12810 3950 12840
rect 3870 12770 3890 12810
rect 3930 12770 3950 12810
rect 3870 12740 3950 12770
rect 3980 12810 4060 12840
rect 3980 12770 4000 12810
rect 4040 12770 4060 12810
rect 3980 12740 4060 12770
rect 4090 12810 4170 12840
rect 4090 12770 4110 12810
rect 4150 12770 4170 12810
rect 4090 12740 4170 12770
rect 4200 12810 4280 12840
rect 4200 12770 4220 12810
rect 4260 12770 4280 12810
rect 4200 12740 4280 12770
rect 4310 12810 4390 12840
rect 4310 12770 4330 12810
rect 4370 12770 4390 12810
rect 4310 12740 4390 12770
rect 4530 12810 4610 12840
rect 4530 12770 4550 12810
rect 4590 12770 4610 12810
rect 4530 12740 4610 12770
rect 4640 12810 4720 12840
rect 4640 12770 4660 12810
rect 4700 12770 4720 12810
rect 4640 12740 4720 12770
rect 4750 12810 4830 12840
rect 4750 12770 4770 12810
rect 4810 12770 4830 12810
rect 4750 12740 4830 12770
rect 4860 12810 4940 12840
rect 5170 12900 5250 12930
rect 5170 12860 5190 12900
rect 5230 12860 5250 12900
rect 5170 12830 5250 12860
rect 5280 12900 5360 12930
rect 5280 12860 5300 12900
rect 5340 12860 5360 12900
rect 5280 12830 5360 12860
rect 5390 12900 5470 12930
rect 5390 12860 5410 12900
rect 5450 12860 5470 12900
rect 5390 12830 5470 12860
rect 5500 12900 5580 12930
rect 5500 12860 5520 12900
rect 5560 12860 5580 12900
rect 5500 12830 5580 12860
rect 5610 12900 5690 12930
rect 5610 12860 5630 12900
rect 5670 12860 5690 12900
rect 5610 12830 5690 12860
rect 5830 12900 5910 12930
rect 5830 12860 5850 12900
rect 5890 12860 5910 12900
rect 5830 12830 5910 12860
rect 5940 12900 6020 12930
rect 5940 12860 5960 12900
rect 6000 12860 6020 12900
rect 5940 12830 6020 12860
rect 6050 12900 6130 12930
rect 6050 12860 6070 12900
rect 6110 12860 6130 12900
rect 6050 12830 6130 12860
rect 6160 12900 6240 12930
rect 6160 12860 6180 12900
rect 6220 12860 6240 12900
rect 6160 12830 6240 12860
rect 6470 12900 6550 12930
rect 6470 12860 6490 12900
rect 6530 12860 6550 12900
rect 6470 12830 6550 12860
rect 6580 12900 6660 12930
rect 6580 12860 6600 12900
rect 6640 12860 6660 12900
rect 6580 12830 6660 12860
rect 6690 12900 6770 12930
rect 6690 12860 6710 12900
rect 6750 12860 6770 12900
rect 6690 12830 6770 12860
rect 6800 12900 6880 12930
rect 6800 12860 6820 12900
rect 6860 12860 6880 12900
rect 6800 12830 6880 12860
rect 6910 12900 6990 12930
rect 6910 12860 6930 12900
rect 6970 12860 6990 12900
rect 6910 12830 6990 12860
rect 7130 12900 7210 12930
rect 7130 12860 7150 12900
rect 7190 12860 7210 12900
rect 7130 12830 7210 12860
rect 7240 12900 7320 12930
rect 7240 12860 7260 12900
rect 7300 12860 7320 12900
rect 7240 12830 7320 12860
rect 7350 12900 7430 12930
rect 7350 12860 7370 12900
rect 7410 12860 7430 12900
rect 7350 12830 7430 12860
rect 7460 12900 7540 12930
rect 7460 12860 7480 12900
rect 7520 12860 7540 12900
rect 7460 12830 7540 12860
rect 7770 12900 7850 12930
rect 7770 12860 7790 12900
rect 7830 12860 7850 12900
rect 7770 12830 7850 12860
rect 7880 12900 7960 12930
rect 7880 12860 7900 12900
rect 7940 12860 7960 12900
rect 7880 12830 7960 12860
rect 7990 12900 8070 12930
rect 7990 12860 8010 12900
rect 8050 12860 8070 12900
rect 7990 12830 8070 12860
rect 8100 12900 8180 12930
rect 8100 12860 8120 12900
rect 8160 12860 8180 12900
rect 8100 12830 8180 12860
rect 8210 12900 8290 12930
rect 8210 12860 8230 12900
rect 8270 12860 8290 12900
rect 8210 12830 8290 12860
rect 8430 12900 8510 12930
rect 8430 12860 8450 12900
rect 8490 12860 8510 12900
rect 8430 12830 8510 12860
rect 8540 12900 8620 12930
rect 8540 12860 8560 12900
rect 8600 12860 8620 12900
rect 8540 12830 8620 12860
rect 8650 12900 8730 12930
rect 8650 12860 8670 12900
rect 8710 12860 8730 12900
rect 8650 12830 8730 12860
rect 8760 12900 8840 12930
rect 8760 12860 8780 12900
rect 8820 12860 8840 12900
rect 8760 12830 8840 12860
rect 4860 12770 4880 12810
rect 4920 12770 4940 12810
rect 4860 12740 4940 12770
rect 9300 13000 9380 13030
rect 9300 12960 9320 13000
rect 9360 12960 9380 13000
rect 9300 12930 9380 12960
rect 9410 13000 9490 13030
rect 9410 12960 9430 13000
rect 9470 12960 9490 13000
rect 9410 12930 9490 12960
rect 9820 13000 9900 13030
rect 9820 12960 9840 13000
rect 9880 12960 9900 13000
rect 9820 12930 9900 12960
rect 9930 13000 10010 13030
rect 9930 12960 9950 13000
rect 9990 12960 10010 13000
rect 9930 12930 10010 12960
rect 10340 13000 10420 13030
rect 10340 12960 10360 13000
rect 10400 12960 10420 13000
rect 10340 12930 10420 12960
rect 10450 13000 10530 13030
rect 10450 12960 10470 13000
rect 10510 12960 10530 13000
rect 10450 12930 10530 12960
rect -640 10210 -560 10240
rect -640 10170 -620 10210
rect -580 10170 -560 10210
rect -640 10110 -560 10170
rect -640 10070 -620 10110
rect -580 10070 -560 10110
rect -640 10040 -560 10070
rect -530 10210 -450 10240
rect -530 10170 -510 10210
rect -470 10170 -450 10210
rect -530 10110 -450 10170
rect -530 10070 -510 10110
rect -470 10070 -450 10110
rect -530 10040 -450 10070
rect -420 10210 -340 10240
rect -420 10170 -400 10210
rect -360 10170 -340 10210
rect -420 10110 -340 10170
rect -420 10070 -400 10110
rect -360 10070 -340 10110
rect -420 10040 -340 10070
rect -120 10210 -40 10240
rect -120 10170 -100 10210
rect -60 10170 -40 10210
rect -120 10110 -40 10170
rect -120 10070 -100 10110
rect -60 10070 -40 10110
rect -120 10040 -40 10070
rect -10 10210 70 10240
rect -10 10170 10 10210
rect 50 10170 70 10210
rect -10 10110 70 10170
rect -10 10070 10 10110
rect 50 10070 70 10110
rect -10 10040 70 10070
rect 100 10210 180 10240
rect 260 10210 340 10240
rect 100 10170 120 10210
rect 160 10170 180 10210
rect 260 10170 280 10210
rect 320 10170 340 10210
rect 100 10110 180 10170
rect 260 10110 340 10170
rect 100 10070 120 10110
rect 160 10070 180 10110
rect 260 10070 280 10110
rect 320 10070 340 10110
rect 100 10040 180 10070
rect 260 10040 340 10070
rect 370 10210 450 10240
rect 370 10170 390 10210
rect 430 10170 450 10210
rect 370 10110 450 10170
rect 370 10070 390 10110
rect 430 10070 450 10110
rect 370 10040 450 10070
rect 480 10210 560 10240
rect 480 10170 500 10210
rect 540 10170 560 10210
rect 480 10110 560 10170
rect 480 10070 500 10110
rect 540 10070 560 10110
rect 480 10040 560 10070
rect 780 10210 860 10240
rect 780 10170 800 10210
rect 840 10170 860 10210
rect 780 10110 860 10170
rect 780 10070 800 10110
rect 840 10070 860 10110
rect 780 10040 860 10070
rect 890 10210 970 10240
rect 890 10170 910 10210
rect 950 10170 970 10210
rect 890 10110 970 10170
rect 890 10070 910 10110
rect 950 10070 970 10110
rect 890 10040 970 10070
rect 1000 10210 1080 10240
rect 1000 10170 1020 10210
rect 1060 10170 1080 10210
rect 1000 10110 1080 10170
rect 1000 10070 1020 10110
rect 1060 10070 1080 10110
rect 1000 10040 1080 10070
rect 1300 10210 1380 10240
rect 1300 10170 1320 10210
rect 1360 10170 1380 10210
rect 1300 10110 1380 10170
rect 1300 10070 1320 10110
rect 1360 10070 1380 10110
rect 1300 10040 1380 10070
rect 1410 10210 1490 10240
rect 1410 10170 1430 10210
rect 1470 10170 1490 10210
rect 1410 10110 1490 10170
rect 1410 10070 1430 10110
rect 1470 10070 1490 10110
rect 1410 10040 1490 10070
rect 1520 10210 1600 10240
rect 1520 10170 1540 10210
rect 1580 10170 1600 10210
rect 1520 10110 1600 10170
rect 1520 10070 1540 10110
rect 1580 10070 1600 10110
rect 1520 10040 1600 10070
rect 1740 10210 1820 10240
rect 1740 10170 1760 10210
rect 1800 10170 1820 10210
rect 1740 10110 1820 10170
rect 1740 10070 1760 10110
rect 1800 10070 1820 10110
rect 1740 10040 1820 10070
rect 1850 10210 1930 10240
rect 1850 10170 1870 10210
rect 1910 10170 1930 10210
rect 1850 10110 1930 10170
rect 1850 10070 1870 10110
rect 1910 10070 1930 10110
rect 1850 10040 1930 10070
rect 2070 10210 2150 10240
rect 2070 10170 2090 10210
rect 2130 10170 2150 10210
rect 2070 10110 2150 10170
rect 2070 10070 2090 10110
rect 2130 10070 2150 10110
rect 2070 10040 2150 10070
rect 2180 10210 2260 10240
rect 2180 10170 2200 10210
rect 2240 10170 2260 10210
rect 2180 10110 2260 10170
rect 2180 10070 2200 10110
rect 2240 10070 2260 10110
rect 2180 10040 2260 10070
rect 2490 10210 2590 10240
rect 2490 10170 2520 10210
rect 2560 10170 2590 10210
rect 2490 10110 2590 10170
rect 2490 10070 2520 10110
rect 2560 10070 2590 10110
rect 2490 10040 2590 10070
rect 2620 10210 2720 10240
rect 2620 10170 2650 10210
rect 2690 10170 2720 10210
rect 2620 10110 2720 10170
rect 2620 10070 2650 10110
rect 2690 10070 2720 10110
rect 2620 10040 2720 10070
rect 2880 10210 2980 10240
rect 2880 10170 2910 10210
rect 2950 10170 2980 10210
rect 2880 10110 2980 10170
rect 2880 10070 2910 10110
rect 2950 10070 2980 10110
rect 2880 10040 2980 10070
rect 3010 10210 3110 10240
rect 3010 10170 3040 10210
rect 3080 10170 3110 10210
rect 3010 10110 3110 10170
rect 3010 10070 3040 10110
rect 3080 10070 3110 10110
rect 3010 10040 3110 10070
rect 3270 10210 3370 10240
rect 3270 10170 3300 10210
rect 3340 10170 3370 10210
rect 3270 10110 3370 10170
rect 3270 10070 3300 10110
rect 3340 10070 3370 10110
rect 3270 10040 3370 10070
rect 3400 10210 3500 10240
rect 3400 10170 3430 10210
rect 3470 10170 3500 10210
rect 3400 10110 3500 10170
rect 3400 10070 3430 10110
rect 3470 10070 3500 10110
rect 3400 10040 3500 10070
rect 3560 10210 3660 10240
rect 3560 10170 3590 10210
rect 3630 10170 3660 10210
rect 3560 10110 3660 10170
rect 3560 10070 3590 10110
rect 3630 10070 3660 10110
rect 3560 10040 3660 10070
rect 3690 10210 3790 10240
rect 3690 10170 3720 10210
rect 3760 10170 3790 10210
rect 3690 10110 3790 10170
rect 3690 10070 3720 10110
rect 3760 10070 3790 10110
rect 3690 10040 3790 10070
rect 5440 8660 5540 8690
rect 5440 8620 5470 8660
rect 5510 8620 5540 8660
rect 5440 8560 5540 8620
rect 5440 8520 5470 8560
rect 5510 8520 5540 8560
rect 5440 8460 5540 8520
rect -640 8410 -560 8440
rect -640 8370 -620 8410
rect -580 8370 -560 8410
rect -640 8310 -560 8370
rect -640 8270 -620 8310
rect -580 8270 -560 8310
rect -640 8240 -560 8270
rect -530 8410 -450 8440
rect -530 8370 -510 8410
rect -470 8370 -450 8410
rect -530 8310 -450 8370
rect -530 8270 -510 8310
rect -470 8270 -450 8310
rect -530 8240 -450 8270
rect -420 8410 -340 8440
rect -420 8370 -400 8410
rect -360 8370 -340 8410
rect -420 8310 -340 8370
rect -420 8270 -400 8310
rect -360 8270 -340 8310
rect -420 8240 -340 8270
rect -120 8410 -40 8440
rect -120 8370 -100 8410
rect -60 8370 -40 8410
rect -120 8310 -40 8370
rect -120 8270 -100 8310
rect -60 8270 -40 8310
rect -120 8240 -40 8270
rect -10 8410 70 8440
rect -10 8370 10 8410
rect 50 8370 70 8410
rect -10 8310 70 8370
rect -10 8270 10 8310
rect 50 8270 70 8310
rect -10 8240 70 8270
rect 100 8410 180 8440
rect 260 8410 340 8440
rect 100 8370 120 8410
rect 160 8370 180 8410
rect 260 8370 280 8410
rect 320 8370 340 8410
rect 100 8310 180 8370
rect 260 8310 340 8370
rect 100 8270 120 8310
rect 160 8270 180 8310
rect 260 8270 280 8310
rect 320 8270 340 8310
rect 100 8240 180 8270
rect 260 8240 340 8270
rect 370 8410 450 8440
rect 370 8370 390 8410
rect 430 8370 450 8410
rect 370 8310 450 8370
rect 370 8270 390 8310
rect 430 8270 450 8310
rect 370 8240 450 8270
rect 480 8410 560 8440
rect 480 8370 500 8410
rect 540 8370 560 8410
rect 480 8310 560 8370
rect 480 8270 500 8310
rect 540 8270 560 8310
rect 480 8240 560 8270
rect 780 8410 860 8440
rect 780 8370 800 8410
rect 840 8370 860 8410
rect 780 8310 860 8370
rect 780 8270 800 8310
rect 840 8270 860 8310
rect 780 8240 860 8270
rect 890 8410 970 8440
rect 890 8370 910 8410
rect 950 8370 970 8410
rect 890 8310 970 8370
rect 890 8270 910 8310
rect 950 8270 970 8310
rect 890 8240 970 8270
rect 1000 8410 1080 8440
rect 1000 8370 1020 8410
rect 1060 8370 1080 8410
rect 1000 8310 1080 8370
rect 1000 8270 1020 8310
rect 1060 8270 1080 8310
rect 1000 8240 1080 8270
rect 1290 8410 1370 8440
rect 1290 8370 1310 8410
rect 1350 8370 1370 8410
rect 1290 8310 1370 8370
rect 1290 8270 1310 8310
rect 1350 8270 1370 8310
rect 1290 8240 1370 8270
rect 1400 8410 1480 8440
rect 1400 8370 1420 8410
rect 1460 8370 1480 8410
rect 1400 8310 1480 8370
rect 1400 8270 1420 8310
rect 1460 8270 1480 8310
rect 1400 8240 1480 8270
rect 1620 8410 1700 8440
rect 1620 8370 1640 8410
rect 1680 8370 1700 8410
rect 1620 8310 1700 8370
rect 1620 8270 1640 8310
rect 1680 8270 1700 8310
rect 1620 8240 1700 8270
rect 1730 8410 1810 8440
rect 1730 8370 1750 8410
rect 1790 8370 1810 8410
rect 1730 8310 1810 8370
rect 1730 8270 1750 8310
rect 1790 8270 1810 8310
rect 1730 8240 1810 8270
rect 1950 8410 2030 8440
rect 1950 8370 1970 8410
rect 2010 8370 2030 8410
rect 1950 8310 2030 8370
rect 1950 8270 1970 8310
rect 2010 8270 2030 8310
rect 1950 8240 2030 8270
rect 2060 8410 2140 8440
rect 2060 8370 2080 8410
rect 2120 8370 2140 8410
rect 2060 8310 2140 8370
rect 2060 8270 2080 8310
rect 2120 8270 2140 8310
rect 2060 8240 2140 8270
rect 2490 8410 2590 8440
rect 2490 8370 2520 8410
rect 2560 8370 2590 8410
rect 2490 8310 2590 8370
rect 2490 8270 2520 8310
rect 2560 8270 2590 8310
rect 2490 8240 2590 8270
rect 2620 8410 2720 8440
rect 2620 8370 2650 8410
rect 2690 8370 2720 8410
rect 2620 8310 2720 8370
rect 2620 8270 2650 8310
rect 2690 8270 2720 8310
rect 2620 8240 2720 8270
rect 2880 8410 2980 8440
rect 2880 8370 2910 8410
rect 2950 8370 2980 8410
rect 2880 8310 2980 8370
rect 2880 8270 2910 8310
rect 2950 8270 2980 8310
rect 2880 8240 2980 8270
rect 3010 8410 3110 8440
rect 3010 8370 3040 8410
rect 3080 8370 3110 8410
rect 3010 8310 3110 8370
rect 3010 8270 3040 8310
rect 3080 8270 3110 8310
rect 3010 8240 3110 8270
rect 3270 8410 3370 8440
rect 3270 8370 3300 8410
rect 3340 8370 3370 8410
rect 3270 8310 3370 8370
rect 3270 8270 3300 8310
rect 3340 8270 3370 8310
rect 3270 8240 3370 8270
rect 3400 8410 3500 8440
rect 3400 8370 3430 8410
rect 3470 8370 3500 8410
rect 3400 8310 3500 8370
rect 3400 8270 3430 8310
rect 3470 8270 3500 8310
rect 3400 8240 3500 8270
rect 3560 8410 3660 8440
rect 3560 8370 3590 8410
rect 3630 8370 3660 8410
rect 3560 8310 3660 8370
rect 3560 8270 3590 8310
rect 3630 8270 3660 8310
rect 3560 8240 3660 8270
rect 3690 8410 3790 8440
rect 3690 8370 3720 8410
rect 3760 8370 3790 8410
rect 3690 8310 3790 8370
rect 3690 8270 3720 8310
rect 3760 8270 3790 8310
rect 3690 8240 3790 8270
rect 3950 8410 4050 8440
rect 3950 8370 3980 8410
rect 4020 8370 4050 8410
rect 3950 8310 4050 8370
rect 3950 8270 3980 8310
rect 4020 8270 4050 8310
rect 3950 8240 4050 8270
rect 4080 8410 4180 8440
rect 4080 8370 4110 8410
rect 4150 8370 4180 8410
rect 4080 8310 4180 8370
rect 4080 8270 4110 8310
rect 4150 8270 4180 8310
rect 5440 8420 5470 8460
rect 5510 8420 5540 8460
rect 5440 8360 5540 8420
rect 5440 8320 5470 8360
rect 5510 8320 5540 8360
rect 5440 8290 5540 8320
rect 5660 8660 5760 8690
rect 5660 8620 5690 8660
rect 5730 8620 5760 8660
rect 5660 8560 5760 8620
rect 5660 8520 5690 8560
rect 5730 8520 5760 8560
rect 5660 8460 5760 8520
rect 5660 8420 5690 8460
rect 5730 8420 5760 8460
rect 5660 8360 5760 8420
rect 5660 8320 5690 8360
rect 5730 8320 5760 8360
rect 5660 8290 5760 8320
rect 5880 8660 5980 8690
rect 5880 8620 5910 8660
rect 5950 8620 5980 8660
rect 5880 8560 5980 8620
rect 5880 8520 5910 8560
rect 5950 8520 5980 8560
rect 5880 8460 5980 8520
rect 5880 8420 5910 8460
rect 5950 8420 5980 8460
rect 5880 8360 5980 8420
rect 5880 8320 5910 8360
rect 5950 8320 5980 8360
rect 5880 8290 5980 8320
rect 6100 8660 6200 8690
rect 6100 8620 6130 8660
rect 6170 8620 6200 8660
rect 6100 8560 6200 8620
rect 6100 8520 6130 8560
rect 6170 8520 6200 8560
rect 6100 8460 6200 8520
rect 6100 8420 6130 8460
rect 6170 8420 6200 8460
rect 6100 8360 6200 8420
rect 6100 8320 6130 8360
rect 6170 8320 6200 8360
rect 6100 8290 6200 8320
rect 6320 8660 6420 8690
rect 6520 8660 6620 8690
rect 6320 8620 6350 8660
rect 6390 8620 6420 8660
rect 6520 8620 6550 8660
rect 6590 8620 6620 8660
rect 6320 8560 6420 8620
rect 6520 8560 6620 8620
rect 6320 8520 6350 8560
rect 6390 8520 6420 8560
rect 6520 8520 6550 8560
rect 6590 8520 6620 8560
rect 6320 8460 6420 8520
rect 6520 8460 6620 8520
rect 6320 8420 6350 8460
rect 6390 8420 6420 8460
rect 6520 8420 6550 8460
rect 6590 8420 6620 8460
rect 6320 8360 6420 8420
rect 6520 8360 6620 8420
rect 6320 8320 6350 8360
rect 6390 8320 6420 8360
rect 6520 8320 6550 8360
rect 6590 8320 6620 8360
rect 6320 8290 6420 8320
rect 6520 8290 6620 8320
rect 6740 8660 6840 8690
rect 6740 8620 6770 8660
rect 6810 8620 6840 8660
rect 6740 8560 6840 8620
rect 6740 8520 6770 8560
rect 6810 8520 6840 8560
rect 6740 8460 6840 8520
rect 6740 8420 6770 8460
rect 6810 8420 6840 8460
rect 6740 8360 6840 8420
rect 6740 8320 6770 8360
rect 6810 8320 6840 8360
rect 6740 8290 6840 8320
rect 6960 8660 7060 8690
rect 6960 8620 6990 8660
rect 7030 8620 7060 8660
rect 6960 8560 7060 8620
rect 6960 8520 6990 8560
rect 7030 8520 7060 8560
rect 6960 8460 7060 8520
rect 6960 8420 6990 8460
rect 7030 8420 7060 8460
rect 6960 8360 7060 8420
rect 6960 8320 6990 8360
rect 7030 8320 7060 8360
rect 6960 8290 7060 8320
rect 7180 8660 7280 8690
rect 7180 8620 7210 8660
rect 7250 8620 7280 8660
rect 7180 8560 7280 8620
rect 7180 8520 7210 8560
rect 7250 8520 7280 8560
rect 7180 8460 7280 8520
rect 7180 8420 7210 8460
rect 7250 8420 7280 8460
rect 7180 8360 7280 8420
rect 7180 8320 7210 8360
rect 7250 8320 7280 8360
rect 7180 8290 7280 8320
rect 7400 8660 7500 8690
rect 7600 8660 7700 8690
rect 7400 8620 7430 8660
rect 7470 8620 7500 8660
rect 7600 8620 7630 8660
rect 7670 8620 7700 8660
rect 7400 8560 7500 8620
rect 7600 8560 7700 8620
rect 7400 8520 7430 8560
rect 7470 8520 7500 8560
rect 7600 8520 7630 8560
rect 7670 8520 7700 8560
rect 7400 8460 7500 8520
rect 7600 8460 7700 8520
rect 7400 8420 7430 8460
rect 7470 8420 7500 8460
rect 7600 8420 7630 8460
rect 7670 8420 7700 8460
rect 7400 8360 7500 8420
rect 7600 8360 7700 8420
rect 7400 8320 7430 8360
rect 7470 8320 7500 8360
rect 7600 8320 7630 8360
rect 7670 8320 7700 8360
rect 7400 8290 7500 8320
rect 7600 8290 7700 8320
rect 7820 8660 7920 8690
rect 7820 8620 7850 8660
rect 7890 8620 7920 8660
rect 7820 8560 7920 8620
rect 7820 8520 7850 8560
rect 7890 8520 7920 8560
rect 7820 8460 7920 8520
rect 7820 8420 7850 8460
rect 7890 8420 7920 8460
rect 7820 8360 7920 8420
rect 7820 8320 7850 8360
rect 7890 8320 7920 8360
rect 7820 8290 7920 8320
rect 8040 8660 8140 8690
rect 8040 8620 8070 8660
rect 8110 8620 8140 8660
rect 8040 8560 8140 8620
rect 8040 8520 8070 8560
rect 8110 8520 8140 8560
rect 8040 8460 8140 8520
rect 8040 8420 8070 8460
rect 8110 8420 8140 8460
rect 8040 8360 8140 8420
rect 8040 8320 8070 8360
rect 8110 8320 8140 8360
rect 8040 8290 8140 8320
rect 8260 8660 8360 8690
rect 8260 8620 8290 8660
rect 8330 8620 8360 8660
rect 8260 8560 8360 8620
rect 8260 8520 8290 8560
rect 8330 8520 8360 8560
rect 8260 8460 8360 8520
rect 8260 8420 8290 8460
rect 8330 8420 8360 8460
rect 8260 8360 8360 8420
rect 8260 8320 8290 8360
rect 8330 8320 8360 8360
rect 8260 8290 8360 8320
rect 8480 8660 8580 8690
rect 8480 8620 8510 8660
rect 8550 8620 8580 8660
rect 8480 8560 8580 8620
rect 8480 8520 8510 8560
rect 8550 8520 8580 8560
rect 8480 8460 8580 8520
rect 8480 8420 8510 8460
rect 8550 8420 8580 8460
rect 8480 8360 8580 8420
rect 8480 8320 8510 8360
rect 8550 8320 8580 8360
rect 8480 8290 8580 8320
rect 4080 8240 4180 8270
rect 5500 6030 5600 6060
rect 5500 5980 5530 6030
rect 5570 5980 5600 6030
rect 5500 5890 5600 5980
rect 5500 5840 5530 5890
rect 5570 5840 5600 5890
rect 5500 5810 5600 5840
rect 5700 6030 5800 6060
rect 5700 5980 5730 6030
rect 5770 5980 5800 6030
rect 5700 5890 5800 5980
rect 5700 5840 5730 5890
rect 5770 5840 5800 5890
rect 5700 5810 5800 5840
rect 5900 6030 6000 6060
rect 5900 5980 5930 6030
rect 5970 5980 6000 6030
rect 5900 5890 6000 5980
rect 5900 5840 5930 5890
rect 5970 5840 6000 5890
rect 5900 5810 6000 5840
rect 6100 6030 6200 6060
rect 6100 5980 6130 6030
rect 6170 5980 6200 6030
rect 6100 5890 6200 5980
rect 6100 5840 6130 5890
rect 6170 5840 6200 5890
rect 6100 5810 6200 5840
rect 6300 6030 6400 6060
rect 6300 5980 6330 6030
rect 6370 5980 6400 6030
rect 6300 5890 6400 5980
rect 6300 5840 6330 5890
rect 6370 5840 6400 5890
rect 6300 5810 6400 5840
rect 6500 6030 6600 6060
rect 6500 5980 6530 6030
rect 6570 5980 6600 6030
rect 6500 5890 6600 5980
rect 6500 5840 6530 5890
rect 6570 5840 6600 5890
rect 6500 5810 6600 5840
rect 6700 6030 6800 6060
rect 6700 5980 6730 6030
rect 6770 5980 6800 6030
rect 6700 5890 6800 5980
rect 6700 5840 6730 5890
rect 6770 5840 6800 5890
rect 6700 5810 6800 5840
rect 6900 6030 7000 6060
rect 6900 5980 6930 6030
rect 6970 5980 7000 6030
rect 6900 5890 7000 5980
rect 6900 5840 6930 5890
rect 6970 5840 7000 5890
rect 6900 5810 7000 5840
rect 7100 6030 7200 6060
rect 7100 5980 7130 6030
rect 7170 5980 7200 6030
rect 7100 5890 7200 5980
rect 7100 5840 7130 5890
rect 7170 5840 7200 5890
rect 7100 5810 7200 5840
rect 7300 6030 7400 6060
rect 7300 5980 7330 6030
rect 7370 5980 7400 6030
rect 7300 5890 7400 5980
rect 7300 5840 7330 5890
rect 7370 5840 7400 5890
rect 7300 5810 7400 5840
rect 7500 6030 7600 6060
rect 7500 5980 7530 6030
rect 7570 5980 7600 6030
rect 7500 5890 7600 5980
rect 7500 5840 7530 5890
rect 7570 5840 7600 5890
rect 7500 5810 7600 5840
rect 5550 5340 5650 5370
rect 5550 5300 5580 5340
rect 5620 5300 5650 5340
rect 5550 5270 5650 5300
rect 5680 5340 5780 5370
rect 5680 5300 5710 5340
rect 5750 5300 5780 5340
rect 5680 5270 5780 5300
rect 5810 5340 5910 5370
rect 5810 5300 5840 5340
rect 5880 5300 5910 5340
rect 5810 5270 5910 5300
rect 5940 5340 6040 5370
rect 5940 5300 5970 5340
rect 6010 5300 6040 5340
rect 5940 5270 6040 5300
rect 6070 5340 6170 5370
rect 6070 5300 6100 5340
rect 6140 5300 6170 5340
rect 6070 5270 6170 5300
rect 6200 5340 6300 5370
rect 6200 5300 6230 5340
rect 6270 5300 6300 5340
rect 6200 5270 6300 5300
rect 6330 5340 6430 5370
rect 6330 5300 6360 5340
rect 6400 5300 6430 5340
rect 6330 5270 6430 5300
rect 6690 5340 6790 5370
rect 6690 5300 6720 5340
rect 6760 5300 6790 5340
rect 6690 5270 6790 5300
rect 6820 5340 6920 5370
rect 6820 5300 6850 5340
rect 6890 5300 6920 5340
rect 6820 5270 6920 5300
rect 6950 5340 7050 5370
rect 6950 5300 6980 5340
rect 7020 5300 7050 5340
rect 6950 5270 7050 5300
rect 7080 5340 7180 5370
rect 7080 5300 7110 5340
rect 7150 5300 7180 5340
rect 7080 5270 7180 5300
rect 7210 5340 7310 5370
rect 7210 5300 7240 5340
rect 7280 5300 7310 5340
rect 7210 5270 7310 5300
rect 7340 5340 7440 5370
rect 7340 5300 7370 5340
rect 7410 5300 7440 5340
rect 7340 5270 7440 5300
rect 7470 5340 7570 5370
rect 7470 5300 7500 5340
rect 7540 5300 7570 5340
rect 7470 5270 7570 5300
rect 7830 5340 7930 5370
rect 7830 5300 7860 5340
rect 7900 5300 7930 5340
rect 7830 5270 7930 5300
rect 7960 5340 8060 5370
rect 7960 5300 7990 5340
rect 8030 5300 8060 5340
rect 7960 5270 8060 5300
rect 8090 5340 8190 5370
rect 8090 5300 8120 5340
rect 8160 5300 8190 5340
rect 8090 5270 8190 5300
rect 8220 5340 8320 5370
rect 8220 5300 8250 5340
rect 8290 5300 8320 5340
rect 8220 5270 8320 5300
rect 8350 5340 8450 5370
rect 8350 5300 8380 5340
rect 8420 5300 8450 5340
rect 8350 5270 8450 5300
rect 8480 5340 8580 5370
rect 8480 5300 8510 5340
rect 8550 5300 8580 5340
rect 8480 5270 8580 5300
rect 8610 5340 8710 5370
rect 8610 5300 8640 5340
rect 8680 5300 8710 5340
rect 8610 5270 8710 5300
rect -1630 3740 -1550 3770
rect -1630 3700 -1610 3740
rect -1570 3700 -1550 3740
rect -1630 3670 -1550 3700
rect -1510 3740 -1430 3770
rect -1510 3700 -1490 3740
rect -1450 3700 -1430 3740
rect -1510 3670 -1430 3700
rect -1390 3740 -1310 3770
rect -1390 3700 -1370 3740
rect -1330 3700 -1310 3740
rect -1390 3670 -1310 3700
rect -1270 3740 -1190 3770
rect -1270 3700 -1250 3740
rect -1210 3700 -1190 3740
rect -1270 3670 -1190 3700
rect -1150 3740 -1070 3770
rect -1150 3700 -1130 3740
rect -1090 3700 -1070 3740
rect -1150 3670 -1070 3700
rect -1030 3740 -950 3770
rect -1030 3700 -1010 3740
rect -970 3700 -950 3740
rect -1030 3670 -950 3700
rect -910 3740 -830 3770
rect -910 3700 -890 3740
rect -850 3700 -830 3740
rect -910 3670 -830 3700
rect -790 3740 -710 3770
rect -790 3700 -770 3740
rect -730 3700 -710 3740
rect -790 3670 -710 3700
rect -670 3740 -590 3770
rect -670 3700 -650 3740
rect -610 3700 -590 3740
rect -670 3670 -590 3700
rect -550 3740 -470 3770
rect -550 3700 -530 3740
rect -490 3700 -470 3740
rect -550 3670 -470 3700
rect -430 3740 -350 3770
rect -430 3700 -410 3740
rect -370 3700 -350 3740
rect -430 3670 -350 3700
rect 930 3740 1010 3770
rect 930 3700 950 3740
rect 990 3700 1010 3740
rect 930 3670 1010 3700
rect 1050 3740 1130 3770
rect 1050 3700 1070 3740
rect 1110 3700 1130 3740
rect 1050 3670 1130 3700
rect 1170 3740 1250 3770
rect 1170 3700 1190 3740
rect 1230 3700 1250 3740
rect 1170 3670 1250 3700
rect 1290 3740 1370 3770
rect 1290 3700 1310 3740
rect 1350 3700 1370 3740
rect 1290 3670 1370 3700
rect 1410 3740 1490 3770
rect 1410 3700 1430 3740
rect 1470 3700 1490 3740
rect 1410 3670 1490 3700
rect 1530 3740 1610 3770
rect 1530 3700 1550 3740
rect 1590 3700 1610 3740
rect 1530 3670 1610 3700
rect 1650 3740 1730 3770
rect 1650 3700 1670 3740
rect 1710 3700 1730 3740
rect 1650 3670 1730 3700
rect 1770 3740 1850 3770
rect 1770 3700 1790 3740
rect 1830 3700 1850 3740
rect 1770 3670 1850 3700
rect 1890 3740 1970 3770
rect 1890 3700 1910 3740
rect 1950 3700 1970 3740
rect 1890 3670 1970 3700
rect 2010 3740 2090 3770
rect 2010 3700 2030 3740
rect 2070 3700 2090 3740
rect 2010 3670 2090 3700
rect 2130 3740 2210 3770
rect 2130 3700 2150 3740
rect 2190 3700 2210 3740
rect 2130 3670 2210 3700
rect -2250 3130 -2170 3160
rect -2250 3090 -2230 3130
rect -2190 3090 -2170 3130
rect -2250 3030 -2170 3090
rect -2250 2990 -2230 3030
rect -2190 2990 -2170 3030
rect -2250 2930 -2170 2990
rect -2250 2890 -2230 2930
rect -2190 2890 -2170 2930
rect -2250 2830 -2170 2890
rect -2250 2790 -2230 2830
rect -2190 2790 -2170 2830
rect -2250 2730 -2170 2790
rect -2250 2690 -2230 2730
rect -2190 2690 -2170 2730
rect -2250 2660 -2170 2690
rect -1170 3130 -1090 3160
rect -1010 3130 -930 3160
rect -1170 3090 -1150 3130
rect -1110 3090 -1090 3130
rect -1010 3090 -990 3130
rect -950 3090 -930 3130
rect -1170 3030 -1090 3090
rect -1010 3030 -930 3090
rect -1170 2990 -1150 3030
rect -1110 2990 -1090 3030
rect -1010 2990 -990 3030
rect -950 2990 -930 3030
rect -1170 2930 -1090 2990
rect -1010 2930 -930 2990
rect -1170 2890 -1150 2930
rect -1110 2890 -1090 2930
rect -1010 2890 -990 2930
rect -950 2890 -930 2930
rect -1170 2830 -1090 2890
rect -1010 2830 -930 2890
rect -1170 2790 -1150 2830
rect -1110 2790 -1090 2830
rect -1010 2790 -990 2830
rect -950 2790 -930 2830
rect -1170 2730 -1090 2790
rect -1010 2730 -930 2790
rect -1170 2690 -1150 2730
rect -1110 2690 -1090 2730
rect -1010 2690 -990 2730
rect -950 2690 -930 2730
rect -1170 2660 -1090 2690
rect -1010 2660 -930 2690
rect 70 3130 150 3160
rect 70 3090 90 3130
rect 130 3090 150 3130
rect 70 3030 150 3090
rect 70 2990 90 3030
rect 130 2990 150 3030
rect 70 2930 150 2990
rect 70 2890 90 2930
rect 130 2890 150 2930
rect 70 2830 150 2890
rect 70 2790 90 2830
rect 130 2790 150 2830
rect 70 2730 150 2790
rect 70 2690 90 2730
rect 130 2690 150 2730
rect 70 2660 150 2690
rect 430 3130 510 3160
rect 430 3090 450 3130
rect 490 3090 510 3130
rect 430 3030 510 3090
rect 430 2990 450 3030
rect 490 2990 510 3030
rect 430 2930 510 2990
rect 430 2890 450 2930
rect 490 2890 510 2930
rect 430 2830 510 2890
rect 430 2790 450 2830
rect 490 2790 510 2830
rect 430 2730 510 2790
rect 430 2690 450 2730
rect 490 2690 510 2730
rect 430 2660 510 2690
rect 1510 3130 1590 3160
rect 1670 3130 1750 3160
rect 1510 3090 1530 3130
rect 1570 3090 1590 3130
rect 1670 3090 1690 3130
rect 1730 3090 1750 3130
rect 1510 3030 1590 3090
rect 1670 3030 1750 3090
rect 1510 2990 1530 3030
rect 1570 2990 1590 3030
rect 1670 2990 1690 3030
rect 1730 2990 1750 3030
rect 1510 2930 1590 2990
rect 1670 2930 1750 2990
rect 1510 2890 1530 2930
rect 1570 2890 1590 2930
rect 1670 2890 1690 2930
rect 1730 2890 1750 2930
rect 1510 2830 1590 2890
rect 1670 2830 1750 2890
rect 1510 2790 1530 2830
rect 1570 2790 1590 2830
rect 1670 2790 1690 2830
rect 1730 2790 1750 2830
rect 1510 2730 1590 2790
rect 1670 2730 1750 2790
rect 1510 2690 1530 2730
rect 1570 2690 1590 2730
rect 1670 2690 1690 2730
rect 1730 2690 1750 2730
rect 1510 2670 1590 2690
rect 1670 2670 1750 2690
rect 1510 2660 1750 2670
rect 2750 3130 2830 3160
rect 2750 3090 2770 3130
rect 2810 3090 2830 3130
rect 2750 3030 2830 3090
rect 2750 2990 2770 3030
rect 2810 2990 2830 3030
rect 2750 2930 2830 2990
rect 2750 2890 2770 2930
rect 2810 2890 2830 2930
rect 2750 2830 2830 2890
rect 2750 2790 2770 2830
rect 2810 2790 2830 2830
rect 2750 2730 2830 2790
rect 2750 2690 2770 2730
rect 2810 2690 2830 2730
rect 2750 2660 2830 2690
rect -1830 2220 -1750 2250
rect -1830 2180 -1810 2220
rect -1770 2180 -1750 2220
rect -1830 2120 -1750 2180
rect -1830 2080 -1810 2120
rect -1770 2080 -1750 2120
rect -1830 2050 -1750 2080
rect 250 2220 330 2250
rect 250 2180 270 2220
rect 310 2180 330 2220
rect 250 2120 330 2180
rect 250 2080 270 2120
rect 310 2080 330 2120
rect 250 2050 330 2080
rect 2330 2220 2410 2250
rect 2330 2180 2350 2220
rect 2390 2180 2410 2220
rect 2330 2120 2410 2180
rect 2330 2080 2350 2120
rect 2390 2080 2410 2120
rect 2330 2050 2410 2080
<< pdiff >>
rect -1300 12490 -1220 12520
rect -1300 12450 -1280 12490
rect -1240 12450 -1220 12490
rect -1300 12420 -1220 12450
rect -1190 12490 -1110 12520
rect -1190 12450 -1170 12490
rect -1130 12450 -1110 12490
rect -1190 12420 -1110 12450
rect -880 12490 -800 12520
rect -880 12450 -860 12490
rect -820 12450 -800 12490
rect -880 12420 -800 12450
rect -770 12490 -690 12520
rect -770 12450 -750 12490
rect -710 12450 -690 12490
rect -770 12420 -690 12450
rect -660 12490 -580 12520
rect -660 12450 -640 12490
rect -600 12450 -580 12490
rect -660 12420 -580 12450
rect -210 12490 -130 12520
rect -210 12450 -190 12490
rect -150 12450 -130 12490
rect -210 12420 -130 12450
rect -100 12490 -20 12520
rect -100 12450 -80 12490
rect -40 12450 -20 12490
rect -100 12420 -20 12450
rect 10 12490 90 12520
rect 10 12450 30 12490
rect 70 12450 90 12490
rect 10 12420 90 12450
rect 230 12490 310 12520
rect 230 12450 250 12490
rect 290 12450 310 12490
rect 230 12420 310 12450
rect 340 12490 420 12520
rect 340 12450 360 12490
rect 400 12450 420 12490
rect 340 12420 420 12450
rect 450 12490 530 12520
rect 450 12450 470 12490
rect 510 12450 530 12490
rect 450 12420 530 12450
rect 560 12490 640 12520
rect 560 12450 580 12490
rect 620 12450 640 12490
rect 560 12420 640 12450
rect 1070 12490 1150 12520
rect 1070 12450 1090 12490
rect 1130 12450 1150 12490
rect 1070 12420 1150 12450
rect 1180 12490 1260 12520
rect 1180 12450 1200 12490
rect 1240 12450 1260 12490
rect 1180 12420 1260 12450
rect 1490 12490 1570 12520
rect 1490 12450 1510 12490
rect 1550 12450 1570 12490
rect 1490 12420 1570 12450
rect 1600 12490 1680 12520
rect 1600 12450 1620 12490
rect 1660 12450 1680 12490
rect 1600 12420 1680 12450
rect 1710 12490 1790 12520
rect 1710 12450 1730 12490
rect 1770 12450 1790 12490
rect 1710 12420 1790 12450
rect 1940 12490 2020 12520
rect 1940 12450 1960 12490
rect 2000 12450 2020 12490
rect 1940 12420 2020 12450
rect 2050 12490 2130 12520
rect 2050 12450 2070 12490
rect 2110 12450 2130 12490
rect 2050 12420 2130 12450
rect 2160 12490 2240 12520
rect 2160 12450 2180 12490
rect 2220 12450 2240 12490
rect 2160 12420 2240 12450
rect 2300 12490 2380 12520
rect 2300 12450 2320 12490
rect 2360 12450 2380 12490
rect 2300 12420 2380 12450
rect 2410 12490 2490 12520
rect 2410 12450 2430 12490
rect 2470 12450 2490 12490
rect 2410 12420 2490 12450
rect 2520 12490 2600 12520
rect 2520 12450 2540 12490
rect 2580 12450 2600 12490
rect 2520 12420 2600 12450
rect 2880 12490 2960 12520
rect 2880 12450 2900 12490
rect 2940 12450 2960 12490
rect 2880 12420 2960 12450
rect 2990 12490 3070 12520
rect 2990 12450 3010 12490
rect 3050 12450 3070 12490
rect 2990 12420 3070 12450
rect 3100 12490 3180 12520
rect 3100 12450 3120 12490
rect 3160 12450 3180 12490
rect 3100 12420 3180 12450
rect 3320 12490 3400 12520
rect 3320 12450 3340 12490
rect 3380 12450 3400 12490
rect 3320 12420 3400 12450
rect 3430 12490 3510 12520
rect 3430 12450 3450 12490
rect 3490 12450 3510 12490
rect 3430 12420 3510 12450
rect 3540 12490 3620 12520
rect 3540 12450 3560 12490
rect 3600 12450 3620 12490
rect 3540 12420 3620 12450
rect 3940 12490 4020 12520
rect 3940 12450 3960 12490
rect 4000 12450 4020 12490
rect 3940 12420 4020 12450
rect 4050 12490 4130 12520
rect 4050 12450 4070 12490
rect 4110 12450 4130 12490
rect 4050 12420 4130 12450
rect 4280 12490 4360 12520
rect 4280 12450 4300 12490
rect 4340 12450 4360 12490
rect 4280 12420 4360 12450
rect 4390 12490 4470 12520
rect 4390 12450 4410 12490
rect 4450 12450 4470 12490
rect 4390 12420 4470 12450
rect 4500 12490 4580 12520
rect 4500 12450 4520 12490
rect 4560 12450 4580 12490
rect 4500 12420 4580 12450
rect 4640 12490 4720 12520
rect 4640 12450 4660 12490
rect 4700 12450 4720 12490
rect 4640 12420 4720 12450
rect 4750 12490 4830 12520
rect 4750 12450 4770 12490
rect 4810 12450 4830 12490
rect 4750 12420 4830 12450
rect 4860 12490 4940 12520
rect 4860 12450 4880 12490
rect 4920 12450 4940 12490
rect 4860 12420 4940 12450
rect 5240 12490 5320 12520
rect 5240 12450 5260 12490
rect 5300 12450 5320 12490
rect 5240 12420 5320 12450
rect 5350 12490 5430 12520
rect 5350 12450 5370 12490
rect 5410 12450 5430 12490
rect 5350 12420 5430 12450
rect 5580 12490 5660 12520
rect 5580 12450 5600 12490
rect 5640 12450 5660 12490
rect 5580 12420 5660 12450
rect 5690 12490 5770 12520
rect 5690 12450 5710 12490
rect 5750 12450 5770 12490
rect 5690 12420 5770 12450
rect 5800 12490 5880 12520
rect 5800 12450 5820 12490
rect 5860 12450 5880 12490
rect 5800 12420 5880 12450
rect 5940 12490 6020 12520
rect 5940 12450 5960 12490
rect 6000 12450 6020 12490
rect 5940 12420 6020 12450
rect 6050 12490 6130 12520
rect 6050 12450 6070 12490
rect 6110 12450 6130 12490
rect 6050 12420 6130 12450
rect 6160 12490 6240 12520
rect 6160 12450 6180 12490
rect 6220 12450 6240 12490
rect 6160 12420 6240 12450
rect 6540 12490 6620 12520
rect 6540 12450 6560 12490
rect 6600 12450 6620 12490
rect 6540 12420 6620 12450
rect 6650 12490 6730 12520
rect 6650 12450 6670 12490
rect 6710 12450 6730 12490
rect 6650 12420 6730 12450
rect 6880 12490 6960 12520
rect 6880 12450 6900 12490
rect 6940 12450 6960 12490
rect 6880 12420 6960 12450
rect 6990 12490 7070 12520
rect 6990 12450 7010 12490
rect 7050 12450 7070 12490
rect 6990 12420 7070 12450
rect 7100 12490 7180 12520
rect 7100 12450 7120 12490
rect 7160 12450 7180 12490
rect 7100 12420 7180 12450
rect 7240 12490 7320 12520
rect 7240 12450 7260 12490
rect 7300 12450 7320 12490
rect 7240 12420 7320 12450
rect 7350 12490 7430 12520
rect 7350 12450 7370 12490
rect 7410 12450 7430 12490
rect 7350 12420 7430 12450
rect 7460 12490 7540 12520
rect 7460 12450 7480 12490
rect 7520 12450 7540 12490
rect 7460 12420 7540 12450
rect 7840 12490 7920 12520
rect 7840 12450 7860 12490
rect 7900 12450 7920 12490
rect 7840 12420 7920 12450
rect 7950 12490 8030 12520
rect 7950 12450 7970 12490
rect 8010 12450 8030 12490
rect 7950 12420 8030 12450
rect 8180 12490 8260 12520
rect 8180 12450 8200 12490
rect 8240 12450 8260 12490
rect 8180 12420 8260 12450
rect 8290 12490 8370 12520
rect 8290 12450 8310 12490
rect 8350 12450 8370 12490
rect 8290 12420 8370 12450
rect 8400 12490 8480 12520
rect 8400 12450 8420 12490
rect 8460 12450 8480 12490
rect 8400 12420 8480 12450
rect 8540 12490 8620 12520
rect 8540 12450 8560 12490
rect 8600 12450 8620 12490
rect 8540 12420 8620 12450
rect 8650 12490 8730 12520
rect 8650 12450 8670 12490
rect 8710 12450 8730 12490
rect 8650 12420 8730 12450
rect 8760 12490 8840 12520
rect 8760 12450 8780 12490
rect 8820 12450 8840 12490
rect 8760 12420 8840 12450
rect 9300 12340 9380 12370
rect 9300 12300 9320 12340
rect 9360 12300 9380 12340
rect 9300 12240 9380 12300
rect 9300 12200 9320 12240
rect 9360 12200 9380 12240
rect 9300 12170 9380 12200
rect 9410 12340 9490 12370
rect 9410 12300 9430 12340
rect 9470 12300 9490 12340
rect 9410 12240 9490 12300
rect 9410 12200 9430 12240
rect 9470 12200 9490 12240
rect 9410 12170 9490 12200
rect 9820 12340 9900 12370
rect 9820 12300 9840 12340
rect 9880 12300 9900 12340
rect 9820 12240 9900 12300
rect 9820 12200 9840 12240
rect 9880 12200 9900 12240
rect 9820 12170 9900 12200
rect 9930 12340 10010 12370
rect 9930 12300 9950 12340
rect 9990 12300 10010 12340
rect 9930 12240 10010 12300
rect 9930 12200 9950 12240
rect 9990 12200 10010 12240
rect 9930 12170 10010 12200
rect 10340 12340 10420 12370
rect 10340 12300 10360 12340
rect 10400 12300 10420 12340
rect 10340 12240 10420 12300
rect 10340 12200 10360 12240
rect 10400 12200 10420 12240
rect 10340 12170 10420 12200
rect 10450 12340 10530 12370
rect 10450 12300 10470 12340
rect 10510 12300 10530 12340
rect 10450 12240 10530 12300
rect 10450 12200 10470 12240
rect 10510 12200 10530 12240
rect 10450 12170 10530 12200
rect 9300 11960 9380 11990
rect 9300 11920 9320 11960
rect 9360 11920 9380 11960
rect 9300 11860 9380 11920
rect 9300 11820 9320 11860
rect 9360 11820 9380 11860
rect 9300 11760 9380 11820
rect 9300 11720 9320 11760
rect 9360 11720 9380 11760
rect 9300 11660 9380 11720
rect 9300 11620 9320 11660
rect 9360 11620 9380 11660
rect 9300 11590 9380 11620
rect 9410 11960 9490 11990
rect 9410 11920 9430 11960
rect 9470 11920 9490 11960
rect 9410 11860 9490 11920
rect 9410 11820 9430 11860
rect 9470 11820 9490 11860
rect 9410 11760 9490 11820
rect 9410 11720 9430 11760
rect 9470 11720 9490 11760
rect 9410 11660 9490 11720
rect 9410 11620 9430 11660
rect 9470 11620 9490 11660
rect 9410 11590 9490 11620
rect 9820 11960 9900 11990
rect 9820 11920 9840 11960
rect 9880 11920 9900 11960
rect 9820 11860 9900 11920
rect 9820 11820 9840 11860
rect 9880 11820 9900 11860
rect 9820 11760 9900 11820
rect 9820 11720 9840 11760
rect 9880 11720 9900 11760
rect 9820 11660 9900 11720
rect 9820 11620 9840 11660
rect 9880 11620 9900 11660
rect 9820 11590 9900 11620
rect 9930 11960 10010 11990
rect 9930 11920 9950 11960
rect 9990 11920 10010 11960
rect 9930 11860 10010 11920
rect 9930 11820 9950 11860
rect 9990 11820 10010 11860
rect 9930 11760 10010 11820
rect 9930 11720 9950 11760
rect 9990 11720 10010 11760
rect 9930 11660 10010 11720
rect 9930 11620 9950 11660
rect 9990 11620 10010 11660
rect 9930 11590 10010 11620
rect 10340 11960 10420 11990
rect 10340 11920 10360 11960
rect 10400 11920 10420 11960
rect 10340 11860 10420 11920
rect 10340 11820 10360 11860
rect 10400 11820 10420 11860
rect 10340 11760 10420 11820
rect 10340 11720 10360 11760
rect 10400 11720 10420 11760
rect 10340 11660 10420 11720
rect 10340 11620 10360 11660
rect 10400 11620 10420 11660
rect 10340 11590 10420 11620
rect 10450 11960 10530 11990
rect 10450 11920 10470 11960
rect 10510 11920 10530 11960
rect 10450 11860 10530 11920
rect 10450 11820 10470 11860
rect 10510 11820 10530 11860
rect 10450 11760 10530 11820
rect 10450 11720 10470 11760
rect 10510 11720 10530 11760
rect 10450 11660 10530 11720
rect 10450 11620 10470 11660
rect 10510 11620 10530 11660
rect 10450 11590 10530 11620
rect 9300 11270 9380 11300
rect 9300 11230 9320 11270
rect 9360 11230 9380 11270
rect 9300 11170 9380 11230
rect 9300 11130 9320 11170
rect 9360 11130 9380 11170
rect 9300 11070 9380 11130
rect 9300 11030 9320 11070
rect 9360 11030 9380 11070
rect 9300 10970 9380 11030
rect 9300 10930 9320 10970
rect 9360 10930 9380 10970
rect 9300 10900 9380 10930
rect 9680 11270 9760 11300
rect 9680 11230 9700 11270
rect 9740 11230 9760 11270
rect 9680 11170 9760 11230
rect 9680 11130 9700 11170
rect 9740 11130 9760 11170
rect 9680 11070 9760 11130
rect 9680 11030 9700 11070
rect 9740 11030 9760 11070
rect 9680 10970 9760 11030
rect 9680 10930 9700 10970
rect 9740 10930 9760 10970
rect 9680 10900 9760 10930
rect 9820 11270 9900 11300
rect 9820 11230 9840 11270
rect 9880 11230 9900 11270
rect 9820 11170 9900 11230
rect 9820 11130 9840 11170
rect 9880 11130 9900 11170
rect 9820 11070 9900 11130
rect 9820 11030 9840 11070
rect 9880 11030 9900 11070
rect 9820 10970 9900 11030
rect 9820 10930 9840 10970
rect 9880 10930 9900 10970
rect 9820 10900 9900 10930
rect 10200 11270 10280 11300
rect 10200 11230 10220 11270
rect 10260 11230 10280 11270
rect 10200 11170 10280 11230
rect 10200 11130 10220 11170
rect 10260 11130 10280 11170
rect 10200 11070 10280 11130
rect 10200 11030 10220 11070
rect 10260 11030 10280 11070
rect 10200 10970 10280 11030
rect 10200 10930 10220 10970
rect 10260 10930 10280 10970
rect 10200 10900 10280 10930
rect 10340 11270 10420 11300
rect 10340 11230 10360 11270
rect 10400 11230 10420 11270
rect 10340 11170 10420 11230
rect 10340 11130 10360 11170
rect 10400 11130 10420 11170
rect 10340 11070 10420 11130
rect 10340 11030 10360 11070
rect 10400 11030 10420 11070
rect 10340 10970 10420 11030
rect 10340 10930 10360 10970
rect 10400 10930 10420 10970
rect 10340 10900 10420 10930
rect 10720 11270 10800 11300
rect 10720 11230 10740 11270
rect 10780 11230 10800 11270
rect 10720 11170 10800 11230
rect 10720 11130 10740 11170
rect 10780 11130 10800 11170
rect 10720 11070 10800 11130
rect 10720 11030 10740 11070
rect 10780 11030 10800 11070
rect 10720 10970 10800 11030
rect 10720 10930 10740 10970
rect 10780 10930 10800 10970
rect 10720 10900 10800 10930
rect 10860 11270 10940 11300
rect 10860 11230 10880 11270
rect 10920 11230 10940 11270
rect 10860 11170 10940 11230
rect 10860 11130 10880 11170
rect 10920 11130 10940 11170
rect 10860 11070 10940 11130
rect 10860 11030 10880 11070
rect 10920 11030 10940 11070
rect 10860 10970 10940 11030
rect 10860 10930 10880 10970
rect 10920 10930 10940 10970
rect 10860 10900 10940 10930
rect 11240 11270 11320 11300
rect 11240 11230 11260 11270
rect 11300 11230 11320 11270
rect 11240 11170 11320 11230
rect 11240 11130 11260 11170
rect 11300 11130 11320 11170
rect 11240 11070 11320 11130
rect 11240 11030 11260 11070
rect 11300 11030 11320 11070
rect 11240 10970 11320 11030
rect 11240 10930 11260 10970
rect 11300 10930 11320 10970
rect 11240 10900 11320 10930
rect -640 9790 -560 9820
rect -640 9750 -620 9790
rect -580 9750 -560 9790
rect -640 9690 -560 9750
rect -640 9650 -620 9690
rect -580 9650 -560 9690
rect -640 9590 -560 9650
rect -640 9550 -620 9590
rect -580 9550 -560 9590
rect -640 9490 -560 9550
rect -640 9450 -620 9490
rect -580 9450 -560 9490
rect -640 9420 -560 9450
rect -530 9790 -450 9820
rect -530 9750 -510 9790
rect -470 9750 -450 9790
rect -530 9690 -450 9750
rect -530 9650 -510 9690
rect -470 9650 -450 9690
rect -530 9590 -450 9650
rect -530 9550 -510 9590
rect -470 9550 -450 9590
rect -530 9490 -450 9550
rect -530 9450 -510 9490
rect -470 9450 -450 9490
rect -530 9420 -450 9450
rect -420 9790 -340 9820
rect -420 9750 -400 9790
rect -360 9750 -340 9790
rect -420 9690 -340 9750
rect -420 9650 -400 9690
rect -360 9650 -340 9690
rect -420 9590 -340 9650
rect -420 9550 -400 9590
rect -360 9550 -340 9590
rect -420 9490 -340 9550
rect -420 9450 -400 9490
rect -360 9450 -340 9490
rect -420 9420 -340 9450
rect -120 9790 -40 9820
rect -120 9750 -100 9790
rect -60 9750 -40 9790
rect -120 9690 -40 9750
rect -120 9650 -100 9690
rect -60 9650 -40 9690
rect -120 9590 -40 9650
rect -120 9550 -100 9590
rect -60 9550 -40 9590
rect -120 9490 -40 9550
rect -120 9450 -100 9490
rect -60 9450 -40 9490
rect -120 9420 -40 9450
rect -10 9790 70 9820
rect -10 9750 10 9790
rect 50 9750 70 9790
rect -10 9690 70 9750
rect -10 9650 10 9690
rect 50 9650 70 9690
rect -10 9590 70 9650
rect -10 9550 10 9590
rect 50 9550 70 9590
rect -10 9490 70 9550
rect -10 9450 10 9490
rect 50 9450 70 9490
rect -10 9420 70 9450
rect 100 9790 180 9820
rect 260 9790 340 9820
rect 100 9750 120 9790
rect 160 9750 180 9790
rect 260 9750 280 9790
rect 320 9750 340 9790
rect 100 9690 180 9750
rect 260 9690 340 9750
rect 100 9650 120 9690
rect 160 9650 180 9690
rect 260 9650 280 9690
rect 320 9650 340 9690
rect 100 9590 180 9650
rect 260 9590 340 9650
rect 100 9550 120 9590
rect 160 9550 180 9590
rect 260 9550 280 9590
rect 320 9550 340 9590
rect 100 9490 180 9550
rect 260 9490 340 9550
rect 100 9450 120 9490
rect 160 9450 180 9490
rect 260 9450 280 9490
rect 320 9450 340 9490
rect 100 9420 180 9450
rect 260 9420 340 9450
rect 370 9790 450 9820
rect 370 9750 390 9790
rect 430 9750 450 9790
rect 370 9690 450 9750
rect 370 9650 390 9690
rect 430 9650 450 9690
rect 370 9590 450 9650
rect 370 9550 390 9590
rect 430 9550 450 9590
rect 370 9490 450 9550
rect 370 9450 390 9490
rect 430 9450 450 9490
rect 370 9420 450 9450
rect 480 9790 560 9820
rect 480 9750 500 9790
rect 540 9750 560 9790
rect 480 9690 560 9750
rect 480 9650 500 9690
rect 540 9650 560 9690
rect 480 9590 560 9650
rect 480 9550 500 9590
rect 540 9550 560 9590
rect 480 9490 560 9550
rect 480 9450 500 9490
rect 540 9450 560 9490
rect 480 9420 560 9450
rect 780 9790 860 9820
rect 780 9750 800 9790
rect 840 9750 860 9790
rect 780 9690 860 9750
rect 780 9650 800 9690
rect 840 9650 860 9690
rect 780 9590 860 9650
rect 780 9550 800 9590
rect 840 9550 860 9590
rect 780 9490 860 9550
rect 780 9450 800 9490
rect 840 9450 860 9490
rect 780 9420 860 9450
rect 890 9790 970 9820
rect 890 9750 910 9790
rect 950 9750 970 9790
rect 890 9690 970 9750
rect 890 9650 910 9690
rect 950 9650 970 9690
rect 890 9590 970 9650
rect 890 9550 910 9590
rect 950 9550 970 9590
rect 890 9490 970 9550
rect 890 9450 910 9490
rect 950 9450 970 9490
rect 890 9420 970 9450
rect 1000 9790 1080 9820
rect 1000 9750 1020 9790
rect 1060 9750 1080 9790
rect 1000 9690 1080 9750
rect 1000 9650 1020 9690
rect 1060 9650 1080 9690
rect 1000 9590 1080 9650
rect 1000 9550 1020 9590
rect 1060 9550 1080 9590
rect 1000 9490 1080 9550
rect 1000 9450 1020 9490
rect 1060 9450 1080 9490
rect 1000 9420 1080 9450
rect 1300 9790 1380 9820
rect 1300 9750 1320 9790
rect 1360 9750 1380 9790
rect 1300 9690 1380 9750
rect 1300 9650 1320 9690
rect 1360 9650 1380 9690
rect 1300 9590 1380 9650
rect 1300 9550 1320 9590
rect 1360 9550 1380 9590
rect 1300 9490 1380 9550
rect 1300 9450 1320 9490
rect 1360 9450 1380 9490
rect 1300 9430 1380 9450
rect 1280 9420 1380 9430
rect 1410 9790 1490 9820
rect 1410 9750 1430 9790
rect 1470 9750 1490 9790
rect 1410 9690 1490 9750
rect 1410 9650 1430 9690
rect 1470 9650 1490 9690
rect 1410 9590 1490 9650
rect 1410 9550 1430 9590
rect 1470 9550 1490 9590
rect 1410 9490 1490 9550
rect 1410 9450 1430 9490
rect 1470 9450 1490 9490
rect 1410 9420 1490 9450
rect 1520 9790 1600 9820
rect 1520 9750 1540 9790
rect 1580 9750 1600 9790
rect 1520 9690 1600 9750
rect 1520 9650 1540 9690
rect 1580 9650 1600 9690
rect 1520 9590 1600 9650
rect 1520 9550 1540 9590
rect 1580 9550 1600 9590
rect 1520 9490 1600 9550
rect 1520 9450 1540 9490
rect 1580 9450 1600 9490
rect 1520 9420 1600 9450
rect 1740 9790 1820 9820
rect 1740 9750 1760 9790
rect 1800 9750 1820 9790
rect 1740 9690 1820 9750
rect 1740 9650 1760 9690
rect 1800 9650 1820 9690
rect 1740 9590 1820 9650
rect 1740 9550 1760 9590
rect 1800 9550 1820 9590
rect 1740 9490 1820 9550
rect 1740 9450 1760 9490
rect 1800 9450 1820 9490
rect 1740 9420 1820 9450
rect 1850 9790 1930 9820
rect 1850 9750 1870 9790
rect 1910 9750 1930 9790
rect 1850 9690 1930 9750
rect 1850 9650 1870 9690
rect 1910 9650 1930 9690
rect 1850 9590 1930 9650
rect 1850 9550 1870 9590
rect 1910 9550 1930 9590
rect 1850 9490 1930 9550
rect 1850 9450 1870 9490
rect 1910 9450 1930 9490
rect 1850 9420 1930 9450
rect 2070 9790 2150 9820
rect 2070 9750 2090 9790
rect 2130 9750 2150 9790
rect 2070 9690 2150 9750
rect 2070 9650 2090 9690
rect 2130 9650 2150 9690
rect 2070 9590 2150 9650
rect 2070 9550 2090 9590
rect 2130 9550 2150 9590
rect 2070 9490 2150 9550
rect 2070 9450 2090 9490
rect 2130 9450 2150 9490
rect 2070 9420 2150 9450
rect 2180 9790 2260 9820
rect 2180 9750 2200 9790
rect 2240 9750 2260 9790
rect 2180 9690 2260 9750
rect 2180 9650 2200 9690
rect 2240 9650 2260 9690
rect 2180 9590 2260 9650
rect 2180 9550 2200 9590
rect 2240 9550 2260 9590
rect 2180 9490 2260 9550
rect 2180 9450 2200 9490
rect 2240 9450 2260 9490
rect 2180 9420 2260 9450
rect 2490 9790 2590 9820
rect 2490 9750 2520 9790
rect 2560 9750 2590 9790
rect 2490 9690 2590 9750
rect 2490 9650 2520 9690
rect 2560 9650 2590 9690
rect 2490 9590 2590 9650
rect 2490 9550 2520 9590
rect 2560 9550 2590 9590
rect 2490 9490 2590 9550
rect 2490 9450 2520 9490
rect 2560 9450 2590 9490
rect 2490 9420 2590 9450
rect 2620 9790 2720 9820
rect 2620 9750 2650 9790
rect 2690 9750 2720 9790
rect 2620 9690 2720 9750
rect 2620 9650 2650 9690
rect 2690 9650 2720 9690
rect 2620 9590 2720 9650
rect 2620 9550 2650 9590
rect 2690 9550 2720 9590
rect 2620 9490 2720 9550
rect 2620 9450 2650 9490
rect 2690 9450 2720 9490
rect 2620 9420 2720 9450
rect 2880 9790 2980 9820
rect 2880 9750 2910 9790
rect 2950 9750 2980 9790
rect 2880 9690 2980 9750
rect 2880 9650 2910 9690
rect 2950 9650 2980 9690
rect 2880 9590 2980 9650
rect 2880 9550 2910 9590
rect 2950 9550 2980 9590
rect 2880 9490 2980 9550
rect 2880 9450 2910 9490
rect 2950 9450 2980 9490
rect 2880 9420 2980 9450
rect 3010 9790 3110 9820
rect 3010 9750 3040 9790
rect 3080 9750 3110 9790
rect 3010 9690 3110 9750
rect 3010 9650 3040 9690
rect 3080 9650 3110 9690
rect 3010 9590 3110 9650
rect 3010 9550 3040 9590
rect 3080 9550 3110 9590
rect 3010 9490 3110 9550
rect 3010 9450 3040 9490
rect 3080 9450 3110 9490
rect 3010 9420 3110 9450
rect 3270 9790 3370 9820
rect 3270 9750 3300 9790
rect 3340 9750 3370 9790
rect 3270 9690 3370 9750
rect 3270 9650 3300 9690
rect 3340 9650 3370 9690
rect 3270 9590 3370 9650
rect 3270 9550 3300 9590
rect 3340 9550 3370 9590
rect 3270 9490 3370 9550
rect 3270 9450 3300 9490
rect 3340 9450 3370 9490
rect 3270 9420 3370 9450
rect 3400 9790 3500 9820
rect 3400 9750 3430 9790
rect 3470 9750 3500 9790
rect 3400 9690 3500 9750
rect 3400 9650 3430 9690
rect 3470 9650 3500 9690
rect 3400 9590 3500 9650
rect 3400 9550 3430 9590
rect 3470 9550 3500 9590
rect 3400 9490 3500 9550
rect 3400 9450 3430 9490
rect 3470 9450 3500 9490
rect 3400 9420 3500 9450
rect 3560 9790 3660 9820
rect 3560 9750 3590 9790
rect 3630 9750 3660 9790
rect 3560 9690 3660 9750
rect 3560 9650 3590 9690
rect 3630 9650 3660 9690
rect 3560 9590 3660 9650
rect 3560 9550 3590 9590
rect 3630 9550 3660 9590
rect 3560 9490 3660 9550
rect 3560 9450 3590 9490
rect 3630 9450 3660 9490
rect 3560 9420 3660 9450
rect 3690 9790 3790 9820
rect 3690 9750 3720 9790
rect 3760 9750 3790 9790
rect 3690 9690 3790 9750
rect 3690 9650 3720 9690
rect 3760 9650 3790 9690
rect 3690 9590 3790 9650
rect 3690 9550 3720 9590
rect 3760 9550 3790 9590
rect 3690 9490 3790 9550
rect 3690 9450 3720 9490
rect 3760 9450 3790 9490
rect 3690 9420 3790 9450
rect 3950 9790 4050 9820
rect 3950 9750 3980 9790
rect 4020 9750 4050 9790
rect 3950 9690 4050 9750
rect 3950 9650 3980 9690
rect 4020 9650 4050 9690
rect 3950 9590 4050 9650
rect 3950 9550 3980 9590
rect 4020 9550 4050 9590
rect 3950 9490 4050 9550
rect 3950 9450 3980 9490
rect 4020 9450 4050 9490
rect 3950 9420 4050 9450
rect 4080 9790 4180 9820
rect 4080 9750 4110 9790
rect 4150 9750 4180 9790
rect 4080 9690 4180 9750
rect 4080 9650 4110 9690
rect 4150 9650 4180 9690
rect 4080 9590 4180 9650
rect 4080 9550 4110 9590
rect 4150 9550 4180 9590
rect 4080 9490 4180 9550
rect 4080 9450 4110 9490
rect 4150 9450 4180 9490
rect 4080 9420 4180 9450
rect 5640 9760 5740 9790
rect 5640 9720 5670 9760
rect 5710 9720 5740 9760
rect 5640 9660 5740 9720
rect 5640 9620 5670 9660
rect 5710 9620 5740 9660
rect 5640 9560 5740 9620
rect 5640 9520 5670 9560
rect 5710 9520 5740 9560
rect 5640 9460 5740 9520
rect 5640 9420 5670 9460
rect 5710 9420 5740 9460
rect 5640 9390 5740 9420
rect 5860 9760 5960 9790
rect 5860 9720 5890 9760
rect 5930 9720 5960 9760
rect 5860 9660 5960 9720
rect 5860 9620 5890 9660
rect 5930 9620 5960 9660
rect 5860 9560 5960 9620
rect 5860 9520 5890 9560
rect 5930 9520 5960 9560
rect 5860 9460 5960 9520
rect 5860 9420 5890 9460
rect 5930 9420 5960 9460
rect 5860 9390 5960 9420
rect 6080 9760 6180 9790
rect 6080 9720 6110 9760
rect 6150 9720 6180 9760
rect 6080 9660 6180 9720
rect 6080 9620 6110 9660
rect 6150 9620 6180 9660
rect 6080 9560 6180 9620
rect 6080 9520 6110 9560
rect 6150 9520 6180 9560
rect 6080 9460 6180 9520
rect 6080 9420 6110 9460
rect 6150 9420 6180 9460
rect 6080 9390 6180 9420
rect 6300 9760 6400 9790
rect 6300 9720 6330 9760
rect 6370 9720 6400 9760
rect 6300 9660 6400 9720
rect 6300 9620 6330 9660
rect 6370 9620 6400 9660
rect 6300 9560 6400 9620
rect 6300 9520 6330 9560
rect 6370 9520 6400 9560
rect 6300 9460 6400 9520
rect 6300 9420 6330 9460
rect 6370 9420 6400 9460
rect 6300 9390 6400 9420
rect 6520 9760 6620 9790
rect 6520 9720 6550 9760
rect 6590 9720 6620 9760
rect 6520 9660 6620 9720
rect 6520 9620 6550 9660
rect 6590 9620 6620 9660
rect 6520 9560 6620 9620
rect 6520 9520 6550 9560
rect 6590 9520 6620 9560
rect 6520 9460 6620 9520
rect 6520 9420 6550 9460
rect 6590 9420 6620 9460
rect 6520 9390 6620 9420
rect 6740 9760 6840 9790
rect 6740 9720 6770 9760
rect 6810 9720 6840 9760
rect 6740 9660 6840 9720
rect 6740 9620 6770 9660
rect 6810 9620 6840 9660
rect 6740 9560 6840 9620
rect 6740 9520 6770 9560
rect 6810 9520 6840 9560
rect 6740 9460 6840 9520
rect 6740 9420 6770 9460
rect 6810 9420 6840 9460
rect 6740 9390 6840 9420
rect 6960 9760 7060 9790
rect 7160 9760 7260 9790
rect 6960 9720 6990 9760
rect 7030 9720 7060 9760
rect 7160 9720 7190 9760
rect 7230 9720 7260 9760
rect 6960 9660 7060 9720
rect 7160 9660 7260 9720
rect 6960 9620 6990 9660
rect 7030 9620 7060 9660
rect 7160 9620 7190 9660
rect 7230 9620 7260 9660
rect 6960 9560 7060 9620
rect 7160 9560 7260 9620
rect 6960 9520 6990 9560
rect 7030 9520 7060 9560
rect 7160 9520 7190 9560
rect 7230 9520 7260 9560
rect 6960 9460 7060 9520
rect 7160 9460 7260 9520
rect 6960 9420 6990 9460
rect 7030 9420 7060 9460
rect 7160 9420 7190 9460
rect 7230 9420 7260 9460
rect 6960 9390 7060 9420
rect 7160 9390 7260 9420
rect 7380 9760 7480 9790
rect 7380 9720 7410 9760
rect 7450 9720 7480 9760
rect 7380 9660 7480 9720
rect 7380 9620 7410 9660
rect 7450 9620 7480 9660
rect 7380 9560 7480 9620
rect 7380 9520 7410 9560
rect 7450 9520 7480 9560
rect 7380 9460 7480 9520
rect 7380 9420 7410 9460
rect 7450 9420 7480 9460
rect 7380 9390 7480 9420
rect 7600 9760 7700 9790
rect 7600 9720 7630 9760
rect 7670 9720 7700 9760
rect 7600 9660 7700 9720
rect 7600 9620 7630 9660
rect 7670 9620 7700 9660
rect 7600 9560 7700 9620
rect 7600 9520 7630 9560
rect 7670 9520 7700 9560
rect 7600 9460 7700 9520
rect 7600 9420 7630 9460
rect 7670 9420 7700 9460
rect 7600 9390 7700 9420
rect 7820 9760 7920 9790
rect 7820 9720 7850 9760
rect 7890 9720 7920 9760
rect 7820 9660 7920 9720
rect 7820 9620 7850 9660
rect 7890 9620 7920 9660
rect 7820 9560 7920 9620
rect 7820 9520 7850 9560
rect 7890 9520 7920 9560
rect 7820 9460 7920 9520
rect 7820 9420 7850 9460
rect 7890 9420 7920 9460
rect 7820 9390 7920 9420
rect 8040 9760 8140 9790
rect 8040 9720 8070 9760
rect 8110 9720 8140 9760
rect 8040 9660 8140 9720
rect 8040 9620 8070 9660
rect 8110 9620 8140 9660
rect 8040 9560 8140 9620
rect 8040 9520 8070 9560
rect 8110 9520 8140 9560
rect 8040 9460 8140 9520
rect 8040 9420 8070 9460
rect 8110 9420 8140 9460
rect 8040 9390 8140 9420
rect 8260 9760 8360 9790
rect 8260 9720 8290 9760
rect 8330 9720 8360 9760
rect 8260 9660 8360 9720
rect 8260 9620 8290 9660
rect 8330 9620 8360 9660
rect 8260 9560 8360 9620
rect 8260 9520 8290 9560
rect 8330 9520 8360 9560
rect 8260 9460 8360 9520
rect 8260 9420 8290 9460
rect 8330 9420 8360 9460
rect 8260 9390 8360 9420
rect 8480 9760 8580 9790
rect 8480 9720 8510 9760
rect 8550 9720 8580 9760
rect 8480 9660 8580 9720
rect 8480 9620 8510 9660
rect 8550 9620 8580 9660
rect 8480 9560 8580 9620
rect 8480 9520 8510 9560
rect 8550 9520 8580 9560
rect 8480 9460 8580 9520
rect 8480 9420 8510 9460
rect 8550 9420 8580 9460
rect 8480 9390 8580 9420
rect -640 9030 -560 9060
rect -640 8990 -620 9030
rect -580 8990 -560 9030
rect -640 8930 -560 8990
rect -640 8890 -620 8930
rect -580 8890 -560 8930
rect -640 8830 -560 8890
rect -640 8790 -620 8830
rect -580 8790 -560 8830
rect -640 8730 -560 8790
rect -640 8690 -620 8730
rect -580 8690 -560 8730
rect -640 8660 -560 8690
rect -530 9030 -450 9060
rect -530 8990 -510 9030
rect -470 8990 -450 9030
rect -530 8930 -450 8990
rect -530 8890 -510 8930
rect -470 8890 -450 8930
rect -530 8830 -450 8890
rect -530 8790 -510 8830
rect -470 8790 -450 8830
rect -530 8730 -450 8790
rect -530 8690 -510 8730
rect -470 8690 -450 8730
rect -530 8660 -450 8690
rect -420 9030 -340 9060
rect -420 8990 -400 9030
rect -360 8990 -340 9030
rect -420 8930 -340 8990
rect -420 8890 -400 8930
rect -360 8890 -340 8930
rect -420 8830 -340 8890
rect -420 8790 -400 8830
rect -360 8790 -340 8830
rect -420 8730 -340 8790
rect -420 8690 -400 8730
rect -360 8690 -340 8730
rect -420 8660 -340 8690
rect -120 9030 -40 9060
rect -120 8990 -100 9030
rect -60 8990 -40 9030
rect -120 8930 -40 8990
rect -120 8890 -100 8930
rect -60 8890 -40 8930
rect -120 8830 -40 8890
rect -120 8790 -100 8830
rect -60 8790 -40 8830
rect -120 8730 -40 8790
rect -120 8690 -100 8730
rect -60 8690 -40 8730
rect -120 8660 -40 8690
rect -10 9030 70 9060
rect -10 8990 10 9030
rect 50 8990 70 9030
rect -10 8930 70 8990
rect -10 8890 10 8930
rect 50 8890 70 8930
rect -10 8830 70 8890
rect -10 8790 10 8830
rect 50 8790 70 8830
rect -10 8730 70 8790
rect -10 8690 10 8730
rect 50 8690 70 8730
rect -10 8660 70 8690
rect 100 9030 180 9060
rect 260 9030 340 9060
rect 100 8990 120 9030
rect 160 8990 180 9030
rect 260 8990 280 9030
rect 320 8990 340 9030
rect 100 8930 180 8990
rect 260 8930 340 8990
rect 100 8890 120 8930
rect 160 8890 180 8930
rect 260 8890 280 8930
rect 320 8890 340 8930
rect 100 8830 180 8890
rect 260 8830 340 8890
rect 100 8790 120 8830
rect 160 8790 180 8830
rect 260 8790 280 8830
rect 320 8790 340 8830
rect 100 8730 180 8790
rect 260 8730 340 8790
rect 100 8690 120 8730
rect 160 8690 180 8730
rect 260 8690 280 8730
rect 320 8690 340 8730
rect 100 8660 180 8690
rect 260 8660 340 8690
rect 370 9030 450 9060
rect 370 8990 390 9030
rect 430 8990 450 9030
rect 370 8930 450 8990
rect 370 8890 390 8930
rect 430 8890 450 8930
rect 370 8830 450 8890
rect 370 8790 390 8830
rect 430 8790 450 8830
rect 370 8730 450 8790
rect 370 8690 390 8730
rect 430 8690 450 8730
rect 370 8660 450 8690
rect 480 9030 560 9060
rect 480 8990 500 9030
rect 540 8990 560 9030
rect 480 8930 560 8990
rect 480 8890 500 8930
rect 540 8890 560 8930
rect 480 8830 560 8890
rect 480 8790 500 8830
rect 540 8790 560 8830
rect 480 8730 560 8790
rect 480 8690 500 8730
rect 540 8690 560 8730
rect 480 8660 560 8690
rect 780 9030 860 9060
rect 780 8990 800 9030
rect 840 8990 860 9030
rect 780 8930 860 8990
rect 780 8890 800 8930
rect 840 8890 860 8930
rect 780 8830 860 8890
rect 780 8790 800 8830
rect 840 8790 860 8830
rect 780 8730 860 8790
rect 780 8690 800 8730
rect 840 8690 860 8730
rect 780 8660 860 8690
rect 890 9030 970 9060
rect 890 8990 910 9030
rect 950 8990 970 9030
rect 890 8930 970 8990
rect 890 8890 910 8930
rect 950 8890 970 8930
rect 890 8830 970 8890
rect 890 8790 910 8830
rect 950 8790 970 8830
rect 890 8730 970 8790
rect 890 8690 910 8730
rect 950 8690 970 8730
rect 890 8660 970 8690
rect 1000 9030 1080 9060
rect 1000 8990 1020 9030
rect 1060 8990 1080 9030
rect 1000 8930 1080 8990
rect 1000 8890 1020 8930
rect 1060 8890 1080 8930
rect 1000 8830 1080 8890
rect 1000 8790 1020 8830
rect 1060 8790 1080 8830
rect 1000 8730 1080 8790
rect 1000 8690 1020 8730
rect 1060 8690 1080 8730
rect 1000 8660 1080 8690
rect 1290 9030 1370 9060
rect 1290 8990 1310 9030
rect 1350 8990 1370 9030
rect 1290 8930 1370 8990
rect 1290 8890 1310 8930
rect 1350 8890 1370 8930
rect 1290 8830 1370 8890
rect 1290 8790 1310 8830
rect 1350 8790 1370 8830
rect 1290 8730 1370 8790
rect 1290 8690 1310 8730
rect 1350 8690 1370 8730
rect 1290 8660 1370 8690
rect 1400 9030 1480 9060
rect 1400 8990 1420 9030
rect 1460 8990 1480 9030
rect 1400 8930 1480 8990
rect 1400 8890 1420 8930
rect 1460 8890 1480 8930
rect 1400 8830 1480 8890
rect 1400 8790 1420 8830
rect 1460 8790 1480 8830
rect 1400 8730 1480 8790
rect 1400 8690 1420 8730
rect 1460 8690 1480 8730
rect 1400 8660 1480 8690
rect 1620 9030 1700 9060
rect 1620 8990 1640 9030
rect 1680 8990 1700 9030
rect 1620 8930 1700 8990
rect 1620 8890 1640 8930
rect 1680 8890 1700 8930
rect 1620 8830 1700 8890
rect 1620 8790 1640 8830
rect 1680 8790 1700 8830
rect 1620 8730 1700 8790
rect 1620 8690 1640 8730
rect 1680 8690 1700 8730
rect 1620 8660 1700 8690
rect 1730 9030 1810 9060
rect 1730 8990 1750 9030
rect 1790 8990 1810 9030
rect 1730 8930 1810 8990
rect 1730 8890 1750 8930
rect 1790 8890 1810 8930
rect 1730 8830 1810 8890
rect 1730 8790 1750 8830
rect 1790 8790 1810 8830
rect 1730 8730 1810 8790
rect 1730 8690 1750 8730
rect 1790 8690 1810 8730
rect 1730 8660 1810 8690
rect 1950 9030 2030 9060
rect 1950 8990 1970 9030
rect 2010 8990 2030 9030
rect 1950 8930 2030 8990
rect 1950 8890 1970 8930
rect 2010 8890 2030 8930
rect 1950 8830 2030 8890
rect 1950 8790 1970 8830
rect 2010 8790 2030 8830
rect 1950 8730 2030 8790
rect 1950 8690 1970 8730
rect 2010 8690 2030 8730
rect 1950 8660 2030 8690
rect 2060 9030 2140 9060
rect 2060 8990 2080 9030
rect 2120 8990 2140 9030
rect 2060 8930 2140 8990
rect 2060 8890 2080 8930
rect 2120 8890 2140 8930
rect 2060 8830 2140 8890
rect 2060 8790 2080 8830
rect 2120 8790 2140 8830
rect 2060 8730 2140 8790
rect 2060 8690 2080 8730
rect 2120 8690 2140 8730
rect 2060 8660 2140 8690
rect 2490 9030 2590 9060
rect 2490 8990 2520 9030
rect 2560 8990 2590 9030
rect 2490 8930 2590 8990
rect 2490 8890 2520 8930
rect 2560 8890 2590 8930
rect 2490 8830 2590 8890
rect 2490 8790 2520 8830
rect 2560 8790 2590 8830
rect 2490 8730 2590 8790
rect 2490 8690 2520 8730
rect 2560 8690 2590 8730
rect 2490 8660 2590 8690
rect 2620 9030 2720 9060
rect 2620 8990 2650 9030
rect 2690 8990 2720 9030
rect 2620 8930 2720 8990
rect 2620 8890 2650 8930
rect 2690 8890 2720 8930
rect 2620 8830 2720 8890
rect 2620 8790 2650 8830
rect 2690 8790 2720 8830
rect 2620 8730 2720 8790
rect 2620 8690 2650 8730
rect 2690 8690 2720 8730
rect 2620 8660 2720 8690
rect 2880 9030 2980 9060
rect 2880 8990 2910 9030
rect 2950 8990 2980 9030
rect 2880 8930 2980 8990
rect 2880 8890 2910 8930
rect 2950 8890 2980 8930
rect 2880 8830 2980 8890
rect 2880 8790 2910 8830
rect 2950 8790 2980 8830
rect 2880 8730 2980 8790
rect 2880 8690 2910 8730
rect 2950 8690 2980 8730
rect 2880 8660 2980 8690
rect 3010 9030 3110 9060
rect 3010 8990 3040 9030
rect 3080 8990 3110 9030
rect 3010 8930 3110 8990
rect 3010 8890 3040 8930
rect 3080 8890 3110 8930
rect 3010 8830 3110 8890
rect 3010 8790 3040 8830
rect 3080 8790 3110 8830
rect 3010 8730 3110 8790
rect 3010 8690 3040 8730
rect 3080 8690 3110 8730
rect 3010 8660 3110 8690
rect 3270 9030 3370 9060
rect 3270 8990 3300 9030
rect 3340 8990 3370 9030
rect 3270 8930 3370 8990
rect 3270 8890 3300 8930
rect 3340 8890 3370 8930
rect 3270 8830 3370 8890
rect 3270 8790 3300 8830
rect 3340 8790 3370 8830
rect 3270 8730 3370 8790
rect 3270 8690 3300 8730
rect 3340 8690 3370 8730
rect 3270 8660 3370 8690
rect 3400 9030 3500 9060
rect 3400 8990 3430 9030
rect 3470 8990 3500 9030
rect 3400 8930 3500 8990
rect 3400 8890 3430 8930
rect 3470 8890 3500 8930
rect 3400 8830 3500 8890
rect 3400 8790 3430 8830
rect 3470 8790 3500 8830
rect 3400 8730 3500 8790
rect 3400 8690 3430 8730
rect 3470 8690 3500 8730
rect 3400 8660 3500 8690
rect 3560 9030 3660 9060
rect 3560 8990 3590 9030
rect 3630 8990 3660 9030
rect 3560 8930 3660 8990
rect 3560 8890 3590 8930
rect 3630 8890 3660 8930
rect 3560 8830 3660 8890
rect 3560 8790 3590 8830
rect 3630 8790 3660 8830
rect 3560 8730 3660 8790
rect 3560 8690 3590 8730
rect 3630 8690 3660 8730
rect 3560 8660 3660 8690
rect 3690 9030 3790 9060
rect 3690 8990 3720 9030
rect 3760 8990 3790 9030
rect 3690 8930 3790 8990
rect 3690 8890 3720 8930
rect 3760 8890 3790 8930
rect 3690 8830 3790 8890
rect 3690 8790 3720 8830
rect 3760 8790 3790 8830
rect 3690 8730 3790 8790
rect 3690 8690 3720 8730
rect 3760 8690 3790 8730
rect 3690 8660 3790 8690
rect -1360 6840 -1280 6870
rect -1360 6800 -1340 6840
rect -1300 6800 -1280 6840
rect -1360 6740 -1280 6800
rect -1360 6700 -1340 6740
rect -1300 6700 -1280 6740
rect -1360 6670 -1280 6700
rect -1250 6840 -1170 6870
rect -1250 6800 -1230 6840
rect -1190 6800 -1170 6840
rect -1250 6740 -1170 6800
rect -1250 6700 -1230 6740
rect -1190 6700 -1170 6740
rect -1250 6670 -1170 6700
rect -1140 6840 -1060 6870
rect -1140 6800 -1120 6840
rect -1080 6800 -1060 6840
rect -1140 6740 -1060 6800
rect -1140 6700 -1120 6740
rect -1080 6700 -1060 6740
rect -1140 6670 -1060 6700
rect -1030 6840 -950 6870
rect -1030 6800 -1010 6840
rect -970 6800 -950 6840
rect -1030 6740 -950 6800
rect -1030 6700 -1010 6740
rect -970 6700 -950 6740
rect -1030 6670 -950 6700
rect -920 6840 -840 6870
rect -920 6800 -900 6840
rect -860 6800 -840 6840
rect -920 6740 -840 6800
rect -920 6700 -900 6740
rect -860 6700 -840 6740
rect -920 6670 -840 6700
rect -810 6840 -730 6870
rect -810 6800 -790 6840
rect -750 6800 -730 6840
rect -810 6740 -730 6800
rect -810 6700 -790 6740
rect -750 6700 -730 6740
rect -810 6670 -730 6700
rect -700 6840 -620 6870
rect -700 6800 -680 6840
rect -640 6800 -620 6840
rect -700 6740 -620 6800
rect -700 6700 -680 6740
rect -640 6700 -620 6740
rect -700 6670 -620 6700
rect -590 6840 -510 6870
rect -590 6800 -570 6840
rect -530 6800 -510 6840
rect -590 6740 -510 6800
rect -590 6700 -570 6740
rect -530 6700 -510 6740
rect -590 6670 -510 6700
rect -480 6840 -400 6870
rect -480 6800 -460 6840
rect -420 6800 -400 6840
rect -480 6740 -400 6800
rect -480 6700 -460 6740
rect -420 6700 -400 6740
rect -480 6670 -400 6700
rect -370 6840 -290 6870
rect -370 6800 -350 6840
rect -310 6800 -290 6840
rect -370 6740 -290 6800
rect -370 6700 -350 6740
rect -310 6700 -290 6740
rect -370 6670 -290 6700
rect -260 6840 -180 6870
rect -260 6800 -240 6840
rect -200 6800 -180 6840
rect -260 6740 -180 6800
rect -260 6700 -240 6740
rect -200 6700 -180 6740
rect -260 6670 -180 6700
rect -150 6840 -70 6870
rect -150 6800 -130 6840
rect -90 6800 -70 6840
rect -150 6740 -70 6800
rect -150 6700 -130 6740
rect -90 6700 -70 6740
rect -150 6670 -70 6700
rect -40 6840 40 6870
rect -40 6800 -20 6840
rect 20 6800 40 6840
rect -40 6740 40 6800
rect -40 6700 -20 6740
rect 20 6700 40 6740
rect -40 6670 40 6700
rect 540 6840 620 6870
rect 540 6800 560 6840
rect 600 6800 620 6840
rect 540 6740 620 6800
rect 540 6700 560 6740
rect 600 6700 620 6740
rect 540 6670 620 6700
rect 650 6840 730 6870
rect 650 6800 670 6840
rect 710 6800 730 6840
rect 650 6740 730 6800
rect 650 6700 670 6740
rect 710 6700 730 6740
rect 650 6670 730 6700
rect 760 6840 840 6870
rect 760 6800 780 6840
rect 820 6800 840 6840
rect 760 6740 840 6800
rect 760 6700 780 6740
rect 820 6700 840 6740
rect 760 6670 840 6700
rect 870 6840 950 6870
rect 870 6800 890 6840
rect 930 6800 950 6840
rect 870 6740 950 6800
rect 870 6700 890 6740
rect 930 6700 950 6740
rect 870 6670 950 6700
rect 980 6840 1060 6870
rect 980 6800 1000 6840
rect 1040 6800 1060 6840
rect 980 6740 1060 6800
rect 980 6700 1000 6740
rect 1040 6700 1060 6740
rect 980 6670 1060 6700
rect 1090 6840 1170 6870
rect 1090 6800 1110 6840
rect 1150 6800 1170 6840
rect 1090 6740 1170 6800
rect 1090 6700 1110 6740
rect 1150 6700 1170 6740
rect 1090 6670 1170 6700
rect 1200 6840 1280 6870
rect 1200 6800 1220 6840
rect 1260 6800 1280 6840
rect 1200 6740 1280 6800
rect 1200 6700 1220 6740
rect 1260 6700 1280 6740
rect 1200 6670 1280 6700
rect 1310 6840 1390 6870
rect 1310 6800 1330 6840
rect 1370 6800 1390 6840
rect 1310 6740 1390 6800
rect 1310 6700 1330 6740
rect 1370 6700 1390 6740
rect 1310 6670 1390 6700
rect 1420 6840 1500 6870
rect 1420 6800 1440 6840
rect 1480 6800 1500 6840
rect 1420 6740 1500 6800
rect 1420 6700 1440 6740
rect 1480 6700 1500 6740
rect 1420 6670 1500 6700
rect 1530 6840 1610 6870
rect 1530 6800 1550 6840
rect 1590 6800 1610 6840
rect 1530 6740 1610 6800
rect 1530 6700 1550 6740
rect 1590 6700 1610 6740
rect 1530 6670 1610 6700
rect 1640 6840 1720 6870
rect 1640 6800 1660 6840
rect 1700 6800 1720 6840
rect 1640 6740 1720 6800
rect 1640 6700 1660 6740
rect 1700 6700 1720 6740
rect 1640 6670 1720 6700
rect 1750 6840 1830 6870
rect 1750 6800 1770 6840
rect 1810 6800 1830 6840
rect 1750 6740 1830 6800
rect 1750 6700 1770 6740
rect 1810 6700 1830 6740
rect 1750 6670 1830 6700
rect 1860 6840 1940 6870
rect 1860 6800 1880 6840
rect 1920 6800 1940 6840
rect 1860 6740 1940 6800
rect 1860 6700 1880 6740
rect 1920 6700 1940 6740
rect 1860 6670 1940 6700
rect -1370 6240 -1290 6270
rect -1370 6200 -1350 6240
rect -1310 6200 -1290 6240
rect -1370 6140 -1290 6200
rect -1370 6100 -1350 6140
rect -1310 6100 -1290 6140
rect -1370 6040 -1290 6100
rect -1370 6000 -1350 6040
rect -1310 6000 -1290 6040
rect -1370 5940 -1290 6000
rect -1370 5900 -1350 5940
rect -1310 5900 -1290 5940
rect -1370 5840 -1290 5900
rect -1370 5800 -1350 5840
rect -1310 5800 -1290 5840
rect -1370 5740 -1290 5800
rect -1370 5700 -1350 5740
rect -1310 5700 -1290 5740
rect -1370 5670 -1290 5700
rect -1190 6240 -1110 6270
rect -1190 6200 -1170 6240
rect -1130 6200 -1110 6240
rect -1190 6140 -1110 6200
rect -1190 6100 -1170 6140
rect -1130 6100 -1110 6140
rect -1190 6040 -1110 6100
rect -1190 6000 -1170 6040
rect -1130 6000 -1110 6040
rect -1190 5940 -1110 6000
rect -1190 5900 -1170 5940
rect -1130 5900 -1110 5940
rect -1190 5840 -1110 5900
rect -1190 5800 -1170 5840
rect -1130 5800 -1110 5840
rect -1190 5740 -1110 5800
rect -1190 5700 -1170 5740
rect -1130 5700 -1110 5740
rect -1190 5670 -1110 5700
rect -1010 6240 -930 6270
rect -1010 6200 -990 6240
rect -950 6200 -930 6240
rect -1010 6140 -930 6200
rect -1010 6100 -990 6140
rect -950 6100 -930 6140
rect -1010 6040 -930 6100
rect -1010 6000 -990 6040
rect -950 6000 -930 6040
rect -1010 5940 -930 6000
rect -1010 5900 -990 5940
rect -950 5900 -930 5940
rect -1010 5840 -930 5900
rect -1010 5800 -990 5840
rect -950 5800 -930 5840
rect -1010 5740 -930 5800
rect -1010 5700 -990 5740
rect -950 5700 -930 5740
rect -1010 5670 -930 5700
rect -830 6240 -750 6270
rect -830 6200 -810 6240
rect -770 6200 -750 6240
rect -830 6140 -750 6200
rect -830 6100 -810 6140
rect -770 6100 -750 6140
rect -830 6040 -750 6100
rect -830 6000 -810 6040
rect -770 6000 -750 6040
rect -830 5940 -750 6000
rect -830 5900 -810 5940
rect -770 5900 -750 5940
rect -830 5840 -750 5900
rect -830 5800 -810 5840
rect -770 5800 -750 5840
rect -830 5740 -750 5800
rect -830 5700 -810 5740
rect -770 5700 -750 5740
rect -830 5670 -750 5700
rect -650 6240 -570 6270
rect -650 6200 -630 6240
rect -590 6200 -570 6240
rect -650 6140 -570 6200
rect -650 6100 -630 6140
rect -590 6100 -570 6140
rect -650 6040 -570 6100
rect -650 6000 -630 6040
rect -590 6000 -570 6040
rect -650 5940 -570 6000
rect -650 5900 -630 5940
rect -590 5900 -570 5940
rect -650 5840 -570 5900
rect -650 5800 -630 5840
rect -590 5800 -570 5840
rect -650 5740 -570 5800
rect -650 5700 -630 5740
rect -590 5700 -570 5740
rect -650 5670 -570 5700
rect -470 6240 -390 6270
rect -470 6200 -450 6240
rect -410 6200 -390 6240
rect -470 6140 -390 6200
rect -470 6100 -450 6140
rect -410 6100 -390 6140
rect -470 6040 -390 6100
rect -470 6000 -450 6040
rect -410 6000 -390 6040
rect -470 5940 -390 6000
rect -470 5900 -450 5940
rect -410 5900 -390 5940
rect -470 5840 -390 5900
rect -470 5800 -450 5840
rect -410 5800 -390 5840
rect -470 5740 -390 5800
rect -470 5700 -450 5740
rect -410 5700 -390 5740
rect -470 5670 -390 5700
rect -290 6240 -210 6270
rect -290 6200 -270 6240
rect -230 6200 -210 6240
rect -290 6140 -210 6200
rect -290 6100 -270 6140
rect -230 6100 -210 6140
rect -290 6040 -210 6100
rect -290 6000 -270 6040
rect -230 6000 -210 6040
rect -290 5940 -210 6000
rect -290 5900 -270 5940
rect -230 5900 -210 5940
rect -290 5840 -210 5900
rect -290 5800 -270 5840
rect -230 5800 -210 5840
rect -290 5740 -210 5800
rect -290 5700 -270 5740
rect -230 5700 -210 5740
rect -290 5670 -210 5700
rect -110 6240 -30 6270
rect -110 6200 -90 6240
rect -50 6200 -30 6240
rect -110 6140 -30 6200
rect -110 6100 -90 6140
rect -50 6100 -30 6140
rect -110 6040 -30 6100
rect -110 6000 -90 6040
rect -50 6000 -30 6040
rect -110 5940 -30 6000
rect -110 5900 -90 5940
rect -50 5900 -30 5940
rect -110 5840 -30 5900
rect -110 5800 -90 5840
rect -50 5800 -30 5840
rect -110 5740 -30 5800
rect -110 5700 -90 5740
rect -50 5700 -30 5740
rect -110 5670 -30 5700
rect 70 6240 150 6270
rect 70 6200 90 6240
rect 130 6200 150 6240
rect 70 6140 150 6200
rect 70 6100 90 6140
rect 130 6100 150 6140
rect 70 6040 150 6100
rect 70 6000 90 6040
rect 130 6000 150 6040
rect 70 5940 150 6000
rect 70 5900 90 5940
rect 130 5900 150 5940
rect 70 5840 150 5900
rect 70 5800 90 5840
rect 130 5800 150 5840
rect 70 5740 150 5800
rect 70 5700 90 5740
rect 130 5700 150 5740
rect 70 5670 150 5700
rect 250 6240 330 6270
rect 250 6200 270 6240
rect 310 6200 330 6240
rect 250 6140 330 6200
rect 250 6100 270 6140
rect 310 6100 330 6140
rect 250 6040 330 6100
rect 250 6000 270 6040
rect 310 6000 330 6040
rect 250 5940 330 6000
rect 250 5900 270 5940
rect 310 5900 330 5940
rect 250 5840 330 5900
rect 250 5800 270 5840
rect 310 5800 330 5840
rect 250 5740 330 5800
rect 250 5700 270 5740
rect 310 5700 330 5740
rect 250 5670 330 5700
rect 430 6240 510 6270
rect 430 6200 450 6240
rect 490 6200 510 6240
rect 430 6140 510 6200
rect 430 6100 450 6140
rect 490 6100 510 6140
rect 430 6040 510 6100
rect 430 6000 450 6040
rect 490 6000 510 6040
rect 430 5940 510 6000
rect 430 5900 450 5940
rect 490 5900 510 5940
rect 430 5840 510 5900
rect 430 5800 450 5840
rect 490 5800 510 5840
rect 430 5740 510 5800
rect 430 5700 450 5740
rect 490 5700 510 5740
rect 430 5670 510 5700
rect 610 6240 690 6270
rect 610 6200 630 6240
rect 670 6200 690 6240
rect 610 6140 690 6200
rect 610 6100 630 6140
rect 670 6100 690 6140
rect 610 6040 690 6100
rect 610 6000 630 6040
rect 670 6000 690 6040
rect 610 5940 690 6000
rect 610 5900 630 5940
rect 670 5900 690 5940
rect 610 5840 690 5900
rect 610 5800 630 5840
rect 670 5800 690 5840
rect 610 5740 690 5800
rect 610 5700 630 5740
rect 670 5700 690 5740
rect 610 5670 690 5700
rect 790 6240 870 6270
rect 790 6200 810 6240
rect 850 6200 870 6240
rect 790 6140 870 6200
rect 790 6100 810 6140
rect 850 6100 870 6140
rect 790 6040 870 6100
rect 790 6000 810 6040
rect 850 6000 870 6040
rect 790 5940 870 6000
rect 790 5900 810 5940
rect 850 5900 870 5940
rect 790 5840 870 5900
rect 790 5800 810 5840
rect 850 5800 870 5840
rect 790 5740 870 5800
rect 790 5700 810 5740
rect 850 5700 870 5740
rect 790 5670 870 5700
rect 970 6240 1050 6270
rect 970 6200 990 6240
rect 1030 6200 1050 6240
rect 970 6140 1050 6200
rect 970 6100 990 6140
rect 1030 6100 1050 6140
rect 970 6040 1050 6100
rect 970 6000 990 6040
rect 1030 6000 1050 6040
rect 970 5940 1050 6000
rect 970 5900 990 5940
rect 1030 5900 1050 5940
rect 970 5840 1050 5900
rect 970 5800 990 5840
rect 1030 5800 1050 5840
rect 970 5740 1050 5800
rect 970 5700 990 5740
rect 1030 5700 1050 5740
rect 970 5670 1050 5700
rect 1150 6240 1230 6270
rect 1150 6200 1170 6240
rect 1210 6200 1230 6240
rect 1150 6140 1230 6200
rect 1150 6100 1170 6140
rect 1210 6100 1230 6140
rect 1150 6040 1230 6100
rect 1150 6000 1170 6040
rect 1210 6000 1230 6040
rect 1150 5940 1230 6000
rect 1150 5900 1170 5940
rect 1210 5900 1230 5940
rect 1150 5840 1230 5900
rect 1150 5800 1170 5840
rect 1210 5800 1230 5840
rect 1150 5740 1230 5800
rect 1150 5700 1170 5740
rect 1210 5700 1230 5740
rect 1150 5670 1230 5700
rect 1330 6240 1410 6270
rect 1330 6200 1350 6240
rect 1390 6200 1410 6240
rect 1330 6140 1410 6200
rect 1330 6100 1350 6140
rect 1390 6100 1410 6140
rect 1330 6040 1410 6100
rect 1330 6000 1350 6040
rect 1390 6000 1410 6040
rect 1330 5940 1410 6000
rect 1330 5900 1350 5940
rect 1390 5900 1410 5940
rect 1330 5840 1410 5900
rect 1330 5800 1350 5840
rect 1390 5800 1410 5840
rect 1330 5740 1410 5800
rect 1330 5700 1350 5740
rect 1390 5700 1410 5740
rect 1330 5670 1410 5700
rect 1510 6240 1590 6270
rect 1510 6200 1530 6240
rect 1570 6200 1590 6240
rect 1510 6140 1590 6200
rect 1510 6100 1530 6140
rect 1570 6100 1590 6140
rect 1510 6040 1590 6100
rect 1510 6000 1530 6040
rect 1570 6000 1590 6040
rect 1510 5940 1590 6000
rect 1510 5900 1530 5940
rect 1570 5900 1590 5940
rect 1510 5840 1590 5900
rect 1510 5800 1530 5840
rect 1570 5800 1590 5840
rect 1510 5740 1590 5800
rect 1510 5700 1530 5740
rect 1570 5700 1590 5740
rect 1510 5670 1590 5700
rect 1690 6240 1770 6270
rect 1690 6200 1710 6240
rect 1750 6200 1770 6240
rect 1690 6140 1770 6200
rect 1690 6100 1710 6140
rect 1750 6100 1770 6140
rect 1690 6040 1770 6100
rect 1690 6000 1710 6040
rect 1750 6000 1770 6040
rect 1690 5940 1770 6000
rect 1690 5900 1710 5940
rect 1750 5900 1770 5940
rect 1690 5840 1770 5900
rect 1690 5800 1710 5840
rect 1750 5800 1770 5840
rect 1690 5740 1770 5800
rect 1690 5700 1710 5740
rect 1750 5700 1770 5740
rect 1690 5670 1770 5700
rect 1870 6240 1950 6270
rect 1870 6200 1890 6240
rect 1930 6200 1950 6240
rect 1870 6140 1950 6200
rect 1870 6100 1890 6140
rect 1930 6100 1950 6140
rect 1870 6040 1950 6100
rect 1870 6000 1890 6040
rect 1930 6000 1950 6040
rect 1870 5940 1950 6000
rect 1870 5900 1890 5940
rect 1930 5900 1950 5940
rect 1870 5840 1950 5900
rect 2490 6040 2580 6070
rect 2490 6000 2520 6040
rect 2560 6000 2580 6040
rect 2490 5940 2580 6000
rect 2490 5900 2520 5940
rect 2560 5900 2580 5940
rect 2490 5870 2580 5900
rect 2610 6040 2690 6070
rect 2610 6000 2630 6040
rect 2670 6000 2690 6040
rect 2610 5940 2690 6000
rect 2610 5900 2630 5940
rect 2670 5900 2690 5940
rect 2610 5870 2690 5900
rect 2720 6040 2800 6070
rect 2720 6000 2740 6040
rect 2780 6000 2800 6040
rect 2720 5940 2800 6000
rect 2720 5900 2740 5940
rect 2780 5900 2800 5940
rect 2720 5870 2800 5900
rect 2830 6040 2910 6070
rect 2830 6000 2850 6040
rect 2890 6000 2910 6040
rect 2830 5940 2910 6000
rect 2830 5900 2850 5940
rect 2890 5900 2910 5940
rect 2830 5870 2910 5900
rect 2940 6040 3020 6070
rect 2940 6000 2960 6040
rect 3000 6000 3020 6040
rect 2940 5940 3020 6000
rect 2940 5900 2960 5940
rect 3000 5900 3020 5940
rect 2940 5870 3020 5900
rect 1870 5800 1890 5840
rect 1930 5800 1950 5840
rect 1870 5740 1950 5800
rect 1870 5700 1890 5740
rect 1930 5700 1950 5740
rect 1870 5670 1950 5700
rect 5550 4760 5650 4790
rect 5550 4720 5580 4760
rect 5620 4720 5650 4760
rect -2470 4680 -2390 4710
rect -2470 4640 -2450 4680
rect -2410 4640 -2390 4680
rect -2470 4580 -2390 4640
rect -2470 4540 -2450 4580
rect -2410 4540 -2390 4580
rect -2470 4510 -2390 4540
rect -2350 4680 -2270 4710
rect -2350 4640 -2330 4680
rect -2290 4640 -2270 4680
rect -2350 4580 -2270 4640
rect -2350 4540 -2330 4580
rect -2290 4540 -2270 4580
rect -2350 4510 -2270 4540
rect -2230 4680 -2150 4710
rect -2230 4640 -2210 4680
rect -2170 4640 -2150 4680
rect -2230 4580 -2150 4640
rect -2230 4540 -2210 4580
rect -2170 4540 -2150 4580
rect -2230 4510 -2150 4540
rect -2110 4680 -2030 4710
rect -2110 4640 -2090 4680
rect -2050 4640 -2030 4680
rect -2110 4580 -2030 4640
rect -2110 4540 -2090 4580
rect -2050 4540 -2030 4580
rect -2110 4510 -2030 4540
rect -1990 4680 -1910 4710
rect -1990 4640 -1970 4680
rect -1930 4640 -1910 4680
rect -1990 4580 -1910 4640
rect -1990 4540 -1970 4580
rect -1930 4540 -1910 4580
rect -1990 4510 -1910 4540
rect -1870 4680 -1790 4710
rect -1870 4640 -1850 4680
rect -1810 4640 -1790 4680
rect -1870 4580 -1790 4640
rect -1870 4540 -1850 4580
rect -1810 4540 -1790 4580
rect -1870 4510 -1790 4540
rect -1750 4680 -1670 4710
rect -1750 4640 -1730 4680
rect -1690 4640 -1670 4680
rect -1750 4580 -1670 4640
rect -1750 4540 -1730 4580
rect -1690 4540 -1670 4580
rect -1750 4510 -1670 4540
rect -1630 4680 -1550 4710
rect -1630 4640 -1610 4680
rect -1570 4640 -1550 4680
rect -1630 4580 -1550 4640
rect -1630 4540 -1610 4580
rect -1570 4540 -1550 4580
rect -1630 4510 -1550 4540
rect -1510 4680 -1430 4710
rect -1510 4640 -1490 4680
rect -1450 4640 -1430 4680
rect -1510 4580 -1430 4640
rect -1510 4540 -1490 4580
rect -1450 4540 -1430 4580
rect -1510 4510 -1430 4540
rect -1390 4680 -1310 4710
rect -1390 4640 -1370 4680
rect -1330 4640 -1310 4680
rect -1390 4580 -1310 4640
rect -1390 4540 -1370 4580
rect -1330 4540 -1310 4580
rect -1390 4510 -1310 4540
rect -1270 4680 -1190 4710
rect -1270 4640 -1250 4680
rect -1210 4640 -1190 4680
rect -1270 4580 -1190 4640
rect -1270 4540 -1250 4580
rect -1210 4540 -1190 4580
rect -1270 4510 -1190 4540
rect -1150 4680 -1070 4710
rect -1150 4640 -1130 4680
rect -1090 4640 -1070 4680
rect -1150 4580 -1070 4640
rect -1150 4540 -1130 4580
rect -1090 4540 -1070 4580
rect -1150 4510 -1070 4540
rect -1030 4680 -950 4710
rect -1030 4640 -1010 4680
rect -970 4640 -950 4680
rect -1030 4580 -950 4640
rect -1030 4540 -1010 4580
rect -970 4540 -950 4580
rect -1030 4510 -950 4540
rect -910 4680 -830 4710
rect -910 4640 -890 4680
rect -850 4640 -830 4680
rect -910 4580 -830 4640
rect -910 4540 -890 4580
rect -850 4540 -830 4580
rect -910 4510 -830 4540
rect -790 4680 -710 4710
rect -790 4640 -770 4680
rect -730 4640 -710 4680
rect -790 4580 -710 4640
rect -790 4540 -770 4580
rect -730 4540 -710 4580
rect -790 4510 -710 4540
rect -670 4680 -590 4710
rect -670 4640 -650 4680
rect -610 4640 -590 4680
rect -670 4580 -590 4640
rect -670 4540 -650 4580
rect -610 4540 -590 4580
rect -670 4510 -590 4540
rect -550 4680 -470 4710
rect -550 4640 -530 4680
rect -490 4640 -470 4680
rect -550 4580 -470 4640
rect -550 4540 -530 4580
rect -490 4540 -470 4580
rect -550 4510 -470 4540
rect -430 4680 -350 4710
rect -430 4640 -410 4680
rect -370 4640 -350 4680
rect -430 4580 -350 4640
rect -430 4540 -410 4580
rect -370 4540 -350 4580
rect -430 4510 -350 4540
rect -310 4680 -230 4710
rect -310 4640 -290 4680
rect -250 4640 -230 4680
rect -310 4580 -230 4640
rect -310 4540 -290 4580
rect -250 4540 -230 4580
rect -310 4510 -230 4540
rect -190 4680 -110 4710
rect -190 4640 -170 4680
rect -130 4640 -110 4680
rect -190 4580 -110 4640
rect -190 4540 -170 4580
rect -130 4540 -110 4580
rect -190 4510 -110 4540
rect -70 4680 10 4710
rect -70 4640 -50 4680
rect -10 4640 10 4680
rect -70 4580 10 4640
rect -70 4540 -50 4580
rect -10 4540 10 4580
rect -70 4510 10 4540
rect 570 4680 650 4710
rect 570 4640 590 4680
rect 630 4640 650 4680
rect 570 4580 650 4640
rect 570 4540 590 4580
rect 630 4540 650 4580
rect 570 4510 650 4540
rect 690 4680 770 4710
rect 690 4640 710 4680
rect 750 4640 770 4680
rect 690 4580 770 4640
rect 690 4540 710 4580
rect 750 4540 770 4580
rect 690 4510 770 4540
rect 810 4680 890 4710
rect 810 4640 830 4680
rect 870 4640 890 4680
rect 810 4580 890 4640
rect 810 4540 830 4580
rect 870 4540 890 4580
rect 810 4510 890 4540
rect 930 4680 1010 4710
rect 930 4640 950 4680
rect 990 4640 1010 4680
rect 930 4580 1010 4640
rect 930 4540 950 4580
rect 990 4540 1010 4580
rect 930 4510 1010 4540
rect 1050 4680 1130 4710
rect 1050 4640 1070 4680
rect 1110 4640 1130 4680
rect 1050 4580 1130 4640
rect 1050 4540 1070 4580
rect 1110 4540 1130 4580
rect 1050 4510 1130 4540
rect 1170 4680 1250 4710
rect 1170 4640 1190 4680
rect 1230 4640 1250 4680
rect 1170 4580 1250 4640
rect 1170 4540 1190 4580
rect 1230 4540 1250 4580
rect 1170 4510 1250 4540
rect 1290 4680 1370 4710
rect 1290 4640 1310 4680
rect 1350 4640 1370 4680
rect 1290 4580 1370 4640
rect 1290 4540 1310 4580
rect 1350 4540 1370 4580
rect 1290 4510 1370 4540
rect 1410 4680 1490 4710
rect 1410 4640 1430 4680
rect 1470 4640 1490 4680
rect 1410 4580 1490 4640
rect 1410 4540 1430 4580
rect 1470 4540 1490 4580
rect 1410 4510 1490 4540
rect 1530 4680 1610 4710
rect 1530 4640 1550 4680
rect 1590 4640 1610 4680
rect 1530 4580 1610 4640
rect 1530 4540 1550 4580
rect 1590 4540 1610 4580
rect 1530 4510 1610 4540
rect 1650 4680 1730 4710
rect 1650 4640 1670 4680
rect 1710 4640 1730 4680
rect 1650 4580 1730 4640
rect 1650 4540 1670 4580
rect 1710 4540 1730 4580
rect 1650 4510 1730 4540
rect 1770 4680 1850 4710
rect 1770 4640 1790 4680
rect 1830 4640 1850 4680
rect 1770 4580 1850 4640
rect 1770 4540 1790 4580
rect 1830 4540 1850 4580
rect 1770 4510 1850 4540
rect 1890 4680 1970 4710
rect 1890 4640 1910 4680
rect 1950 4640 1970 4680
rect 1890 4580 1970 4640
rect 1890 4540 1910 4580
rect 1950 4540 1970 4580
rect 1890 4510 1970 4540
rect 2010 4680 2090 4710
rect 2010 4640 2030 4680
rect 2070 4640 2090 4680
rect 2010 4580 2090 4640
rect 2010 4540 2030 4580
rect 2070 4540 2090 4580
rect 2010 4510 2090 4540
rect 2130 4680 2210 4710
rect 2130 4640 2150 4680
rect 2190 4640 2210 4680
rect 2130 4580 2210 4640
rect 2130 4540 2150 4580
rect 2190 4540 2210 4580
rect 2130 4510 2210 4540
rect 2250 4680 2330 4710
rect 2250 4640 2270 4680
rect 2310 4640 2330 4680
rect 2250 4580 2330 4640
rect 2250 4540 2270 4580
rect 2310 4540 2330 4580
rect 2250 4510 2330 4540
rect 2370 4680 2450 4710
rect 2370 4640 2390 4680
rect 2430 4640 2450 4680
rect 2370 4580 2450 4640
rect 2370 4540 2390 4580
rect 2430 4540 2450 4580
rect 2370 4510 2450 4540
rect 2490 4680 2570 4710
rect 2490 4640 2510 4680
rect 2550 4640 2570 4680
rect 2490 4580 2570 4640
rect 2490 4540 2510 4580
rect 2550 4540 2570 4580
rect 2490 4510 2570 4540
rect 2610 4680 2690 4710
rect 2610 4640 2630 4680
rect 2670 4640 2690 4680
rect 2610 4580 2690 4640
rect 2610 4540 2630 4580
rect 2670 4540 2690 4580
rect 2610 4510 2690 4540
rect 2730 4680 2810 4710
rect 2730 4640 2750 4680
rect 2790 4640 2810 4680
rect 2730 4580 2810 4640
rect 2730 4540 2750 4580
rect 2790 4540 2810 4580
rect 2730 4510 2810 4540
rect 2850 4680 2930 4710
rect 2850 4640 2870 4680
rect 2910 4640 2930 4680
rect 2850 4580 2930 4640
rect 2850 4540 2870 4580
rect 2910 4540 2930 4580
rect 2850 4510 2930 4540
rect 2970 4680 3050 4710
rect 2970 4640 2990 4680
rect 3030 4640 3050 4680
rect 2970 4580 3050 4640
rect 5550 4660 5650 4720
rect 5550 4620 5580 4660
rect 5620 4620 5650 4660
rect 5550 4590 5650 4620
rect 5680 4760 5780 4790
rect 5680 4720 5710 4760
rect 5750 4720 5780 4760
rect 5680 4660 5780 4720
rect 5680 4620 5710 4660
rect 5750 4620 5780 4660
rect 5680 4590 5780 4620
rect 5810 4760 5910 4790
rect 5810 4720 5840 4760
rect 5880 4720 5910 4760
rect 5810 4660 5910 4720
rect 5810 4620 5840 4660
rect 5880 4620 5910 4660
rect 5810 4590 5910 4620
rect 5940 4760 6040 4790
rect 5940 4720 5970 4760
rect 6010 4720 6040 4760
rect 5940 4660 6040 4720
rect 5940 4620 5970 4660
rect 6010 4620 6040 4660
rect 5940 4590 6040 4620
rect 6070 4760 6170 4790
rect 6070 4720 6100 4760
rect 6140 4720 6170 4760
rect 6070 4660 6170 4720
rect 6070 4620 6100 4660
rect 6140 4620 6170 4660
rect 6070 4590 6170 4620
rect 6200 4760 6300 4790
rect 6200 4720 6230 4760
rect 6270 4720 6300 4760
rect 6200 4660 6300 4720
rect 6200 4620 6230 4660
rect 6270 4620 6300 4660
rect 6200 4590 6300 4620
rect 6330 4760 6430 4790
rect 6330 4720 6360 4760
rect 6400 4720 6430 4760
rect 6330 4660 6430 4720
rect 6330 4620 6360 4660
rect 6400 4620 6430 4660
rect 6330 4590 6430 4620
rect 6690 4760 6790 4790
rect 6690 4720 6720 4760
rect 6760 4720 6790 4760
rect 6690 4660 6790 4720
rect 6690 4620 6720 4660
rect 6760 4620 6790 4660
rect 6690 4590 6790 4620
rect 6820 4760 6920 4790
rect 6820 4720 6850 4760
rect 6890 4720 6920 4760
rect 6820 4660 6920 4720
rect 6820 4620 6850 4660
rect 6890 4620 6920 4660
rect 6820 4590 6920 4620
rect 6950 4760 7050 4790
rect 6950 4720 6980 4760
rect 7020 4720 7050 4760
rect 6950 4660 7050 4720
rect 6950 4620 6980 4660
rect 7020 4620 7050 4660
rect 6950 4590 7050 4620
rect 7080 4760 7180 4790
rect 7080 4720 7110 4760
rect 7150 4720 7180 4760
rect 7080 4660 7180 4720
rect 7080 4620 7110 4660
rect 7150 4620 7180 4660
rect 7080 4590 7180 4620
rect 7210 4760 7310 4790
rect 7210 4720 7240 4760
rect 7280 4720 7310 4760
rect 7210 4660 7310 4720
rect 7210 4620 7240 4660
rect 7280 4620 7310 4660
rect 7210 4590 7310 4620
rect 7340 4760 7440 4790
rect 7340 4720 7370 4760
rect 7410 4720 7440 4760
rect 7340 4660 7440 4720
rect 7340 4620 7370 4660
rect 7410 4620 7440 4660
rect 7340 4590 7440 4620
rect 7470 4760 7570 4790
rect 7470 4720 7500 4760
rect 7540 4720 7570 4760
rect 7470 4660 7570 4720
rect 7470 4620 7500 4660
rect 7540 4620 7570 4660
rect 7470 4590 7570 4620
rect 7830 4760 7930 4790
rect 7830 4720 7860 4760
rect 7900 4720 7930 4760
rect 7830 4660 7930 4720
rect 7830 4620 7860 4660
rect 7900 4620 7930 4660
rect 7830 4590 7930 4620
rect 7960 4760 8060 4790
rect 7960 4720 7990 4760
rect 8030 4720 8060 4760
rect 7960 4660 8060 4720
rect 7960 4620 7990 4660
rect 8030 4620 8060 4660
rect 7960 4590 8060 4620
rect 8090 4760 8190 4790
rect 8090 4720 8120 4760
rect 8160 4720 8190 4760
rect 8090 4660 8190 4720
rect 8090 4620 8120 4660
rect 8160 4620 8190 4660
rect 8090 4590 8190 4620
rect 8220 4760 8320 4790
rect 8220 4720 8250 4760
rect 8290 4720 8320 4760
rect 8220 4660 8320 4720
rect 8220 4620 8250 4660
rect 8290 4620 8320 4660
rect 8220 4590 8320 4620
rect 8350 4760 8450 4790
rect 8350 4720 8380 4760
rect 8420 4720 8450 4760
rect 8350 4660 8450 4720
rect 8350 4620 8380 4660
rect 8420 4620 8450 4660
rect 8350 4590 8450 4620
rect 8480 4760 8580 4790
rect 8480 4720 8510 4760
rect 8550 4720 8580 4760
rect 8480 4660 8580 4720
rect 8480 4620 8510 4660
rect 8550 4620 8580 4660
rect 8480 4590 8580 4620
rect 8610 4760 8710 4790
rect 8610 4720 8640 4760
rect 8680 4720 8710 4760
rect 8610 4660 8710 4720
rect 8610 4620 8640 4660
rect 8680 4620 8710 4660
rect 8610 4590 8710 4620
rect 2970 4540 2990 4580
rect 3030 4540 3050 4580
rect 2970 4510 3050 4540
rect 5620 4110 5720 4140
rect 5620 4070 5650 4110
rect 5690 4070 5720 4110
rect 5620 4010 5720 4070
rect 5620 3970 5650 4010
rect 5690 3970 5720 4010
rect 5620 3910 5720 3970
rect 5620 3870 5650 3910
rect 5690 3870 5720 3910
rect 5620 3810 5720 3870
rect 5620 3770 5650 3810
rect 5690 3770 5720 3810
rect 5620 3710 5720 3770
rect 5620 3670 5650 3710
rect 5690 3670 5720 3710
rect 5620 3640 5720 3670
rect 5820 4110 5920 4140
rect 5820 4070 5850 4110
rect 5890 4070 5920 4110
rect 5820 4010 5920 4070
rect 5820 3970 5850 4010
rect 5890 3970 5920 4010
rect 5820 3910 5920 3970
rect 5820 3870 5850 3910
rect 5890 3870 5920 3910
rect 5820 3810 5920 3870
rect 5820 3770 5850 3810
rect 5890 3770 5920 3810
rect 5820 3710 5920 3770
rect 5820 3670 5850 3710
rect 5890 3670 5920 3710
rect 5820 3640 5920 3670
rect 6020 4110 6120 4140
rect 6020 4070 6050 4110
rect 6090 4070 6120 4110
rect 6020 4010 6120 4070
rect 6020 3970 6050 4010
rect 6090 3970 6120 4010
rect 6020 3910 6120 3970
rect 6020 3870 6050 3910
rect 6090 3870 6120 3910
rect 6020 3810 6120 3870
rect 6020 3770 6050 3810
rect 6090 3770 6120 3810
rect 6020 3710 6120 3770
rect 6020 3670 6050 3710
rect 6090 3670 6120 3710
rect 6020 3640 6120 3670
rect 6220 4110 6320 4140
rect 6220 4070 6250 4110
rect 6290 4070 6320 4110
rect 6220 4010 6320 4070
rect 6220 3970 6250 4010
rect 6290 3970 6320 4010
rect 6220 3910 6320 3970
rect 6220 3870 6250 3910
rect 6290 3870 6320 3910
rect 6220 3810 6320 3870
rect 6220 3770 6250 3810
rect 6290 3770 6320 3810
rect 6220 3710 6320 3770
rect 6220 3670 6250 3710
rect 6290 3670 6320 3710
rect 6220 3640 6320 3670
rect 6420 4110 6520 4140
rect 6420 4070 6450 4110
rect 6490 4070 6520 4110
rect 6420 4010 6520 4070
rect 6420 3970 6450 4010
rect 6490 3970 6520 4010
rect 6420 3910 6520 3970
rect 6420 3870 6450 3910
rect 6490 3870 6520 3910
rect 6420 3810 6520 3870
rect 6420 3770 6450 3810
rect 6490 3770 6520 3810
rect 6420 3710 6520 3770
rect 6420 3670 6450 3710
rect 6490 3670 6520 3710
rect 6420 3640 6520 3670
rect 6620 4110 6720 4140
rect 6620 4070 6650 4110
rect 6690 4070 6720 4110
rect 6620 4010 6720 4070
rect 6620 3970 6650 4010
rect 6690 3970 6720 4010
rect 6620 3910 6720 3970
rect 6620 3870 6650 3910
rect 6690 3870 6720 3910
rect 6620 3810 6720 3870
rect 6620 3770 6650 3810
rect 6690 3770 6720 3810
rect 6620 3710 6720 3770
rect 6620 3670 6650 3710
rect 6690 3670 6720 3710
rect 6620 3640 6720 3670
rect 6820 4110 6920 4140
rect 6820 4070 6850 4110
rect 6890 4070 6920 4110
rect 6820 4010 6920 4070
rect 6820 3970 6850 4010
rect 6890 3970 6920 4010
rect 6820 3910 6920 3970
rect 6820 3870 6850 3910
rect 6890 3870 6920 3910
rect 6820 3810 6920 3870
rect 6820 3770 6850 3810
rect 6890 3770 6920 3810
rect 6820 3710 6920 3770
rect 6820 3670 6850 3710
rect 6890 3670 6920 3710
rect 6820 3640 6920 3670
rect 7020 4110 7120 4140
rect 7020 4070 7050 4110
rect 7090 4070 7120 4110
rect 7020 4010 7120 4070
rect 7020 3970 7050 4010
rect 7090 3970 7120 4010
rect 7020 3910 7120 3970
rect 7020 3870 7050 3910
rect 7090 3870 7120 3910
rect 7020 3810 7120 3870
rect 7020 3770 7050 3810
rect 7090 3770 7120 3810
rect 7020 3710 7120 3770
rect 7020 3670 7050 3710
rect 7090 3670 7120 3710
rect 7020 3640 7120 3670
rect 7220 4110 7320 4140
rect 7220 4070 7250 4110
rect 7290 4070 7320 4110
rect 7220 4010 7320 4070
rect 7220 3970 7250 4010
rect 7290 3970 7320 4010
rect 7220 3910 7320 3970
rect 7220 3870 7250 3910
rect 7290 3870 7320 3910
rect 7220 3810 7320 3870
rect 7220 3770 7250 3810
rect 7290 3770 7320 3810
rect 7220 3710 7320 3770
rect 7220 3670 7250 3710
rect 7290 3670 7320 3710
rect 7220 3640 7320 3670
rect 7420 4110 7520 4140
rect 7420 4070 7450 4110
rect 7490 4070 7520 4110
rect 7420 4010 7520 4070
rect 7420 3970 7450 4010
rect 7490 3970 7520 4010
rect 7420 3910 7520 3970
rect 7420 3870 7450 3910
rect 7490 3870 7520 3910
rect 7420 3810 7520 3870
rect 7420 3770 7450 3810
rect 7490 3770 7520 3810
rect 7420 3710 7520 3770
rect 7420 3670 7450 3710
rect 7490 3670 7520 3710
rect 7420 3640 7520 3670
rect 7620 4110 7720 4140
rect 7620 4070 7650 4110
rect 7690 4070 7720 4110
rect 7620 4010 7720 4070
rect 7620 3970 7650 4010
rect 7690 3970 7720 4010
rect 7620 3910 7720 3970
rect 7620 3870 7650 3910
rect 7690 3870 7720 3910
rect 7620 3810 7720 3870
rect 7620 3770 7650 3810
rect 7690 3770 7720 3810
rect 7620 3710 7720 3770
rect 7620 3670 7650 3710
rect 7690 3670 7720 3710
rect 7620 3640 7720 3670
rect -1410 1198 -730 1250
rect -1410 1164 -1358 1198
rect -1324 1164 -1268 1198
rect -1234 1164 -1178 1198
rect -1144 1164 -1088 1198
rect -1054 1164 -998 1198
rect -964 1164 -908 1198
rect -874 1164 -818 1198
rect -784 1164 -730 1198
rect -1410 1108 -730 1164
rect -1410 1074 -1358 1108
rect -1324 1074 -1268 1108
rect -1234 1074 -1178 1108
rect -1144 1074 -1088 1108
rect -1054 1074 -998 1108
rect -964 1074 -908 1108
rect -874 1074 -818 1108
rect -784 1074 -730 1108
rect -1410 1018 -730 1074
rect -1410 984 -1358 1018
rect -1324 984 -1268 1018
rect -1234 984 -1178 1018
rect -1144 984 -1088 1018
rect -1054 984 -998 1018
rect -964 984 -908 1018
rect -874 984 -818 1018
rect -784 984 -730 1018
rect -1410 928 -730 984
rect -1410 894 -1358 928
rect -1324 894 -1268 928
rect -1234 894 -1178 928
rect -1144 894 -1088 928
rect -1054 894 -998 928
rect -964 894 -908 928
rect -874 894 -818 928
rect -784 894 -730 928
rect -1410 838 -730 894
rect -1410 804 -1358 838
rect -1324 804 -1268 838
rect -1234 804 -1178 838
rect -1144 804 -1088 838
rect -1054 804 -998 838
rect -964 804 -908 838
rect -874 804 -818 838
rect -784 804 -730 838
rect -1410 748 -730 804
rect -1410 714 -1358 748
rect -1324 714 -1268 748
rect -1234 714 -1178 748
rect -1144 714 -1088 748
rect -1054 714 -998 748
rect -964 714 -908 748
rect -874 714 -818 748
rect -784 714 -730 748
rect -1410 658 -730 714
rect -1410 624 -1358 658
rect -1324 624 -1268 658
rect -1234 624 -1178 658
rect -1144 624 -1088 658
rect -1054 624 -998 658
rect -964 624 -908 658
rect -874 624 -818 658
rect -784 624 -730 658
rect -1410 570 -730 624
rect -50 1198 630 1250
rect -50 1164 2 1198
rect 36 1164 92 1198
rect 126 1164 182 1198
rect 216 1164 272 1198
rect 306 1164 362 1198
rect 396 1164 452 1198
rect 486 1164 542 1198
rect 576 1164 630 1198
rect -50 1108 630 1164
rect -50 1074 2 1108
rect 36 1074 92 1108
rect 126 1074 182 1108
rect 216 1074 272 1108
rect 306 1074 362 1108
rect 396 1074 452 1108
rect 486 1074 542 1108
rect 576 1074 630 1108
rect -50 1018 630 1074
rect -50 984 2 1018
rect 36 984 92 1018
rect 126 984 182 1018
rect 216 984 272 1018
rect 306 984 362 1018
rect 396 984 452 1018
rect 486 984 542 1018
rect 576 984 630 1018
rect -50 928 630 984
rect -50 894 2 928
rect 36 894 92 928
rect 126 894 182 928
rect 216 894 272 928
rect 306 894 362 928
rect 396 894 452 928
rect 486 894 542 928
rect 576 894 630 928
rect -50 838 630 894
rect -50 804 2 838
rect 36 804 92 838
rect 126 804 182 838
rect 216 804 272 838
rect 306 804 362 838
rect 396 804 452 838
rect 486 804 542 838
rect 576 804 630 838
rect -50 748 630 804
rect -50 714 2 748
rect 36 714 92 748
rect 126 714 182 748
rect 216 714 272 748
rect 306 714 362 748
rect 396 714 452 748
rect 486 714 542 748
rect 576 714 630 748
rect -50 658 630 714
rect -50 624 2 658
rect 36 624 92 658
rect 126 624 182 658
rect 216 624 272 658
rect 306 624 362 658
rect 396 624 452 658
rect 486 624 542 658
rect 576 624 630 658
rect -50 570 630 624
rect 1310 1198 1990 1250
rect 1310 1164 1362 1198
rect 1396 1164 1452 1198
rect 1486 1164 1542 1198
rect 1576 1164 1632 1198
rect 1666 1164 1722 1198
rect 1756 1164 1812 1198
rect 1846 1164 1902 1198
rect 1936 1164 1990 1198
rect 1310 1108 1990 1164
rect 1310 1074 1362 1108
rect 1396 1074 1452 1108
rect 1486 1074 1542 1108
rect 1576 1074 1632 1108
rect 1666 1074 1722 1108
rect 1756 1074 1812 1108
rect 1846 1074 1902 1108
rect 1936 1074 1990 1108
rect 1310 1018 1990 1074
rect 1310 984 1362 1018
rect 1396 984 1452 1018
rect 1486 984 1542 1018
rect 1576 984 1632 1018
rect 1666 984 1722 1018
rect 1756 984 1812 1018
rect 1846 984 1902 1018
rect 1936 984 1990 1018
rect 1310 928 1990 984
rect 1310 894 1362 928
rect 1396 894 1452 928
rect 1486 894 1542 928
rect 1576 894 1632 928
rect 1666 894 1722 928
rect 1756 894 1812 928
rect 1846 894 1902 928
rect 1936 894 1990 928
rect 1310 838 1990 894
rect 1310 804 1362 838
rect 1396 804 1452 838
rect 1486 804 1542 838
rect 1576 804 1632 838
rect 1666 804 1722 838
rect 1756 804 1812 838
rect 1846 804 1902 838
rect 1936 804 1990 838
rect 1310 748 1990 804
rect 1310 714 1362 748
rect 1396 714 1452 748
rect 1486 714 1542 748
rect 1576 714 1632 748
rect 1666 714 1722 748
rect 1756 714 1812 748
rect 1846 714 1902 748
rect 1936 714 1990 748
rect 1310 658 1990 714
rect 1310 624 1362 658
rect 1396 624 1452 658
rect 1486 624 1542 658
rect 1576 624 1632 658
rect 1666 624 1722 658
rect 1756 624 1812 658
rect 1846 624 1902 658
rect 1936 624 1990 658
rect 1310 570 1990 624
rect -1410 -162 -730 -110
rect -1410 -196 -1358 -162
rect -1324 -196 -1268 -162
rect -1234 -196 -1178 -162
rect -1144 -196 -1088 -162
rect -1054 -196 -998 -162
rect -964 -196 -908 -162
rect -874 -196 -818 -162
rect -784 -196 -730 -162
rect -1410 -252 -730 -196
rect -1410 -286 -1358 -252
rect -1324 -286 -1268 -252
rect -1234 -286 -1178 -252
rect -1144 -286 -1088 -252
rect -1054 -286 -998 -252
rect -964 -286 -908 -252
rect -874 -286 -818 -252
rect -784 -286 -730 -252
rect -1410 -342 -730 -286
rect -1410 -376 -1358 -342
rect -1324 -376 -1268 -342
rect -1234 -376 -1178 -342
rect -1144 -376 -1088 -342
rect -1054 -376 -998 -342
rect -964 -376 -908 -342
rect -874 -376 -818 -342
rect -784 -376 -730 -342
rect -1410 -432 -730 -376
rect -1410 -466 -1358 -432
rect -1324 -466 -1268 -432
rect -1234 -466 -1178 -432
rect -1144 -466 -1088 -432
rect -1054 -466 -998 -432
rect -964 -466 -908 -432
rect -874 -466 -818 -432
rect -784 -466 -730 -432
rect -1410 -522 -730 -466
rect -1410 -556 -1358 -522
rect -1324 -556 -1268 -522
rect -1234 -556 -1178 -522
rect -1144 -556 -1088 -522
rect -1054 -556 -998 -522
rect -964 -556 -908 -522
rect -874 -556 -818 -522
rect -784 -556 -730 -522
rect -1410 -612 -730 -556
rect -1410 -646 -1358 -612
rect -1324 -646 -1268 -612
rect -1234 -646 -1178 -612
rect -1144 -646 -1088 -612
rect -1054 -646 -998 -612
rect -964 -646 -908 -612
rect -874 -646 -818 -612
rect -784 -646 -730 -612
rect -1410 -702 -730 -646
rect -1410 -736 -1358 -702
rect -1324 -736 -1268 -702
rect -1234 -736 -1178 -702
rect -1144 -736 -1088 -702
rect -1054 -736 -998 -702
rect -964 -736 -908 -702
rect -874 -736 -818 -702
rect -784 -736 -730 -702
rect -1410 -790 -730 -736
rect -50 -162 630 -110
rect -50 -196 2 -162
rect 36 -196 92 -162
rect 126 -196 182 -162
rect 216 -196 272 -162
rect 306 -196 362 -162
rect 396 -196 452 -162
rect 486 -196 542 -162
rect 576 -196 630 -162
rect -50 -252 630 -196
rect -50 -286 2 -252
rect 36 -286 92 -252
rect 126 -286 182 -252
rect 216 -286 272 -252
rect 306 -286 362 -252
rect 396 -286 452 -252
rect 486 -286 542 -252
rect 576 -286 630 -252
rect -50 -342 630 -286
rect -50 -376 2 -342
rect 36 -376 92 -342
rect 126 -376 182 -342
rect 216 -376 272 -342
rect 306 -376 362 -342
rect 396 -376 452 -342
rect 486 -376 542 -342
rect 576 -376 630 -342
rect -50 -432 630 -376
rect -50 -466 2 -432
rect 36 -466 92 -432
rect 126 -466 182 -432
rect 216 -466 272 -432
rect 306 -466 362 -432
rect 396 -466 452 -432
rect 486 -466 542 -432
rect 576 -466 630 -432
rect -50 -522 630 -466
rect -50 -556 2 -522
rect 36 -556 92 -522
rect 126 -556 182 -522
rect 216 -556 272 -522
rect 306 -556 362 -522
rect 396 -556 452 -522
rect 486 -556 542 -522
rect 576 -556 630 -522
rect -50 -612 630 -556
rect -50 -646 2 -612
rect 36 -646 92 -612
rect 126 -646 182 -612
rect 216 -646 272 -612
rect 306 -646 362 -612
rect 396 -646 452 -612
rect 486 -646 542 -612
rect 576 -646 630 -612
rect -50 -702 630 -646
rect -50 -736 2 -702
rect 36 -736 92 -702
rect 126 -736 182 -702
rect 216 -736 272 -702
rect 306 -736 362 -702
rect 396 -736 452 -702
rect 486 -736 542 -702
rect 576 -736 630 -702
rect -50 -790 630 -736
rect 1310 -162 1990 -110
rect 1310 -196 1362 -162
rect 1396 -196 1452 -162
rect 1486 -196 1542 -162
rect 1576 -196 1632 -162
rect 1666 -196 1722 -162
rect 1756 -196 1812 -162
rect 1846 -196 1902 -162
rect 1936 -196 1990 -162
rect 1310 -252 1990 -196
rect 1310 -286 1362 -252
rect 1396 -286 1452 -252
rect 1486 -286 1542 -252
rect 1576 -286 1632 -252
rect 1666 -286 1722 -252
rect 1756 -286 1812 -252
rect 1846 -286 1902 -252
rect 1936 -286 1990 -252
rect 1310 -342 1990 -286
rect 1310 -376 1362 -342
rect 1396 -376 1452 -342
rect 1486 -376 1542 -342
rect 1576 -376 1632 -342
rect 1666 -376 1722 -342
rect 1756 -376 1812 -342
rect 1846 -376 1902 -342
rect 1936 -376 1990 -342
rect 1310 -432 1990 -376
rect 1310 -466 1362 -432
rect 1396 -466 1452 -432
rect 1486 -466 1542 -432
rect 1576 -466 1632 -432
rect 1666 -466 1722 -432
rect 1756 -466 1812 -432
rect 1846 -466 1902 -432
rect 1936 -466 1990 -432
rect 1310 -522 1990 -466
rect 1310 -556 1362 -522
rect 1396 -556 1452 -522
rect 1486 -556 1542 -522
rect 1576 -556 1632 -522
rect 1666 -556 1722 -522
rect 1756 -556 1812 -522
rect 1846 -556 1902 -522
rect 1936 -556 1990 -522
rect 1310 -612 1990 -556
rect 1310 -646 1362 -612
rect 1396 -646 1452 -612
rect 1486 -646 1542 -612
rect 1576 -646 1632 -612
rect 1666 -646 1722 -612
rect 1756 -646 1812 -612
rect 1846 -646 1902 -612
rect 1936 -646 1990 -612
rect 1310 -702 1990 -646
rect 1310 -736 1362 -702
rect 1396 -736 1452 -702
rect 1486 -736 1542 -702
rect 1576 -736 1632 -702
rect 1666 -736 1722 -702
rect 1756 -736 1812 -702
rect 1846 -736 1902 -702
rect 1936 -736 1990 -702
rect 1310 -790 1990 -736
rect -1410 -1522 -730 -1470
rect -1410 -1556 -1358 -1522
rect -1324 -1556 -1268 -1522
rect -1234 -1556 -1178 -1522
rect -1144 -1556 -1088 -1522
rect -1054 -1556 -998 -1522
rect -964 -1556 -908 -1522
rect -874 -1556 -818 -1522
rect -784 -1556 -730 -1522
rect -1410 -1612 -730 -1556
rect -1410 -1646 -1358 -1612
rect -1324 -1646 -1268 -1612
rect -1234 -1646 -1178 -1612
rect -1144 -1646 -1088 -1612
rect -1054 -1646 -998 -1612
rect -964 -1646 -908 -1612
rect -874 -1646 -818 -1612
rect -784 -1646 -730 -1612
rect -1410 -1702 -730 -1646
rect -1410 -1736 -1358 -1702
rect -1324 -1736 -1268 -1702
rect -1234 -1736 -1178 -1702
rect -1144 -1736 -1088 -1702
rect -1054 -1736 -998 -1702
rect -964 -1736 -908 -1702
rect -874 -1736 -818 -1702
rect -784 -1736 -730 -1702
rect -1410 -1792 -730 -1736
rect -1410 -1826 -1358 -1792
rect -1324 -1826 -1268 -1792
rect -1234 -1826 -1178 -1792
rect -1144 -1826 -1088 -1792
rect -1054 -1826 -998 -1792
rect -964 -1826 -908 -1792
rect -874 -1826 -818 -1792
rect -784 -1826 -730 -1792
rect -1410 -1882 -730 -1826
rect -1410 -1916 -1358 -1882
rect -1324 -1916 -1268 -1882
rect -1234 -1916 -1178 -1882
rect -1144 -1916 -1088 -1882
rect -1054 -1916 -998 -1882
rect -964 -1916 -908 -1882
rect -874 -1916 -818 -1882
rect -784 -1916 -730 -1882
rect -1410 -1972 -730 -1916
rect -1410 -2006 -1358 -1972
rect -1324 -2006 -1268 -1972
rect -1234 -2006 -1178 -1972
rect -1144 -2006 -1088 -1972
rect -1054 -2006 -998 -1972
rect -964 -2006 -908 -1972
rect -874 -2006 -818 -1972
rect -784 -2006 -730 -1972
rect -1410 -2062 -730 -2006
rect -1410 -2096 -1358 -2062
rect -1324 -2096 -1268 -2062
rect -1234 -2096 -1178 -2062
rect -1144 -2096 -1088 -2062
rect -1054 -2096 -998 -2062
rect -964 -2096 -908 -2062
rect -874 -2096 -818 -2062
rect -784 -2096 -730 -2062
rect -1410 -2150 -730 -2096
rect -50 -1522 630 -1470
rect -50 -1556 2 -1522
rect 36 -1556 92 -1522
rect 126 -1556 182 -1522
rect 216 -1556 272 -1522
rect 306 -1556 362 -1522
rect 396 -1556 452 -1522
rect 486 -1556 542 -1522
rect 576 -1556 630 -1522
rect -50 -1612 630 -1556
rect -50 -1646 2 -1612
rect 36 -1646 92 -1612
rect 126 -1646 182 -1612
rect 216 -1646 272 -1612
rect 306 -1646 362 -1612
rect 396 -1646 452 -1612
rect 486 -1646 542 -1612
rect 576 -1646 630 -1612
rect -50 -1702 630 -1646
rect -50 -1736 2 -1702
rect 36 -1736 92 -1702
rect 126 -1736 182 -1702
rect 216 -1736 272 -1702
rect 306 -1736 362 -1702
rect 396 -1736 452 -1702
rect 486 -1736 542 -1702
rect 576 -1736 630 -1702
rect -50 -1792 630 -1736
rect -50 -1826 2 -1792
rect 36 -1826 92 -1792
rect 126 -1826 182 -1792
rect 216 -1826 272 -1792
rect 306 -1826 362 -1792
rect 396 -1826 452 -1792
rect 486 -1826 542 -1792
rect 576 -1826 630 -1792
rect -50 -1882 630 -1826
rect -50 -1916 2 -1882
rect 36 -1916 92 -1882
rect 126 -1916 182 -1882
rect 216 -1916 272 -1882
rect 306 -1916 362 -1882
rect 396 -1916 452 -1882
rect 486 -1916 542 -1882
rect 576 -1916 630 -1882
rect -50 -1972 630 -1916
rect -50 -2006 2 -1972
rect 36 -2006 92 -1972
rect 126 -2006 182 -1972
rect 216 -2006 272 -1972
rect 306 -2006 362 -1972
rect 396 -2006 452 -1972
rect 486 -2006 542 -1972
rect 576 -2006 630 -1972
rect -50 -2062 630 -2006
rect -50 -2096 2 -2062
rect 36 -2096 92 -2062
rect 126 -2096 182 -2062
rect 216 -2096 272 -2062
rect 306 -2096 362 -2062
rect 396 -2096 452 -2062
rect 486 -2096 542 -2062
rect 576 -2096 630 -2062
rect -50 -2150 630 -2096
rect 1310 -1522 1990 -1470
rect 1310 -1556 1362 -1522
rect 1396 -1556 1452 -1522
rect 1486 -1556 1542 -1522
rect 1576 -1556 1632 -1522
rect 1666 -1556 1722 -1522
rect 1756 -1556 1812 -1522
rect 1846 -1556 1902 -1522
rect 1936 -1556 1990 -1522
rect 1310 -1612 1990 -1556
rect 1310 -1646 1362 -1612
rect 1396 -1646 1452 -1612
rect 1486 -1646 1542 -1612
rect 1576 -1646 1632 -1612
rect 1666 -1646 1722 -1612
rect 1756 -1646 1812 -1612
rect 1846 -1646 1902 -1612
rect 1936 -1646 1990 -1612
rect 1310 -1702 1990 -1646
rect 1310 -1736 1362 -1702
rect 1396 -1736 1452 -1702
rect 1486 -1736 1542 -1702
rect 1576 -1736 1632 -1702
rect 1666 -1736 1722 -1702
rect 1756 -1736 1812 -1702
rect 1846 -1736 1902 -1702
rect 1936 -1736 1990 -1702
rect 1310 -1792 1990 -1736
rect 1310 -1826 1362 -1792
rect 1396 -1826 1452 -1792
rect 1486 -1826 1542 -1792
rect 1576 -1826 1632 -1792
rect 1666 -1826 1722 -1792
rect 1756 -1826 1812 -1792
rect 1846 -1826 1902 -1792
rect 1936 -1826 1990 -1792
rect 1310 -1882 1990 -1826
rect 1310 -1916 1362 -1882
rect 1396 -1916 1452 -1882
rect 1486 -1916 1542 -1882
rect 1576 -1916 1632 -1882
rect 1666 -1916 1722 -1882
rect 1756 -1916 1812 -1882
rect 1846 -1916 1902 -1882
rect 1936 -1916 1990 -1882
rect 1310 -1972 1990 -1916
rect 1310 -2006 1362 -1972
rect 1396 -2006 1452 -1972
rect 1486 -2006 1542 -1972
rect 1576 -2006 1632 -1972
rect 1666 -2006 1722 -1972
rect 1756 -2006 1812 -1972
rect 1846 -2006 1902 -1972
rect 1936 -2006 1990 -1972
rect 1310 -2062 1990 -2006
rect 1310 -2096 1362 -2062
rect 1396 -2096 1452 -2062
rect 1486 -2096 1542 -2062
rect 1576 -2096 1632 -2062
rect 1666 -2096 1722 -2062
rect 1756 -2096 1812 -2062
rect 1846 -2096 1902 -2062
rect 1936 -2096 1990 -2062
rect 1310 -2150 1990 -2096
<< ndiffc >>
rect 9320 13720 9360 13760
rect 9320 13620 9360 13660
rect 9430 13720 9470 13760
rect 9430 13620 9470 13660
rect 9840 13720 9880 13760
rect 9840 13620 9880 13660
rect 9950 13720 9990 13760
rect 9950 13620 9990 13660
rect 10360 13720 10400 13760
rect 10360 13620 10400 13660
rect 10470 13720 10510 13760
rect 10470 13620 10510 13660
rect 10960 13720 11000 13760
rect 10960 13620 11000 13660
rect 11070 13720 11110 13760
rect 11070 13620 11110 13660
rect 9320 13340 9360 13380
rect 9320 13240 9360 13280
rect 9430 13340 9470 13380
rect 9430 13240 9470 13280
rect 9840 13340 9880 13380
rect 9840 13240 9880 13280
rect 9950 13340 9990 13380
rect 9950 13240 9990 13280
rect 10360 13340 10400 13380
rect 10360 13240 10400 13280
rect 10470 13340 10510 13380
rect 10470 13240 10510 13280
rect -1440 12770 -1400 12810
rect -1330 12770 -1290 12810
rect -1220 12770 -1180 12810
rect -1110 12770 -1070 12810
rect -1000 12770 -960 12810
rect -860 12770 -820 12810
rect -750 12770 -710 12810
rect -640 12770 -600 12810
rect -410 12770 -370 12810
rect -300 12770 -260 12810
rect -190 12770 -150 12810
rect -80 12770 -40 12810
rect 30 12770 70 12810
rect 250 12770 290 12810
rect 360 12770 400 12810
rect 470 12770 510 12810
rect 580 12770 620 12810
rect 690 12770 730 12810
rect 930 12770 970 12810
rect 1040 12770 1080 12810
rect 1150 12770 1190 12810
rect 1260 12770 1300 12810
rect 1370 12770 1410 12810
rect 1510 12770 1550 12810
rect 1620 12770 1660 12810
rect 1730 12770 1770 12810
rect 2070 12770 2110 12810
rect 2180 12770 2220 12810
rect 2430 12770 2470 12810
rect 2540 12770 2580 12810
rect 2680 12770 2720 12810
rect 2790 12770 2830 12810
rect 2900 12770 2940 12810
rect 3010 12770 3050 12810
rect 3120 12770 3160 12810
rect 3340 12770 3380 12810
rect 3450 12770 3490 12810
rect 3560 12770 3600 12810
rect 3670 12770 3710 12810
rect 3890 12770 3930 12810
rect 4000 12770 4040 12810
rect 4110 12770 4150 12810
rect 4220 12770 4260 12810
rect 4330 12770 4370 12810
rect 4550 12770 4590 12810
rect 4660 12770 4700 12810
rect 4770 12770 4810 12810
rect 5190 12860 5230 12900
rect 5300 12860 5340 12900
rect 5410 12860 5450 12900
rect 5520 12860 5560 12900
rect 5630 12860 5670 12900
rect 5850 12860 5890 12900
rect 5960 12860 6000 12900
rect 6070 12860 6110 12900
rect 6180 12860 6220 12900
rect 6490 12860 6530 12900
rect 6600 12860 6640 12900
rect 6710 12860 6750 12900
rect 6820 12860 6860 12900
rect 6930 12860 6970 12900
rect 7150 12860 7190 12900
rect 7260 12860 7300 12900
rect 7370 12860 7410 12900
rect 7480 12860 7520 12900
rect 7790 12860 7830 12900
rect 7900 12860 7940 12900
rect 8010 12860 8050 12900
rect 8120 12860 8160 12900
rect 8230 12860 8270 12900
rect 8450 12860 8490 12900
rect 8560 12860 8600 12900
rect 8670 12860 8710 12900
rect 8780 12860 8820 12900
rect 4880 12770 4920 12810
rect 9320 12960 9360 13000
rect 9430 12960 9470 13000
rect 9840 12960 9880 13000
rect 9950 12960 9990 13000
rect 10360 12960 10400 13000
rect 10470 12960 10510 13000
rect -620 10170 -580 10210
rect -620 10070 -580 10110
rect -510 10170 -470 10210
rect -510 10070 -470 10110
rect -400 10170 -360 10210
rect -400 10070 -360 10110
rect -100 10170 -60 10210
rect -100 10070 -60 10110
rect 10 10170 50 10210
rect 10 10070 50 10110
rect 120 10170 160 10210
rect 280 10170 320 10210
rect 120 10070 160 10110
rect 280 10070 320 10110
rect 390 10170 430 10210
rect 390 10070 430 10110
rect 500 10170 540 10210
rect 500 10070 540 10110
rect 800 10170 840 10210
rect 800 10070 840 10110
rect 910 10170 950 10210
rect 910 10070 950 10110
rect 1020 10170 1060 10210
rect 1020 10070 1060 10110
rect 1320 10170 1360 10210
rect 1320 10070 1360 10110
rect 1430 10170 1470 10210
rect 1430 10070 1470 10110
rect 1540 10170 1580 10210
rect 1540 10070 1580 10110
rect 1760 10170 1800 10210
rect 1760 10070 1800 10110
rect 1870 10170 1910 10210
rect 1870 10070 1910 10110
rect 2090 10170 2130 10210
rect 2090 10070 2130 10110
rect 2200 10170 2240 10210
rect 2200 10070 2240 10110
rect 2520 10170 2560 10210
rect 2520 10070 2560 10110
rect 2650 10170 2690 10210
rect 2650 10070 2690 10110
rect 2910 10170 2950 10210
rect 2910 10070 2950 10110
rect 3040 10170 3080 10210
rect 3040 10070 3080 10110
rect 3300 10170 3340 10210
rect 3300 10070 3340 10110
rect 3430 10170 3470 10210
rect 3430 10070 3470 10110
rect 3590 10170 3630 10210
rect 3590 10070 3630 10110
rect 3720 10170 3760 10210
rect 3720 10070 3760 10110
rect 5470 8620 5510 8660
rect 5470 8520 5510 8560
rect -620 8370 -580 8410
rect -620 8270 -580 8310
rect -510 8370 -470 8410
rect -510 8270 -470 8310
rect -400 8370 -360 8410
rect -400 8270 -360 8310
rect -100 8370 -60 8410
rect -100 8270 -60 8310
rect 10 8370 50 8410
rect 10 8270 50 8310
rect 120 8370 160 8410
rect 280 8370 320 8410
rect 120 8270 160 8310
rect 280 8270 320 8310
rect 390 8370 430 8410
rect 390 8270 430 8310
rect 500 8370 540 8410
rect 500 8270 540 8310
rect 800 8370 840 8410
rect 800 8270 840 8310
rect 910 8370 950 8410
rect 910 8270 950 8310
rect 1020 8370 1060 8410
rect 1020 8270 1060 8310
rect 1310 8370 1350 8410
rect 1310 8270 1350 8310
rect 1420 8370 1460 8410
rect 1420 8270 1460 8310
rect 1640 8370 1680 8410
rect 1640 8270 1680 8310
rect 1750 8370 1790 8410
rect 1750 8270 1790 8310
rect 1970 8370 2010 8410
rect 1970 8270 2010 8310
rect 2080 8370 2120 8410
rect 2080 8270 2120 8310
rect 2520 8370 2560 8410
rect 2520 8270 2560 8310
rect 2650 8370 2690 8410
rect 2650 8270 2690 8310
rect 2910 8370 2950 8410
rect 2910 8270 2950 8310
rect 3040 8370 3080 8410
rect 3040 8270 3080 8310
rect 3300 8370 3340 8410
rect 3300 8270 3340 8310
rect 3430 8370 3470 8410
rect 3430 8270 3470 8310
rect 3590 8370 3630 8410
rect 3590 8270 3630 8310
rect 3720 8370 3760 8410
rect 3720 8270 3760 8310
rect 3980 8370 4020 8410
rect 3980 8270 4020 8310
rect 4110 8370 4150 8410
rect 4110 8270 4150 8310
rect 5470 8420 5510 8460
rect 5470 8320 5510 8360
rect 5690 8620 5730 8660
rect 5690 8520 5730 8560
rect 5690 8420 5730 8460
rect 5690 8320 5730 8360
rect 5910 8620 5950 8660
rect 5910 8520 5950 8560
rect 5910 8420 5950 8460
rect 5910 8320 5950 8360
rect 6130 8620 6170 8660
rect 6130 8520 6170 8560
rect 6130 8420 6170 8460
rect 6130 8320 6170 8360
rect 6350 8620 6390 8660
rect 6550 8620 6590 8660
rect 6350 8520 6390 8560
rect 6550 8520 6590 8560
rect 6350 8420 6390 8460
rect 6550 8420 6590 8460
rect 6350 8320 6390 8360
rect 6550 8320 6590 8360
rect 6770 8620 6810 8660
rect 6770 8520 6810 8560
rect 6770 8420 6810 8460
rect 6770 8320 6810 8360
rect 6990 8620 7030 8660
rect 6990 8520 7030 8560
rect 6990 8420 7030 8460
rect 6990 8320 7030 8360
rect 7210 8620 7250 8660
rect 7210 8520 7250 8560
rect 7210 8420 7250 8460
rect 7210 8320 7250 8360
rect 7430 8620 7470 8660
rect 7630 8620 7670 8660
rect 7430 8520 7470 8560
rect 7630 8520 7670 8560
rect 7430 8420 7470 8460
rect 7630 8420 7670 8460
rect 7430 8320 7470 8360
rect 7630 8320 7670 8360
rect 7850 8620 7890 8660
rect 7850 8520 7890 8560
rect 7850 8420 7890 8460
rect 7850 8320 7890 8360
rect 8070 8620 8110 8660
rect 8070 8520 8110 8560
rect 8070 8420 8110 8460
rect 8070 8320 8110 8360
rect 8290 8620 8330 8660
rect 8290 8520 8330 8560
rect 8290 8420 8330 8460
rect 8290 8320 8330 8360
rect 8510 8620 8550 8660
rect 8510 8520 8550 8560
rect 8510 8420 8550 8460
rect 8510 8320 8550 8360
rect 5530 5980 5570 6030
rect 5530 5840 5570 5890
rect 5730 5980 5770 6030
rect 5730 5840 5770 5890
rect 5930 5980 5970 6030
rect 5930 5840 5970 5890
rect 6130 5980 6170 6030
rect 6130 5840 6170 5890
rect 6330 5980 6370 6030
rect 6330 5840 6370 5890
rect 6530 5980 6570 6030
rect 6530 5840 6570 5890
rect 6730 5980 6770 6030
rect 6730 5840 6770 5890
rect 6930 5980 6970 6030
rect 6930 5840 6970 5890
rect 7130 5980 7170 6030
rect 7130 5840 7170 5890
rect 7330 5980 7370 6030
rect 7330 5840 7370 5890
rect 7530 5980 7570 6030
rect 7530 5840 7570 5890
rect 5580 5300 5620 5340
rect 5710 5300 5750 5340
rect 5840 5300 5880 5340
rect 5970 5300 6010 5340
rect 6100 5300 6140 5340
rect 6230 5300 6270 5340
rect 6360 5300 6400 5340
rect 6720 5300 6760 5340
rect 6850 5300 6890 5340
rect 6980 5300 7020 5340
rect 7110 5300 7150 5340
rect 7240 5300 7280 5340
rect 7370 5300 7410 5340
rect 7500 5300 7540 5340
rect 7860 5300 7900 5340
rect 7990 5300 8030 5340
rect 8120 5300 8160 5340
rect 8250 5300 8290 5340
rect 8380 5300 8420 5340
rect 8510 5300 8550 5340
rect 8640 5300 8680 5340
rect -1610 3700 -1570 3740
rect -1490 3700 -1450 3740
rect -1370 3700 -1330 3740
rect -1250 3700 -1210 3740
rect -1130 3700 -1090 3740
rect -1010 3700 -970 3740
rect -890 3700 -850 3740
rect -770 3700 -730 3740
rect -650 3700 -610 3740
rect -530 3700 -490 3740
rect -410 3700 -370 3740
rect 950 3700 990 3740
rect 1070 3700 1110 3740
rect 1190 3700 1230 3740
rect 1310 3700 1350 3740
rect 1430 3700 1470 3740
rect 1550 3700 1590 3740
rect 1670 3700 1710 3740
rect 1790 3700 1830 3740
rect 1910 3700 1950 3740
rect 2030 3700 2070 3740
rect 2150 3700 2190 3740
rect -2230 3090 -2190 3130
rect -2230 2990 -2190 3030
rect -2230 2890 -2190 2930
rect -2230 2790 -2190 2830
rect -2230 2690 -2190 2730
rect -1150 3090 -1110 3130
rect -990 3090 -950 3130
rect -1150 2990 -1110 3030
rect -990 2990 -950 3030
rect -1150 2890 -1110 2930
rect -990 2890 -950 2930
rect -1150 2790 -1110 2830
rect -990 2790 -950 2830
rect -1150 2690 -1110 2730
rect -990 2690 -950 2730
rect 90 3090 130 3130
rect 90 2990 130 3030
rect 90 2890 130 2930
rect 90 2790 130 2830
rect 90 2690 130 2730
rect 450 3090 490 3130
rect 450 2990 490 3030
rect 450 2890 490 2930
rect 450 2790 490 2830
rect 450 2690 490 2730
rect 1530 3090 1570 3130
rect 1690 3090 1730 3130
rect 1530 2990 1570 3030
rect 1690 2990 1730 3030
rect 1530 2890 1570 2930
rect 1690 2890 1730 2930
rect 1530 2790 1570 2830
rect 1690 2790 1730 2830
rect 1530 2690 1570 2730
rect 1690 2690 1730 2730
rect 2770 3090 2810 3130
rect 2770 2990 2810 3030
rect 2770 2890 2810 2930
rect 2770 2790 2810 2830
rect 2770 2690 2810 2730
rect -1810 2180 -1770 2220
rect -1810 2080 -1770 2120
rect 270 2180 310 2220
rect 270 2080 310 2120
rect 2350 2180 2390 2220
rect 2350 2080 2390 2120
<< pdiffc >>
rect -1280 12450 -1240 12490
rect -1170 12450 -1130 12490
rect -860 12450 -820 12490
rect -750 12450 -710 12490
rect -640 12450 -600 12490
rect -190 12450 -150 12490
rect -80 12450 -40 12490
rect 30 12450 70 12490
rect 250 12450 290 12490
rect 360 12450 400 12490
rect 470 12450 510 12490
rect 580 12450 620 12490
rect 1090 12450 1130 12490
rect 1200 12450 1240 12490
rect 1510 12450 1550 12490
rect 1620 12450 1660 12490
rect 1730 12450 1770 12490
rect 1960 12450 2000 12490
rect 2070 12450 2110 12490
rect 2180 12450 2220 12490
rect 2320 12450 2360 12490
rect 2430 12450 2470 12490
rect 2540 12450 2580 12490
rect 2900 12450 2940 12490
rect 3010 12450 3050 12490
rect 3120 12450 3160 12490
rect 3340 12450 3380 12490
rect 3450 12450 3490 12490
rect 3560 12450 3600 12490
rect 3960 12450 4000 12490
rect 4070 12450 4110 12490
rect 4300 12450 4340 12490
rect 4410 12450 4450 12490
rect 4520 12450 4560 12490
rect 4660 12450 4700 12490
rect 4770 12450 4810 12490
rect 4880 12450 4920 12490
rect 5260 12450 5300 12490
rect 5370 12450 5410 12490
rect 5600 12450 5640 12490
rect 5710 12450 5750 12490
rect 5820 12450 5860 12490
rect 5960 12450 6000 12490
rect 6070 12450 6110 12490
rect 6180 12450 6220 12490
rect 6560 12450 6600 12490
rect 6670 12450 6710 12490
rect 6900 12450 6940 12490
rect 7010 12450 7050 12490
rect 7120 12450 7160 12490
rect 7260 12450 7300 12490
rect 7370 12450 7410 12490
rect 7480 12450 7520 12490
rect 7860 12450 7900 12490
rect 7970 12450 8010 12490
rect 8200 12450 8240 12490
rect 8310 12450 8350 12490
rect 8420 12450 8460 12490
rect 8560 12450 8600 12490
rect 8670 12450 8710 12490
rect 8780 12450 8820 12490
rect 9320 12300 9360 12340
rect 9320 12200 9360 12240
rect 9430 12300 9470 12340
rect 9430 12200 9470 12240
rect 9840 12300 9880 12340
rect 9840 12200 9880 12240
rect 9950 12300 9990 12340
rect 9950 12200 9990 12240
rect 10360 12300 10400 12340
rect 10360 12200 10400 12240
rect 10470 12300 10510 12340
rect 10470 12200 10510 12240
rect 9320 11920 9360 11960
rect 9320 11820 9360 11860
rect 9320 11720 9360 11760
rect 9320 11620 9360 11660
rect 9430 11920 9470 11960
rect 9430 11820 9470 11860
rect 9430 11720 9470 11760
rect 9430 11620 9470 11660
rect 9840 11920 9880 11960
rect 9840 11820 9880 11860
rect 9840 11720 9880 11760
rect 9840 11620 9880 11660
rect 9950 11920 9990 11960
rect 9950 11820 9990 11860
rect 9950 11720 9990 11760
rect 9950 11620 9990 11660
rect 10360 11920 10400 11960
rect 10360 11820 10400 11860
rect 10360 11720 10400 11760
rect 10360 11620 10400 11660
rect 10470 11920 10510 11960
rect 10470 11820 10510 11860
rect 10470 11720 10510 11760
rect 10470 11620 10510 11660
rect 9320 11230 9360 11270
rect 9320 11130 9360 11170
rect 9320 11030 9360 11070
rect 9320 10930 9360 10970
rect 9700 11230 9740 11270
rect 9700 11130 9740 11170
rect 9700 11030 9740 11070
rect 9700 10930 9740 10970
rect 9840 11230 9880 11270
rect 9840 11130 9880 11170
rect 9840 11030 9880 11070
rect 9840 10930 9880 10970
rect 10220 11230 10260 11270
rect 10220 11130 10260 11170
rect 10220 11030 10260 11070
rect 10220 10930 10260 10970
rect 10360 11230 10400 11270
rect 10360 11130 10400 11170
rect 10360 11030 10400 11070
rect 10360 10930 10400 10970
rect 10740 11230 10780 11270
rect 10740 11130 10780 11170
rect 10740 11030 10780 11070
rect 10740 10930 10780 10970
rect 10880 11230 10920 11270
rect 10880 11130 10920 11170
rect 10880 11030 10920 11070
rect 10880 10930 10920 10970
rect 11260 11230 11300 11270
rect 11260 11130 11300 11170
rect 11260 11030 11300 11070
rect 11260 10930 11300 10970
rect -620 9750 -580 9790
rect -620 9650 -580 9690
rect -620 9550 -580 9590
rect -620 9450 -580 9490
rect -510 9750 -470 9790
rect -510 9650 -470 9690
rect -510 9550 -470 9590
rect -510 9450 -470 9490
rect -400 9750 -360 9790
rect -400 9650 -360 9690
rect -400 9550 -360 9590
rect -400 9450 -360 9490
rect -100 9750 -60 9790
rect -100 9650 -60 9690
rect -100 9550 -60 9590
rect -100 9450 -60 9490
rect 10 9750 50 9790
rect 10 9650 50 9690
rect 10 9550 50 9590
rect 10 9450 50 9490
rect 120 9750 160 9790
rect 280 9750 320 9790
rect 120 9650 160 9690
rect 280 9650 320 9690
rect 120 9550 160 9590
rect 280 9550 320 9590
rect 120 9450 160 9490
rect 280 9450 320 9490
rect 390 9750 430 9790
rect 390 9650 430 9690
rect 390 9550 430 9590
rect 390 9450 430 9490
rect 500 9750 540 9790
rect 500 9650 540 9690
rect 500 9550 540 9590
rect 500 9450 540 9490
rect 800 9750 840 9790
rect 800 9650 840 9690
rect 800 9550 840 9590
rect 800 9450 840 9490
rect 910 9750 950 9790
rect 910 9650 950 9690
rect 910 9550 950 9590
rect 910 9450 950 9490
rect 1020 9750 1060 9790
rect 1020 9650 1060 9690
rect 1020 9550 1060 9590
rect 1020 9450 1060 9490
rect 1320 9750 1360 9790
rect 1320 9650 1360 9690
rect 1320 9550 1360 9590
rect 1320 9450 1360 9490
rect 1430 9750 1470 9790
rect 1430 9650 1470 9690
rect 1430 9550 1470 9590
rect 1430 9450 1470 9490
rect 1540 9750 1580 9790
rect 1540 9650 1580 9690
rect 1540 9550 1580 9590
rect 1540 9450 1580 9490
rect 1760 9750 1800 9790
rect 1760 9650 1800 9690
rect 1760 9550 1800 9590
rect 1760 9450 1800 9490
rect 1870 9750 1910 9790
rect 1870 9650 1910 9690
rect 1870 9550 1910 9590
rect 1870 9450 1910 9490
rect 2090 9750 2130 9790
rect 2090 9650 2130 9690
rect 2090 9550 2130 9590
rect 2090 9450 2130 9490
rect 2200 9750 2240 9790
rect 2200 9650 2240 9690
rect 2200 9550 2240 9590
rect 2200 9450 2240 9490
rect 2520 9750 2560 9790
rect 2520 9650 2560 9690
rect 2520 9550 2560 9590
rect 2520 9450 2560 9490
rect 2650 9750 2690 9790
rect 2650 9650 2690 9690
rect 2650 9550 2690 9590
rect 2650 9450 2690 9490
rect 2910 9750 2950 9790
rect 2910 9650 2950 9690
rect 2910 9550 2950 9590
rect 2910 9450 2950 9490
rect 3040 9750 3080 9790
rect 3040 9650 3080 9690
rect 3040 9550 3080 9590
rect 3040 9450 3080 9490
rect 3300 9750 3340 9790
rect 3300 9650 3340 9690
rect 3300 9550 3340 9590
rect 3300 9450 3340 9490
rect 3430 9750 3470 9790
rect 3430 9650 3470 9690
rect 3430 9550 3470 9590
rect 3430 9450 3470 9490
rect 3590 9750 3630 9790
rect 3590 9650 3630 9690
rect 3590 9550 3630 9590
rect 3590 9450 3630 9490
rect 3720 9750 3760 9790
rect 3720 9650 3760 9690
rect 3720 9550 3760 9590
rect 3720 9450 3760 9490
rect 3980 9750 4020 9790
rect 3980 9650 4020 9690
rect 3980 9550 4020 9590
rect 3980 9450 4020 9490
rect 4110 9750 4150 9790
rect 4110 9650 4150 9690
rect 4110 9550 4150 9590
rect 4110 9450 4150 9490
rect 5670 9720 5710 9760
rect 5670 9620 5710 9660
rect 5670 9520 5710 9560
rect 5670 9420 5710 9460
rect 5890 9720 5930 9760
rect 5890 9620 5930 9660
rect 5890 9520 5930 9560
rect 5890 9420 5930 9460
rect 6110 9720 6150 9760
rect 6110 9620 6150 9660
rect 6110 9520 6150 9560
rect 6110 9420 6150 9460
rect 6330 9720 6370 9760
rect 6330 9620 6370 9660
rect 6330 9520 6370 9560
rect 6330 9420 6370 9460
rect 6550 9720 6590 9760
rect 6550 9620 6590 9660
rect 6550 9520 6590 9560
rect 6550 9420 6590 9460
rect 6770 9720 6810 9760
rect 6770 9620 6810 9660
rect 6770 9520 6810 9560
rect 6770 9420 6810 9460
rect 6990 9720 7030 9760
rect 7190 9720 7230 9760
rect 6990 9620 7030 9660
rect 7190 9620 7230 9660
rect 6990 9520 7030 9560
rect 7190 9520 7230 9560
rect 6990 9420 7030 9460
rect 7190 9420 7230 9460
rect 7410 9720 7450 9760
rect 7410 9620 7450 9660
rect 7410 9520 7450 9560
rect 7410 9420 7450 9460
rect 7630 9720 7670 9760
rect 7630 9620 7670 9660
rect 7630 9520 7670 9560
rect 7630 9420 7670 9460
rect 7850 9720 7890 9760
rect 7850 9620 7890 9660
rect 7850 9520 7890 9560
rect 7850 9420 7890 9460
rect 8070 9720 8110 9760
rect 8070 9620 8110 9660
rect 8070 9520 8110 9560
rect 8070 9420 8110 9460
rect 8290 9720 8330 9760
rect 8290 9620 8330 9660
rect 8290 9520 8330 9560
rect 8290 9420 8330 9460
rect 8510 9720 8550 9760
rect 8510 9620 8550 9660
rect 8510 9520 8550 9560
rect 8510 9420 8550 9460
rect -620 8990 -580 9030
rect -620 8890 -580 8930
rect -620 8790 -580 8830
rect -620 8690 -580 8730
rect -510 8990 -470 9030
rect -510 8890 -470 8930
rect -510 8790 -470 8830
rect -510 8690 -470 8730
rect -400 8990 -360 9030
rect -400 8890 -360 8930
rect -400 8790 -360 8830
rect -400 8690 -360 8730
rect -100 8990 -60 9030
rect -100 8890 -60 8930
rect -100 8790 -60 8830
rect -100 8690 -60 8730
rect 10 8990 50 9030
rect 10 8890 50 8930
rect 10 8790 50 8830
rect 10 8690 50 8730
rect 120 8990 160 9030
rect 280 8990 320 9030
rect 120 8890 160 8930
rect 280 8890 320 8930
rect 120 8790 160 8830
rect 280 8790 320 8830
rect 120 8690 160 8730
rect 280 8690 320 8730
rect 390 8990 430 9030
rect 390 8890 430 8930
rect 390 8790 430 8830
rect 390 8690 430 8730
rect 500 8990 540 9030
rect 500 8890 540 8930
rect 500 8790 540 8830
rect 500 8690 540 8730
rect 800 8990 840 9030
rect 800 8890 840 8930
rect 800 8790 840 8830
rect 800 8690 840 8730
rect 910 8990 950 9030
rect 910 8890 950 8930
rect 910 8790 950 8830
rect 910 8690 950 8730
rect 1020 8990 1060 9030
rect 1020 8890 1060 8930
rect 1020 8790 1060 8830
rect 1020 8690 1060 8730
rect 1310 8990 1350 9030
rect 1310 8890 1350 8930
rect 1310 8790 1350 8830
rect 1310 8690 1350 8730
rect 1420 8990 1460 9030
rect 1420 8890 1460 8930
rect 1420 8790 1460 8830
rect 1420 8690 1460 8730
rect 1640 8990 1680 9030
rect 1640 8890 1680 8930
rect 1640 8790 1680 8830
rect 1640 8690 1680 8730
rect 1750 8990 1790 9030
rect 1750 8890 1790 8930
rect 1750 8790 1790 8830
rect 1750 8690 1790 8730
rect 1970 8990 2010 9030
rect 1970 8890 2010 8930
rect 1970 8790 2010 8830
rect 1970 8690 2010 8730
rect 2080 8990 2120 9030
rect 2080 8890 2120 8930
rect 2080 8790 2120 8830
rect 2080 8690 2120 8730
rect 2520 8990 2560 9030
rect 2520 8890 2560 8930
rect 2520 8790 2560 8830
rect 2520 8690 2560 8730
rect 2650 8990 2690 9030
rect 2650 8890 2690 8930
rect 2650 8790 2690 8830
rect 2650 8690 2690 8730
rect 2910 8990 2950 9030
rect 2910 8890 2950 8930
rect 2910 8790 2950 8830
rect 2910 8690 2950 8730
rect 3040 8990 3080 9030
rect 3040 8890 3080 8930
rect 3040 8790 3080 8830
rect 3040 8690 3080 8730
rect 3300 8990 3340 9030
rect 3300 8890 3340 8930
rect 3300 8790 3340 8830
rect 3300 8690 3340 8730
rect 3430 8990 3470 9030
rect 3430 8890 3470 8930
rect 3430 8790 3470 8830
rect 3430 8690 3470 8730
rect 3590 8990 3630 9030
rect 3590 8890 3630 8930
rect 3590 8790 3630 8830
rect 3590 8690 3630 8730
rect 3720 8990 3760 9030
rect 3720 8890 3760 8930
rect 3720 8790 3760 8830
rect 3720 8690 3760 8730
rect -1340 6800 -1300 6840
rect -1340 6700 -1300 6740
rect -1230 6800 -1190 6840
rect -1230 6700 -1190 6740
rect -1120 6800 -1080 6840
rect -1120 6700 -1080 6740
rect -1010 6800 -970 6840
rect -1010 6700 -970 6740
rect -900 6800 -860 6840
rect -900 6700 -860 6740
rect -790 6800 -750 6840
rect -790 6700 -750 6740
rect -680 6800 -640 6840
rect -680 6700 -640 6740
rect -570 6800 -530 6840
rect -570 6700 -530 6740
rect -460 6800 -420 6840
rect -460 6700 -420 6740
rect -350 6800 -310 6840
rect -350 6700 -310 6740
rect -240 6800 -200 6840
rect -240 6700 -200 6740
rect -130 6800 -90 6840
rect -130 6700 -90 6740
rect -20 6800 20 6840
rect -20 6700 20 6740
rect 560 6800 600 6840
rect 560 6700 600 6740
rect 670 6800 710 6840
rect 670 6700 710 6740
rect 780 6800 820 6840
rect 780 6700 820 6740
rect 890 6800 930 6840
rect 890 6700 930 6740
rect 1000 6800 1040 6840
rect 1000 6700 1040 6740
rect 1110 6800 1150 6840
rect 1110 6700 1150 6740
rect 1220 6800 1260 6840
rect 1220 6700 1260 6740
rect 1330 6800 1370 6840
rect 1330 6700 1370 6740
rect 1440 6800 1480 6840
rect 1440 6700 1480 6740
rect 1550 6800 1590 6840
rect 1550 6700 1590 6740
rect 1660 6800 1700 6840
rect 1660 6700 1700 6740
rect 1770 6800 1810 6840
rect 1770 6700 1810 6740
rect 1880 6800 1920 6840
rect 1880 6700 1920 6740
rect -1350 6200 -1310 6240
rect -1350 6100 -1310 6140
rect -1350 6000 -1310 6040
rect -1350 5900 -1310 5940
rect -1350 5800 -1310 5840
rect -1350 5700 -1310 5740
rect -1170 6200 -1130 6240
rect -1170 6100 -1130 6140
rect -1170 6000 -1130 6040
rect -1170 5900 -1130 5940
rect -1170 5800 -1130 5840
rect -1170 5700 -1130 5740
rect -990 6200 -950 6240
rect -990 6100 -950 6140
rect -990 6000 -950 6040
rect -990 5900 -950 5940
rect -990 5800 -950 5840
rect -990 5700 -950 5740
rect -810 6200 -770 6240
rect -810 6100 -770 6140
rect -810 6000 -770 6040
rect -810 5900 -770 5940
rect -810 5800 -770 5840
rect -810 5700 -770 5740
rect -630 6200 -590 6240
rect -630 6100 -590 6140
rect -630 6000 -590 6040
rect -630 5900 -590 5940
rect -630 5800 -590 5840
rect -630 5700 -590 5740
rect -450 6200 -410 6240
rect -450 6100 -410 6140
rect -450 6000 -410 6040
rect -450 5900 -410 5940
rect -450 5800 -410 5840
rect -450 5700 -410 5740
rect -270 6200 -230 6240
rect -270 6100 -230 6140
rect -270 6000 -230 6040
rect -270 5900 -230 5940
rect -270 5800 -230 5840
rect -270 5700 -230 5740
rect -90 6200 -50 6240
rect -90 6100 -50 6140
rect -90 6000 -50 6040
rect -90 5900 -50 5940
rect -90 5800 -50 5840
rect -90 5700 -50 5740
rect 90 6200 130 6240
rect 90 6100 130 6140
rect 90 6000 130 6040
rect 90 5900 130 5940
rect 90 5800 130 5840
rect 90 5700 130 5740
rect 270 6200 310 6240
rect 270 6100 310 6140
rect 270 6000 310 6040
rect 270 5900 310 5940
rect 270 5800 310 5840
rect 270 5700 310 5740
rect 450 6200 490 6240
rect 450 6100 490 6140
rect 450 6000 490 6040
rect 450 5900 490 5940
rect 450 5800 490 5840
rect 450 5700 490 5740
rect 630 6200 670 6240
rect 630 6100 670 6140
rect 630 6000 670 6040
rect 630 5900 670 5940
rect 630 5800 670 5840
rect 630 5700 670 5740
rect 810 6200 850 6240
rect 810 6100 850 6140
rect 810 6000 850 6040
rect 810 5900 850 5940
rect 810 5800 850 5840
rect 810 5700 850 5740
rect 990 6200 1030 6240
rect 990 6100 1030 6140
rect 990 6000 1030 6040
rect 990 5900 1030 5940
rect 990 5800 1030 5840
rect 990 5700 1030 5740
rect 1170 6200 1210 6240
rect 1170 6100 1210 6140
rect 1170 6000 1210 6040
rect 1170 5900 1210 5940
rect 1170 5800 1210 5840
rect 1170 5700 1210 5740
rect 1350 6200 1390 6240
rect 1350 6100 1390 6140
rect 1350 6000 1390 6040
rect 1350 5900 1390 5940
rect 1350 5800 1390 5840
rect 1350 5700 1390 5740
rect 1530 6200 1570 6240
rect 1530 6100 1570 6140
rect 1530 6000 1570 6040
rect 1530 5900 1570 5940
rect 1530 5800 1570 5840
rect 1530 5700 1570 5740
rect 1710 6200 1750 6240
rect 1710 6100 1750 6140
rect 1710 6000 1750 6040
rect 1710 5900 1750 5940
rect 1710 5800 1750 5840
rect 1710 5700 1750 5740
rect 1890 6200 1930 6240
rect 1890 6100 1930 6140
rect 1890 6000 1930 6040
rect 1890 5900 1930 5940
rect 2520 6000 2560 6040
rect 2520 5900 2560 5940
rect 2630 6000 2670 6040
rect 2630 5900 2670 5940
rect 2740 6000 2780 6040
rect 2740 5900 2780 5940
rect 2850 6000 2890 6040
rect 2850 5900 2890 5940
rect 2960 6000 3000 6040
rect 2960 5900 3000 5940
rect 1890 5800 1930 5840
rect 1890 5700 1930 5740
rect 5580 4720 5620 4760
rect -2450 4640 -2410 4680
rect -2450 4540 -2410 4580
rect -2330 4640 -2290 4680
rect -2330 4540 -2290 4580
rect -2210 4640 -2170 4680
rect -2210 4540 -2170 4580
rect -2090 4640 -2050 4680
rect -2090 4540 -2050 4580
rect -1970 4640 -1930 4680
rect -1970 4540 -1930 4580
rect -1850 4640 -1810 4680
rect -1850 4540 -1810 4580
rect -1730 4640 -1690 4680
rect -1730 4540 -1690 4580
rect -1610 4640 -1570 4680
rect -1610 4540 -1570 4580
rect -1490 4640 -1450 4680
rect -1490 4540 -1450 4580
rect -1370 4640 -1330 4680
rect -1370 4540 -1330 4580
rect -1250 4640 -1210 4680
rect -1250 4540 -1210 4580
rect -1130 4640 -1090 4680
rect -1130 4540 -1090 4580
rect -1010 4640 -970 4680
rect -1010 4540 -970 4580
rect -890 4640 -850 4680
rect -890 4540 -850 4580
rect -770 4640 -730 4680
rect -770 4540 -730 4580
rect -650 4640 -610 4680
rect -650 4540 -610 4580
rect -530 4640 -490 4680
rect -530 4540 -490 4580
rect -410 4640 -370 4680
rect -410 4540 -370 4580
rect -290 4640 -250 4680
rect -290 4540 -250 4580
rect -170 4640 -130 4680
rect -170 4540 -130 4580
rect -50 4640 -10 4680
rect -50 4540 -10 4580
rect 590 4640 630 4680
rect 590 4540 630 4580
rect 710 4640 750 4680
rect 710 4540 750 4580
rect 830 4640 870 4680
rect 830 4540 870 4580
rect 950 4640 990 4680
rect 950 4540 990 4580
rect 1070 4640 1110 4680
rect 1070 4540 1110 4580
rect 1190 4640 1230 4680
rect 1190 4540 1230 4580
rect 1310 4640 1350 4680
rect 1310 4540 1350 4580
rect 1430 4640 1470 4680
rect 1430 4540 1470 4580
rect 1550 4640 1590 4680
rect 1550 4540 1590 4580
rect 1670 4640 1710 4680
rect 1670 4540 1710 4580
rect 1790 4640 1830 4680
rect 1790 4540 1830 4580
rect 1910 4640 1950 4680
rect 1910 4540 1950 4580
rect 2030 4640 2070 4680
rect 2030 4540 2070 4580
rect 2150 4640 2190 4680
rect 2150 4540 2190 4580
rect 2270 4640 2310 4680
rect 2270 4540 2310 4580
rect 2390 4640 2430 4680
rect 2390 4540 2430 4580
rect 2510 4640 2550 4680
rect 2510 4540 2550 4580
rect 2630 4640 2670 4680
rect 2630 4540 2670 4580
rect 2750 4640 2790 4680
rect 2750 4540 2790 4580
rect 2870 4640 2910 4680
rect 2870 4540 2910 4580
rect 2990 4640 3030 4680
rect 5580 4620 5620 4660
rect 5710 4720 5750 4760
rect 5710 4620 5750 4660
rect 5840 4720 5880 4760
rect 5840 4620 5880 4660
rect 5970 4720 6010 4760
rect 5970 4620 6010 4660
rect 6100 4720 6140 4760
rect 6100 4620 6140 4660
rect 6230 4720 6270 4760
rect 6230 4620 6270 4660
rect 6360 4720 6400 4760
rect 6360 4620 6400 4660
rect 6720 4720 6760 4760
rect 6720 4620 6760 4660
rect 6850 4720 6890 4760
rect 6850 4620 6890 4660
rect 6980 4720 7020 4760
rect 6980 4620 7020 4660
rect 7110 4720 7150 4760
rect 7110 4620 7150 4660
rect 7240 4720 7280 4760
rect 7240 4620 7280 4660
rect 7370 4720 7410 4760
rect 7370 4620 7410 4660
rect 7500 4720 7540 4760
rect 7500 4620 7540 4660
rect 7860 4720 7900 4760
rect 7860 4620 7900 4660
rect 7990 4720 8030 4760
rect 7990 4620 8030 4660
rect 8120 4720 8160 4760
rect 8120 4620 8160 4660
rect 8250 4720 8290 4760
rect 8250 4620 8290 4660
rect 8380 4720 8420 4760
rect 8380 4620 8420 4660
rect 8510 4720 8550 4760
rect 8510 4620 8550 4660
rect 8640 4720 8680 4760
rect 8640 4620 8680 4660
rect 2990 4540 3030 4580
rect 5650 4070 5690 4110
rect 5650 3970 5690 4010
rect 5650 3870 5690 3910
rect 5650 3770 5690 3810
rect 5650 3670 5690 3710
rect 5850 4070 5890 4110
rect 5850 3970 5890 4010
rect 5850 3870 5890 3910
rect 5850 3770 5890 3810
rect 5850 3670 5890 3710
rect 6050 4070 6090 4110
rect 6050 3970 6090 4010
rect 6050 3870 6090 3910
rect 6050 3770 6090 3810
rect 6050 3670 6090 3710
rect 6250 4070 6290 4110
rect 6250 3970 6290 4010
rect 6250 3870 6290 3910
rect 6250 3770 6290 3810
rect 6250 3670 6290 3710
rect 6450 4070 6490 4110
rect 6450 3970 6490 4010
rect 6450 3870 6490 3910
rect 6450 3770 6490 3810
rect 6450 3670 6490 3710
rect 6650 4070 6690 4110
rect 6650 3970 6690 4010
rect 6650 3870 6690 3910
rect 6650 3770 6690 3810
rect 6650 3670 6690 3710
rect 6850 4070 6890 4110
rect 6850 3970 6890 4010
rect 6850 3870 6890 3910
rect 6850 3770 6890 3810
rect 6850 3670 6890 3710
rect 7050 4070 7090 4110
rect 7050 3970 7090 4010
rect 7050 3870 7090 3910
rect 7050 3770 7090 3810
rect 7050 3670 7090 3710
rect 7250 4070 7290 4110
rect 7250 3970 7290 4010
rect 7250 3870 7290 3910
rect 7250 3770 7290 3810
rect 7250 3670 7290 3710
rect 7450 4070 7490 4110
rect 7450 3970 7490 4010
rect 7450 3870 7490 3910
rect 7450 3770 7490 3810
rect 7450 3670 7490 3710
rect 7650 4070 7690 4110
rect 7650 3970 7690 4010
rect 7650 3870 7690 3910
rect 7650 3770 7690 3810
rect 7650 3670 7690 3710
rect -1358 1164 -1324 1198
rect -1268 1164 -1234 1198
rect -1178 1164 -1144 1198
rect -1088 1164 -1054 1198
rect -998 1164 -964 1198
rect -908 1164 -874 1198
rect -818 1164 -784 1198
rect -1358 1074 -1324 1108
rect -1268 1074 -1234 1108
rect -1178 1074 -1144 1108
rect -1088 1074 -1054 1108
rect -998 1074 -964 1108
rect -908 1074 -874 1108
rect -818 1074 -784 1108
rect -1358 984 -1324 1018
rect -1268 984 -1234 1018
rect -1178 984 -1144 1018
rect -1088 984 -1054 1018
rect -998 984 -964 1018
rect -908 984 -874 1018
rect -818 984 -784 1018
rect -1358 894 -1324 928
rect -1268 894 -1234 928
rect -1178 894 -1144 928
rect -1088 894 -1054 928
rect -998 894 -964 928
rect -908 894 -874 928
rect -818 894 -784 928
rect -1358 804 -1324 838
rect -1268 804 -1234 838
rect -1178 804 -1144 838
rect -1088 804 -1054 838
rect -998 804 -964 838
rect -908 804 -874 838
rect -818 804 -784 838
rect -1358 714 -1324 748
rect -1268 714 -1234 748
rect -1178 714 -1144 748
rect -1088 714 -1054 748
rect -998 714 -964 748
rect -908 714 -874 748
rect -818 714 -784 748
rect -1358 624 -1324 658
rect -1268 624 -1234 658
rect -1178 624 -1144 658
rect -1088 624 -1054 658
rect -998 624 -964 658
rect -908 624 -874 658
rect -818 624 -784 658
rect 2 1164 36 1198
rect 92 1164 126 1198
rect 182 1164 216 1198
rect 272 1164 306 1198
rect 362 1164 396 1198
rect 452 1164 486 1198
rect 542 1164 576 1198
rect 2 1074 36 1108
rect 92 1074 126 1108
rect 182 1074 216 1108
rect 272 1074 306 1108
rect 362 1074 396 1108
rect 452 1074 486 1108
rect 542 1074 576 1108
rect 2 984 36 1018
rect 92 984 126 1018
rect 182 984 216 1018
rect 272 984 306 1018
rect 362 984 396 1018
rect 452 984 486 1018
rect 542 984 576 1018
rect 2 894 36 928
rect 92 894 126 928
rect 182 894 216 928
rect 272 894 306 928
rect 362 894 396 928
rect 452 894 486 928
rect 542 894 576 928
rect 2 804 36 838
rect 92 804 126 838
rect 182 804 216 838
rect 272 804 306 838
rect 362 804 396 838
rect 452 804 486 838
rect 542 804 576 838
rect 2 714 36 748
rect 92 714 126 748
rect 182 714 216 748
rect 272 714 306 748
rect 362 714 396 748
rect 452 714 486 748
rect 542 714 576 748
rect 2 624 36 658
rect 92 624 126 658
rect 182 624 216 658
rect 272 624 306 658
rect 362 624 396 658
rect 452 624 486 658
rect 542 624 576 658
rect 1362 1164 1396 1198
rect 1452 1164 1486 1198
rect 1542 1164 1576 1198
rect 1632 1164 1666 1198
rect 1722 1164 1756 1198
rect 1812 1164 1846 1198
rect 1902 1164 1936 1198
rect 1362 1074 1396 1108
rect 1452 1074 1486 1108
rect 1542 1074 1576 1108
rect 1632 1074 1666 1108
rect 1722 1074 1756 1108
rect 1812 1074 1846 1108
rect 1902 1074 1936 1108
rect 1362 984 1396 1018
rect 1452 984 1486 1018
rect 1542 984 1576 1018
rect 1632 984 1666 1018
rect 1722 984 1756 1018
rect 1812 984 1846 1018
rect 1902 984 1936 1018
rect 1362 894 1396 928
rect 1452 894 1486 928
rect 1542 894 1576 928
rect 1632 894 1666 928
rect 1722 894 1756 928
rect 1812 894 1846 928
rect 1902 894 1936 928
rect 1362 804 1396 838
rect 1452 804 1486 838
rect 1542 804 1576 838
rect 1632 804 1666 838
rect 1722 804 1756 838
rect 1812 804 1846 838
rect 1902 804 1936 838
rect 1362 714 1396 748
rect 1452 714 1486 748
rect 1542 714 1576 748
rect 1632 714 1666 748
rect 1722 714 1756 748
rect 1812 714 1846 748
rect 1902 714 1936 748
rect 1362 624 1396 658
rect 1452 624 1486 658
rect 1542 624 1576 658
rect 1632 624 1666 658
rect 1722 624 1756 658
rect 1812 624 1846 658
rect 1902 624 1936 658
rect -1358 -196 -1324 -162
rect -1268 -196 -1234 -162
rect -1178 -196 -1144 -162
rect -1088 -196 -1054 -162
rect -998 -196 -964 -162
rect -908 -196 -874 -162
rect -818 -196 -784 -162
rect -1358 -286 -1324 -252
rect -1268 -286 -1234 -252
rect -1178 -286 -1144 -252
rect -1088 -286 -1054 -252
rect -998 -286 -964 -252
rect -908 -286 -874 -252
rect -818 -286 -784 -252
rect -1358 -376 -1324 -342
rect -1268 -376 -1234 -342
rect -1178 -376 -1144 -342
rect -1088 -376 -1054 -342
rect -998 -376 -964 -342
rect -908 -376 -874 -342
rect -818 -376 -784 -342
rect -1358 -466 -1324 -432
rect -1268 -466 -1234 -432
rect -1178 -466 -1144 -432
rect -1088 -466 -1054 -432
rect -998 -466 -964 -432
rect -908 -466 -874 -432
rect -818 -466 -784 -432
rect -1358 -556 -1324 -522
rect -1268 -556 -1234 -522
rect -1178 -556 -1144 -522
rect -1088 -556 -1054 -522
rect -998 -556 -964 -522
rect -908 -556 -874 -522
rect -818 -556 -784 -522
rect -1358 -646 -1324 -612
rect -1268 -646 -1234 -612
rect -1178 -646 -1144 -612
rect -1088 -646 -1054 -612
rect -998 -646 -964 -612
rect -908 -646 -874 -612
rect -818 -646 -784 -612
rect -1358 -736 -1324 -702
rect -1268 -736 -1234 -702
rect -1178 -736 -1144 -702
rect -1088 -736 -1054 -702
rect -998 -736 -964 -702
rect -908 -736 -874 -702
rect -818 -736 -784 -702
rect 2 -196 36 -162
rect 92 -196 126 -162
rect 182 -196 216 -162
rect 272 -196 306 -162
rect 362 -196 396 -162
rect 452 -196 486 -162
rect 542 -196 576 -162
rect 2 -286 36 -252
rect 92 -286 126 -252
rect 182 -286 216 -252
rect 272 -286 306 -252
rect 362 -286 396 -252
rect 452 -286 486 -252
rect 542 -286 576 -252
rect 2 -376 36 -342
rect 92 -376 126 -342
rect 182 -376 216 -342
rect 272 -376 306 -342
rect 362 -376 396 -342
rect 452 -376 486 -342
rect 542 -376 576 -342
rect 2 -466 36 -432
rect 92 -466 126 -432
rect 182 -466 216 -432
rect 272 -466 306 -432
rect 362 -466 396 -432
rect 452 -466 486 -432
rect 542 -466 576 -432
rect 2 -556 36 -522
rect 92 -556 126 -522
rect 182 -556 216 -522
rect 272 -556 306 -522
rect 362 -556 396 -522
rect 452 -556 486 -522
rect 542 -556 576 -522
rect 2 -646 36 -612
rect 92 -646 126 -612
rect 182 -646 216 -612
rect 272 -646 306 -612
rect 362 -646 396 -612
rect 452 -646 486 -612
rect 542 -646 576 -612
rect 2 -736 36 -702
rect 92 -736 126 -702
rect 182 -736 216 -702
rect 272 -736 306 -702
rect 362 -736 396 -702
rect 452 -736 486 -702
rect 542 -736 576 -702
rect 1362 -196 1396 -162
rect 1452 -196 1486 -162
rect 1542 -196 1576 -162
rect 1632 -196 1666 -162
rect 1722 -196 1756 -162
rect 1812 -196 1846 -162
rect 1902 -196 1936 -162
rect 1362 -286 1396 -252
rect 1452 -286 1486 -252
rect 1542 -286 1576 -252
rect 1632 -286 1666 -252
rect 1722 -286 1756 -252
rect 1812 -286 1846 -252
rect 1902 -286 1936 -252
rect 1362 -376 1396 -342
rect 1452 -376 1486 -342
rect 1542 -376 1576 -342
rect 1632 -376 1666 -342
rect 1722 -376 1756 -342
rect 1812 -376 1846 -342
rect 1902 -376 1936 -342
rect 1362 -466 1396 -432
rect 1452 -466 1486 -432
rect 1542 -466 1576 -432
rect 1632 -466 1666 -432
rect 1722 -466 1756 -432
rect 1812 -466 1846 -432
rect 1902 -466 1936 -432
rect 1362 -556 1396 -522
rect 1452 -556 1486 -522
rect 1542 -556 1576 -522
rect 1632 -556 1666 -522
rect 1722 -556 1756 -522
rect 1812 -556 1846 -522
rect 1902 -556 1936 -522
rect 1362 -646 1396 -612
rect 1452 -646 1486 -612
rect 1542 -646 1576 -612
rect 1632 -646 1666 -612
rect 1722 -646 1756 -612
rect 1812 -646 1846 -612
rect 1902 -646 1936 -612
rect 1362 -736 1396 -702
rect 1452 -736 1486 -702
rect 1542 -736 1576 -702
rect 1632 -736 1666 -702
rect 1722 -736 1756 -702
rect 1812 -736 1846 -702
rect 1902 -736 1936 -702
rect -1358 -1556 -1324 -1522
rect -1268 -1556 -1234 -1522
rect -1178 -1556 -1144 -1522
rect -1088 -1556 -1054 -1522
rect -998 -1556 -964 -1522
rect -908 -1556 -874 -1522
rect -818 -1556 -784 -1522
rect -1358 -1646 -1324 -1612
rect -1268 -1646 -1234 -1612
rect -1178 -1646 -1144 -1612
rect -1088 -1646 -1054 -1612
rect -998 -1646 -964 -1612
rect -908 -1646 -874 -1612
rect -818 -1646 -784 -1612
rect -1358 -1736 -1324 -1702
rect -1268 -1736 -1234 -1702
rect -1178 -1736 -1144 -1702
rect -1088 -1736 -1054 -1702
rect -998 -1736 -964 -1702
rect -908 -1736 -874 -1702
rect -818 -1736 -784 -1702
rect -1358 -1826 -1324 -1792
rect -1268 -1826 -1234 -1792
rect -1178 -1826 -1144 -1792
rect -1088 -1826 -1054 -1792
rect -998 -1826 -964 -1792
rect -908 -1826 -874 -1792
rect -818 -1826 -784 -1792
rect -1358 -1916 -1324 -1882
rect -1268 -1916 -1234 -1882
rect -1178 -1916 -1144 -1882
rect -1088 -1916 -1054 -1882
rect -998 -1916 -964 -1882
rect -908 -1916 -874 -1882
rect -818 -1916 -784 -1882
rect -1358 -2006 -1324 -1972
rect -1268 -2006 -1234 -1972
rect -1178 -2006 -1144 -1972
rect -1088 -2006 -1054 -1972
rect -998 -2006 -964 -1972
rect -908 -2006 -874 -1972
rect -818 -2006 -784 -1972
rect -1358 -2096 -1324 -2062
rect -1268 -2096 -1234 -2062
rect -1178 -2096 -1144 -2062
rect -1088 -2096 -1054 -2062
rect -998 -2096 -964 -2062
rect -908 -2096 -874 -2062
rect -818 -2096 -784 -2062
rect 2 -1556 36 -1522
rect 92 -1556 126 -1522
rect 182 -1556 216 -1522
rect 272 -1556 306 -1522
rect 362 -1556 396 -1522
rect 452 -1556 486 -1522
rect 542 -1556 576 -1522
rect 2 -1646 36 -1612
rect 92 -1646 126 -1612
rect 182 -1646 216 -1612
rect 272 -1646 306 -1612
rect 362 -1646 396 -1612
rect 452 -1646 486 -1612
rect 542 -1646 576 -1612
rect 2 -1736 36 -1702
rect 92 -1736 126 -1702
rect 182 -1736 216 -1702
rect 272 -1736 306 -1702
rect 362 -1736 396 -1702
rect 452 -1736 486 -1702
rect 542 -1736 576 -1702
rect 2 -1826 36 -1792
rect 92 -1826 126 -1792
rect 182 -1826 216 -1792
rect 272 -1826 306 -1792
rect 362 -1826 396 -1792
rect 452 -1826 486 -1792
rect 542 -1826 576 -1792
rect 2 -1916 36 -1882
rect 92 -1916 126 -1882
rect 182 -1916 216 -1882
rect 272 -1916 306 -1882
rect 362 -1916 396 -1882
rect 452 -1916 486 -1882
rect 542 -1916 576 -1882
rect 2 -2006 36 -1972
rect 92 -2006 126 -1972
rect 182 -2006 216 -1972
rect 272 -2006 306 -1972
rect 362 -2006 396 -1972
rect 452 -2006 486 -1972
rect 542 -2006 576 -1972
rect 2 -2096 36 -2062
rect 92 -2096 126 -2062
rect 182 -2096 216 -2062
rect 272 -2096 306 -2062
rect 362 -2096 396 -2062
rect 452 -2096 486 -2062
rect 542 -2096 576 -2062
rect 1362 -1556 1396 -1522
rect 1452 -1556 1486 -1522
rect 1542 -1556 1576 -1522
rect 1632 -1556 1666 -1522
rect 1722 -1556 1756 -1522
rect 1812 -1556 1846 -1522
rect 1902 -1556 1936 -1522
rect 1362 -1646 1396 -1612
rect 1452 -1646 1486 -1612
rect 1542 -1646 1576 -1612
rect 1632 -1646 1666 -1612
rect 1722 -1646 1756 -1612
rect 1812 -1646 1846 -1612
rect 1902 -1646 1936 -1612
rect 1362 -1736 1396 -1702
rect 1452 -1736 1486 -1702
rect 1542 -1736 1576 -1702
rect 1632 -1736 1666 -1702
rect 1722 -1736 1756 -1702
rect 1812 -1736 1846 -1702
rect 1902 -1736 1936 -1702
rect 1362 -1826 1396 -1792
rect 1452 -1826 1486 -1792
rect 1542 -1826 1576 -1792
rect 1632 -1826 1666 -1792
rect 1722 -1826 1756 -1792
rect 1812 -1826 1846 -1792
rect 1902 -1826 1936 -1792
rect 1362 -1916 1396 -1882
rect 1452 -1916 1486 -1882
rect 1542 -1916 1576 -1882
rect 1632 -1916 1666 -1882
rect 1722 -1916 1756 -1882
rect 1812 -1916 1846 -1882
rect 1902 -1916 1936 -1882
rect 1362 -2006 1396 -1972
rect 1452 -2006 1486 -1972
rect 1542 -2006 1576 -1972
rect 1632 -2006 1666 -1972
rect 1722 -2006 1756 -1972
rect 1812 -2006 1846 -1972
rect 1902 -2006 1936 -1972
rect 1362 -2096 1396 -2062
rect 1452 -2096 1486 -2062
rect 1542 -2096 1576 -2062
rect 1632 -2096 1666 -2062
rect 1722 -2096 1756 -2062
rect 1812 -2096 1846 -2062
rect 1902 -2096 1936 -2062
<< psubdiff >>
rect 9200 13850 10330 13890
rect 10470 13850 11230 13890
rect 9200 13470 9240 13850
rect 11190 13470 11230 13850
rect 5030 12900 5110 12930
rect 5030 12860 5050 12900
rect 5090 12860 5110 12900
rect 1790 12810 1870 12840
rect 1790 12770 1810 12810
rect 1850 12770 1870 12810
rect 1790 12740 1870 12770
rect 3240 12810 3320 12840
rect 3240 12770 3260 12810
rect 3300 12770 3320 12810
rect 3240 12740 3320 12770
rect 5030 12830 5110 12860
rect 6330 12900 6410 12930
rect 6330 12860 6350 12900
rect 6390 12860 6410 12900
rect 6330 12830 6410 12860
rect 7630 12900 7710 12930
rect 7630 12860 7650 12900
rect 7690 12860 7710 12900
rect 7630 12830 7710 12860
rect 9200 12770 9240 13210
rect 11190 12770 11230 13210
rect 9200 12730 10330 12770
rect 10470 12730 11230 12770
rect -720 10210 -640 10240
rect -720 10170 -700 10210
rect -660 10170 -640 10210
rect -720 10110 -640 10170
rect -720 10070 -700 10110
rect -660 10070 -640 10110
rect -720 10040 -640 10070
rect 180 10210 260 10240
rect 180 10170 200 10210
rect 240 10170 260 10210
rect 180 10110 260 10170
rect 180 10070 200 10110
rect 240 10070 260 10110
rect 180 10040 260 10070
rect 1080 10210 1160 10240
rect 1080 10170 1100 10210
rect 1140 10170 1160 10210
rect 1080 10110 1160 10170
rect 1080 10070 1100 10110
rect 1140 10070 1160 10110
rect 1080 10040 1160 10070
rect 1220 10210 1300 10240
rect 1220 10170 1240 10210
rect 1280 10170 1300 10210
rect 1220 10110 1300 10170
rect 1220 10070 1240 10110
rect 1280 10070 1300 10110
rect 1220 10040 1300 10070
rect 1660 10210 1740 10240
rect 1660 10170 1680 10210
rect 1720 10170 1740 10210
rect 1660 10110 1740 10170
rect 1660 10070 1680 10110
rect 1720 10070 1740 10110
rect 1660 10040 1740 10070
rect 1990 10210 2070 10240
rect 1990 10170 2010 10210
rect 2050 10170 2070 10210
rect 1990 10110 2070 10170
rect 1990 10070 2010 10110
rect 2050 10070 2070 10110
rect 1990 10040 2070 10070
rect 2410 10210 2490 10240
rect 2410 10170 2430 10210
rect 2470 10170 2490 10210
rect 2410 10110 2490 10170
rect 2410 10070 2430 10110
rect 2470 10070 2490 10110
rect 2410 10040 2490 10070
rect 2800 10210 2880 10240
rect 2800 10170 2820 10210
rect 2860 10170 2880 10210
rect 2800 10110 2880 10170
rect 2800 10070 2820 10110
rect 2860 10070 2880 10110
rect 2800 10040 2880 10070
rect 3190 10210 3270 10240
rect 3190 10170 3210 10210
rect 3250 10170 3270 10210
rect 3190 10110 3270 10170
rect 3190 10070 3210 10110
rect 3250 10070 3270 10110
rect 3190 10040 3270 10070
rect 5340 8660 5440 8690
rect 5340 8620 5370 8660
rect 5410 8620 5440 8660
rect 5340 8560 5440 8620
rect 5340 8520 5370 8560
rect 5410 8520 5440 8560
rect 5340 8460 5440 8520
rect -720 8410 -640 8440
rect -720 8370 -700 8410
rect -660 8370 -640 8410
rect -720 8310 -640 8370
rect -720 8270 -700 8310
rect -660 8270 -640 8310
rect -720 8240 -640 8270
rect 180 8410 260 8440
rect 180 8370 200 8410
rect 240 8370 260 8410
rect 180 8310 260 8370
rect 180 8270 200 8310
rect 240 8270 260 8310
rect 180 8240 260 8270
rect 1080 8410 1160 8440
rect 1080 8370 1100 8410
rect 1140 8370 1160 8410
rect 1080 8310 1160 8370
rect 1080 8270 1100 8310
rect 1140 8270 1160 8310
rect 1080 8240 1160 8270
rect 1480 8410 1560 8440
rect 1480 8370 1500 8410
rect 1540 8370 1560 8410
rect 1480 8310 1560 8370
rect 1480 8270 1500 8310
rect 1540 8270 1560 8310
rect 1480 8240 1560 8270
rect 1810 8410 1890 8440
rect 1810 8370 1830 8410
rect 1870 8370 1890 8410
rect 1810 8310 1890 8370
rect 1810 8270 1830 8310
rect 1870 8270 1890 8310
rect 1810 8240 1890 8270
rect 2140 8410 2220 8440
rect 2140 8370 2160 8410
rect 2200 8370 2220 8410
rect 2140 8310 2220 8370
rect 2140 8270 2160 8310
rect 2200 8270 2220 8310
rect 2140 8240 2220 8270
rect 2390 8410 2490 8440
rect 2390 8370 2420 8410
rect 2460 8370 2490 8410
rect 2390 8310 2490 8370
rect 2390 8270 2420 8310
rect 2460 8270 2490 8310
rect 2390 8240 2490 8270
rect 3170 8410 3270 8440
rect 3170 8370 3200 8410
rect 3240 8370 3270 8410
rect 3170 8310 3270 8370
rect 3170 8270 3200 8310
rect 3240 8270 3270 8310
rect 3170 8240 3270 8270
rect 3850 8410 3950 8440
rect 3850 8370 3880 8410
rect 3920 8370 3950 8410
rect 3850 8310 3950 8370
rect 3850 8270 3880 8310
rect 3920 8270 3950 8310
rect 3850 8240 3950 8270
rect 5340 8420 5370 8460
rect 5410 8420 5440 8460
rect 5340 8360 5440 8420
rect 5340 8320 5370 8360
rect 5410 8320 5440 8360
rect 5340 8290 5440 8320
rect 6420 8660 6520 8690
rect 6420 8620 6450 8660
rect 6490 8620 6520 8660
rect 6420 8560 6520 8620
rect 6420 8520 6450 8560
rect 6490 8520 6520 8560
rect 6420 8460 6520 8520
rect 6420 8420 6450 8460
rect 6490 8420 6520 8460
rect 6420 8360 6520 8420
rect 6420 8320 6450 8360
rect 6490 8320 6520 8360
rect 6420 8290 6520 8320
rect 7500 8660 7600 8690
rect 7500 8620 7530 8660
rect 7570 8620 7600 8660
rect 7500 8560 7600 8620
rect 7500 8520 7530 8560
rect 7570 8520 7600 8560
rect 7500 8460 7600 8520
rect 7500 8420 7530 8460
rect 7570 8420 7600 8460
rect 7500 8360 7600 8420
rect 7500 8320 7530 8360
rect 7570 8320 7600 8360
rect 7500 8290 7600 8320
rect 8580 8660 8680 8690
rect 8580 8620 8610 8660
rect 8650 8620 8680 8660
rect 8580 8560 8680 8620
rect 8580 8520 8610 8560
rect 8650 8520 8680 8560
rect 8580 8460 8680 8520
rect 8580 8420 8610 8460
rect 8650 8420 8680 8460
rect 8580 8360 8680 8420
rect 8580 8320 8610 8360
rect 8650 8320 8680 8360
rect 8580 8290 8680 8320
rect 5400 6030 5500 6060
rect 5400 5980 5430 6030
rect 5470 5980 5500 6030
rect 5400 5890 5500 5980
rect 5400 5840 5430 5890
rect 5470 5840 5500 5890
rect 5400 5810 5500 5840
rect 7600 6030 7700 6060
rect 7600 5980 7630 6030
rect 7670 5980 7700 6030
rect 7600 5890 7700 5980
rect 7600 5840 7630 5890
rect 7670 5840 7700 5890
rect 7600 5810 7700 5840
rect 5450 5340 5550 5370
rect 5450 5300 5480 5340
rect 5520 5300 5550 5340
rect 5450 5270 5550 5300
rect 6430 5340 6530 5370
rect 6430 5300 6460 5340
rect 6500 5300 6530 5340
rect 6430 5270 6530 5300
rect 7730 5340 7830 5370
rect 7730 5300 7760 5340
rect 7800 5300 7830 5340
rect 7730 5270 7830 5300
rect 8710 5340 8810 5370
rect 8710 5300 8740 5340
rect 8780 5300 8810 5340
rect 8710 5270 8810 5300
rect -190 3810 -110 3840
rect -190 3770 -170 3810
rect -130 3770 -110 3810
rect -190 3730 -110 3770
rect -190 3690 -170 3730
rect -130 3690 -110 3730
rect -190 3650 -110 3690
rect -190 3610 -170 3650
rect -130 3610 -110 3650
rect -190 3580 -110 3610
rect 690 3810 770 3840
rect 690 3770 710 3810
rect 750 3770 770 3810
rect 690 3730 770 3770
rect 690 3690 710 3730
rect 750 3690 770 3730
rect 690 3650 770 3690
rect 690 3610 710 3650
rect 750 3610 770 3650
rect 690 3580 770 3610
rect -1090 3130 -1010 3160
rect -1090 3090 -1070 3130
rect -1030 3090 -1010 3130
rect -1090 3030 -1010 3090
rect -1090 2990 -1070 3030
rect -1030 2990 -1010 3030
rect -1090 2930 -1010 2990
rect -1090 2890 -1070 2930
rect -1030 2890 -1010 2930
rect -1090 2830 -1010 2890
rect -1090 2790 -1070 2830
rect -1030 2790 -1010 2830
rect -1090 2730 -1010 2790
rect -1090 2690 -1070 2730
rect -1030 2690 -1010 2730
rect -1090 2660 -1010 2690
rect 1590 3130 1670 3160
rect 1590 3090 1610 3130
rect 1650 3090 1670 3130
rect 1590 3030 1670 3090
rect 1590 2990 1610 3030
rect 1650 2990 1670 3030
rect 1590 2930 1670 2990
rect 1590 2890 1610 2930
rect 1650 2890 1670 2930
rect 1590 2830 1670 2890
rect 1590 2790 1610 2830
rect 1650 2790 1670 2830
rect 1590 2730 1670 2790
rect 1590 2690 1610 2730
rect 1650 2690 1670 2730
rect 1590 2670 1670 2690
rect 2410 2220 2490 2250
rect 2410 2180 2430 2220
rect 2470 2180 2490 2220
rect 2410 2120 2490 2180
rect 2410 2080 2430 2120
rect 2470 2080 2490 2120
rect 2410 2050 2490 2080
rect -1714 1519 -426 1554
rect -1714 1496 -1580 1519
rect -1714 1462 -1681 1496
rect -1647 1485 -1580 1496
rect -1546 1485 -1490 1519
rect -1456 1485 -1400 1519
rect -1366 1485 -1310 1519
rect -1276 1485 -1220 1519
rect -1186 1485 -1130 1519
rect -1096 1485 -1040 1519
rect -1006 1485 -950 1519
rect -916 1485 -860 1519
rect -826 1485 -770 1519
rect -736 1485 -680 1519
rect -646 1485 -590 1519
rect -556 1496 -426 1519
rect -556 1485 -494 1496
rect -1647 1462 -494 1485
rect -460 1462 -426 1496
rect -1714 1453 -426 1462
rect -1714 1406 -1613 1453
rect -1714 1372 -1681 1406
rect -1647 1372 -1613 1406
rect -527 1406 -426 1453
rect -1714 1316 -1613 1372
rect -1714 1282 -1681 1316
rect -1647 1282 -1613 1316
rect -1714 1226 -1613 1282
rect -1714 1192 -1681 1226
rect -1647 1192 -1613 1226
rect -1714 1136 -1613 1192
rect -1714 1102 -1681 1136
rect -1647 1102 -1613 1136
rect -1714 1046 -1613 1102
rect -1714 1012 -1681 1046
rect -1647 1012 -1613 1046
rect -1714 956 -1613 1012
rect -1714 922 -1681 956
rect -1647 922 -1613 956
rect -1714 866 -1613 922
rect -1714 832 -1681 866
rect -1647 832 -1613 866
rect -1714 776 -1613 832
rect -1714 742 -1681 776
rect -1647 742 -1613 776
rect -1714 686 -1613 742
rect -1714 652 -1681 686
rect -1647 652 -1613 686
rect -1714 596 -1613 652
rect -1714 562 -1681 596
rect -1647 562 -1613 596
rect -1714 506 -1613 562
rect -1714 472 -1681 506
rect -1647 472 -1613 506
rect -1714 416 -1613 472
rect -527 1372 -494 1406
rect -460 1372 -426 1406
rect -527 1316 -426 1372
rect -527 1282 -494 1316
rect -460 1282 -426 1316
rect -527 1226 -426 1282
rect -527 1192 -494 1226
rect -460 1192 -426 1226
rect -527 1136 -426 1192
rect -527 1102 -494 1136
rect -460 1102 -426 1136
rect -527 1046 -426 1102
rect -527 1012 -494 1046
rect -460 1012 -426 1046
rect -527 956 -426 1012
rect -527 922 -494 956
rect -460 922 -426 956
rect -527 866 -426 922
rect -527 832 -494 866
rect -460 832 -426 866
rect -527 776 -426 832
rect -527 742 -494 776
rect -460 742 -426 776
rect -527 686 -426 742
rect -527 652 -494 686
rect -460 652 -426 686
rect -527 596 -426 652
rect -527 562 -494 596
rect -460 562 -426 596
rect -527 506 -426 562
rect -527 472 -494 506
rect -460 472 -426 506
rect -1714 382 -1681 416
rect -1647 382 -1613 416
rect -1714 367 -1613 382
rect -527 416 -426 472
rect -527 382 -494 416
rect -460 382 -426 416
rect -527 367 -426 382
rect -1714 332 -426 367
rect -1714 298 -1580 332
rect -1546 298 -1490 332
rect -1456 298 -1400 332
rect -1366 298 -1310 332
rect -1276 298 -1220 332
rect -1186 298 -1130 332
rect -1096 298 -1040 332
rect -1006 298 -950 332
rect -916 298 -860 332
rect -826 298 -770 332
rect -736 298 -680 332
rect -646 298 -590 332
rect -556 298 -426 332
rect -1714 266 -426 298
rect -354 1519 934 1554
rect -354 1496 -220 1519
rect -354 1462 -321 1496
rect -287 1485 -220 1496
rect -186 1485 -130 1519
rect -96 1485 -40 1519
rect -6 1485 50 1519
rect 84 1485 140 1519
rect 174 1485 230 1519
rect 264 1485 320 1519
rect 354 1485 410 1519
rect 444 1485 500 1519
rect 534 1485 590 1519
rect 624 1485 680 1519
rect 714 1485 770 1519
rect 804 1496 934 1519
rect 804 1485 866 1496
rect -287 1462 866 1485
rect 900 1462 934 1496
rect -354 1453 934 1462
rect -354 1406 -253 1453
rect -354 1372 -321 1406
rect -287 1372 -253 1406
rect 833 1406 934 1453
rect -354 1316 -253 1372
rect -354 1282 -321 1316
rect -287 1282 -253 1316
rect -354 1226 -253 1282
rect -354 1192 -321 1226
rect -287 1192 -253 1226
rect -354 1136 -253 1192
rect -354 1102 -321 1136
rect -287 1102 -253 1136
rect -354 1046 -253 1102
rect -354 1012 -321 1046
rect -287 1012 -253 1046
rect -354 956 -253 1012
rect -354 922 -321 956
rect -287 922 -253 956
rect -354 866 -253 922
rect -354 832 -321 866
rect -287 832 -253 866
rect -354 776 -253 832
rect -354 742 -321 776
rect -287 742 -253 776
rect -354 686 -253 742
rect -354 652 -321 686
rect -287 652 -253 686
rect -354 596 -253 652
rect -354 562 -321 596
rect -287 562 -253 596
rect -354 506 -253 562
rect -354 472 -321 506
rect -287 472 -253 506
rect -354 416 -253 472
rect 833 1372 866 1406
rect 900 1372 934 1406
rect 833 1316 934 1372
rect 833 1282 866 1316
rect 900 1282 934 1316
rect 833 1226 934 1282
rect 833 1192 866 1226
rect 900 1192 934 1226
rect 833 1136 934 1192
rect 833 1102 866 1136
rect 900 1102 934 1136
rect 833 1046 934 1102
rect 833 1012 866 1046
rect 900 1012 934 1046
rect 833 956 934 1012
rect 833 922 866 956
rect 900 922 934 956
rect 833 866 934 922
rect 833 832 866 866
rect 900 832 934 866
rect 833 776 934 832
rect 833 742 866 776
rect 900 742 934 776
rect 833 686 934 742
rect 833 652 866 686
rect 900 652 934 686
rect 833 596 934 652
rect 833 562 866 596
rect 900 562 934 596
rect 833 506 934 562
rect 833 472 866 506
rect 900 472 934 506
rect -354 382 -321 416
rect -287 382 -253 416
rect -354 367 -253 382
rect 833 416 934 472
rect 833 382 866 416
rect 900 382 934 416
rect 833 367 934 382
rect -354 332 934 367
rect -354 298 -220 332
rect -186 298 -130 332
rect -96 298 -40 332
rect -6 298 50 332
rect 84 298 140 332
rect 174 298 230 332
rect 264 298 320 332
rect 354 298 410 332
rect 444 298 500 332
rect 534 298 590 332
rect 624 298 680 332
rect 714 298 770 332
rect 804 298 934 332
rect -354 266 934 298
rect 1006 1519 2294 1554
rect 1006 1496 1140 1519
rect 1006 1462 1039 1496
rect 1073 1485 1140 1496
rect 1174 1485 1230 1519
rect 1264 1485 1320 1519
rect 1354 1485 1410 1519
rect 1444 1485 1500 1519
rect 1534 1485 1590 1519
rect 1624 1485 1680 1519
rect 1714 1485 1770 1519
rect 1804 1485 1860 1519
rect 1894 1485 1950 1519
rect 1984 1485 2040 1519
rect 2074 1485 2130 1519
rect 2164 1496 2294 1519
rect 2164 1485 2226 1496
rect 1073 1462 2226 1485
rect 2260 1462 2294 1496
rect 1006 1453 2294 1462
rect 1006 1406 1107 1453
rect 1006 1372 1039 1406
rect 1073 1372 1107 1406
rect 2193 1406 2294 1453
rect 1006 1316 1107 1372
rect 1006 1282 1039 1316
rect 1073 1282 1107 1316
rect 1006 1226 1107 1282
rect 1006 1192 1039 1226
rect 1073 1192 1107 1226
rect 1006 1136 1107 1192
rect 1006 1102 1039 1136
rect 1073 1102 1107 1136
rect 1006 1046 1107 1102
rect 1006 1012 1039 1046
rect 1073 1012 1107 1046
rect 1006 956 1107 1012
rect 1006 922 1039 956
rect 1073 922 1107 956
rect 1006 866 1107 922
rect 1006 832 1039 866
rect 1073 832 1107 866
rect 1006 776 1107 832
rect 1006 742 1039 776
rect 1073 742 1107 776
rect 1006 686 1107 742
rect 1006 652 1039 686
rect 1073 652 1107 686
rect 1006 596 1107 652
rect 1006 562 1039 596
rect 1073 562 1107 596
rect 1006 506 1107 562
rect 1006 472 1039 506
rect 1073 472 1107 506
rect 1006 416 1107 472
rect 2193 1372 2226 1406
rect 2260 1372 2294 1406
rect 2193 1316 2294 1372
rect 2193 1282 2226 1316
rect 2260 1282 2294 1316
rect 2193 1226 2294 1282
rect 2193 1192 2226 1226
rect 2260 1192 2294 1226
rect 2193 1136 2294 1192
rect 2193 1102 2226 1136
rect 2260 1102 2294 1136
rect 2193 1046 2294 1102
rect 2193 1012 2226 1046
rect 2260 1012 2294 1046
rect 2193 956 2294 1012
rect 2193 922 2226 956
rect 2260 922 2294 956
rect 2193 866 2294 922
rect 2193 832 2226 866
rect 2260 832 2294 866
rect 2193 776 2294 832
rect 2193 742 2226 776
rect 2260 742 2294 776
rect 2193 686 2294 742
rect 2193 652 2226 686
rect 2260 652 2294 686
rect 2193 596 2294 652
rect 2193 562 2226 596
rect 2260 562 2294 596
rect 2193 506 2294 562
rect 2193 472 2226 506
rect 2260 472 2294 506
rect 1006 382 1039 416
rect 1073 382 1107 416
rect 1006 367 1107 382
rect 2193 416 2294 472
rect 2193 382 2226 416
rect 2260 382 2294 416
rect 2193 367 2294 382
rect 1006 332 2294 367
rect 1006 298 1140 332
rect 1174 298 1230 332
rect 1264 298 1320 332
rect 1354 298 1410 332
rect 1444 298 1500 332
rect 1534 298 1590 332
rect 1624 298 1680 332
rect 1714 298 1770 332
rect 1804 298 1860 332
rect 1894 298 1950 332
rect 1984 298 2040 332
rect 2074 298 2130 332
rect 2164 298 2294 332
rect 1006 266 2294 298
rect -1714 159 -426 194
rect -1714 136 -1580 159
rect -1714 102 -1681 136
rect -1647 125 -1580 136
rect -1546 125 -1490 159
rect -1456 125 -1400 159
rect -1366 125 -1310 159
rect -1276 125 -1220 159
rect -1186 125 -1130 159
rect -1096 125 -1040 159
rect -1006 125 -950 159
rect -916 125 -860 159
rect -826 125 -770 159
rect -736 125 -680 159
rect -646 125 -590 159
rect -556 136 -426 159
rect -556 125 -494 136
rect -1647 102 -494 125
rect -460 102 -426 136
rect -1714 93 -426 102
rect -1714 46 -1613 93
rect -1714 12 -1681 46
rect -1647 12 -1613 46
rect -527 46 -426 93
rect -1714 -44 -1613 12
rect -1714 -78 -1681 -44
rect -1647 -78 -1613 -44
rect -3040 -1390 -2960 -1360
rect -3040 -1430 -3020 -1390
rect -2980 -1430 -2960 -1390
rect -3040 -1460 -2960 -1430
rect -1714 -134 -1613 -78
rect -1714 -168 -1681 -134
rect -1647 -168 -1613 -134
rect -1714 -224 -1613 -168
rect -1714 -258 -1681 -224
rect -1647 -258 -1613 -224
rect -1714 -314 -1613 -258
rect -1714 -348 -1681 -314
rect -1647 -348 -1613 -314
rect -1714 -404 -1613 -348
rect -1714 -438 -1681 -404
rect -1647 -438 -1613 -404
rect -1714 -494 -1613 -438
rect -1714 -528 -1681 -494
rect -1647 -528 -1613 -494
rect -1714 -584 -1613 -528
rect -1714 -618 -1681 -584
rect -1647 -618 -1613 -584
rect -1714 -674 -1613 -618
rect -1714 -708 -1681 -674
rect -1647 -708 -1613 -674
rect -1714 -764 -1613 -708
rect -1714 -798 -1681 -764
rect -1647 -798 -1613 -764
rect -1714 -854 -1613 -798
rect -1714 -888 -1681 -854
rect -1647 -888 -1613 -854
rect -1714 -944 -1613 -888
rect -527 12 -494 46
rect -460 12 -426 46
rect -527 -44 -426 12
rect -527 -78 -494 -44
rect -460 -78 -426 -44
rect -527 -134 -426 -78
rect -527 -168 -494 -134
rect -460 -168 -426 -134
rect -527 -224 -426 -168
rect -527 -258 -494 -224
rect -460 -258 -426 -224
rect -527 -314 -426 -258
rect -527 -348 -494 -314
rect -460 -348 -426 -314
rect -527 -404 -426 -348
rect -527 -438 -494 -404
rect -460 -438 -426 -404
rect -527 -494 -426 -438
rect -527 -528 -494 -494
rect -460 -528 -426 -494
rect -527 -584 -426 -528
rect -527 -618 -494 -584
rect -460 -618 -426 -584
rect -527 -674 -426 -618
rect -527 -708 -494 -674
rect -460 -708 -426 -674
rect -527 -764 -426 -708
rect -527 -798 -494 -764
rect -460 -798 -426 -764
rect -527 -854 -426 -798
rect -527 -888 -494 -854
rect -460 -888 -426 -854
rect -1714 -978 -1681 -944
rect -1647 -978 -1613 -944
rect -1714 -993 -1613 -978
rect -527 -944 -426 -888
rect -527 -978 -494 -944
rect -460 -978 -426 -944
rect -527 -993 -426 -978
rect -1714 -1028 -426 -993
rect -1714 -1062 -1580 -1028
rect -1546 -1062 -1490 -1028
rect -1456 -1062 -1400 -1028
rect -1366 -1062 -1310 -1028
rect -1276 -1062 -1220 -1028
rect -1186 -1062 -1130 -1028
rect -1096 -1062 -1040 -1028
rect -1006 -1062 -950 -1028
rect -916 -1062 -860 -1028
rect -826 -1062 -770 -1028
rect -736 -1062 -680 -1028
rect -646 -1062 -590 -1028
rect -556 -1062 -426 -1028
rect -1714 -1094 -426 -1062
rect -354 159 934 194
rect -354 136 -220 159
rect -354 102 -321 136
rect -287 125 -220 136
rect -186 125 -130 159
rect -96 125 -40 159
rect -6 125 50 159
rect 84 125 140 159
rect 174 125 230 159
rect 264 125 320 159
rect 354 125 410 159
rect 444 125 500 159
rect 534 125 590 159
rect 624 125 680 159
rect 714 125 770 159
rect 804 136 934 159
rect 804 125 866 136
rect -287 102 866 125
rect 900 102 934 136
rect -354 93 934 102
rect -354 46 -253 93
rect -354 12 -321 46
rect -287 12 -253 46
rect 833 46 934 93
rect -354 -44 -253 12
rect -354 -78 -321 -44
rect -287 -78 -253 -44
rect -354 -134 -253 -78
rect -354 -168 -321 -134
rect -287 -168 -253 -134
rect -354 -224 -253 -168
rect -354 -258 -321 -224
rect -287 -258 -253 -224
rect -354 -314 -253 -258
rect -354 -348 -321 -314
rect -287 -348 -253 -314
rect -354 -404 -253 -348
rect -354 -438 -321 -404
rect -287 -438 -253 -404
rect -354 -494 -253 -438
rect -354 -528 -321 -494
rect -287 -528 -253 -494
rect -354 -584 -253 -528
rect -354 -618 -321 -584
rect -287 -618 -253 -584
rect -354 -674 -253 -618
rect -354 -708 -321 -674
rect -287 -708 -253 -674
rect -354 -764 -253 -708
rect -354 -798 -321 -764
rect -287 -798 -253 -764
rect -354 -854 -253 -798
rect -354 -888 -321 -854
rect -287 -888 -253 -854
rect -354 -944 -253 -888
rect 833 12 866 46
rect 900 12 934 46
rect 833 -44 934 12
rect 833 -78 866 -44
rect 900 -78 934 -44
rect 833 -134 934 -78
rect 833 -168 866 -134
rect 900 -168 934 -134
rect 833 -224 934 -168
rect 833 -258 866 -224
rect 900 -258 934 -224
rect 833 -314 934 -258
rect 833 -348 866 -314
rect 900 -348 934 -314
rect 833 -404 934 -348
rect 833 -438 866 -404
rect 900 -438 934 -404
rect 833 -494 934 -438
rect 833 -528 866 -494
rect 900 -528 934 -494
rect 833 -584 934 -528
rect 833 -618 866 -584
rect 900 -618 934 -584
rect 833 -674 934 -618
rect 833 -708 866 -674
rect 900 -708 934 -674
rect 833 -764 934 -708
rect 833 -798 866 -764
rect 900 -798 934 -764
rect 833 -854 934 -798
rect 833 -888 866 -854
rect 900 -888 934 -854
rect -354 -978 -321 -944
rect -287 -978 -253 -944
rect -354 -993 -253 -978
rect 833 -944 934 -888
rect 833 -978 866 -944
rect 900 -978 934 -944
rect 833 -993 934 -978
rect -354 -1028 934 -993
rect -354 -1062 -220 -1028
rect -186 -1062 -130 -1028
rect -96 -1062 -40 -1028
rect -6 -1062 50 -1028
rect 84 -1062 140 -1028
rect 174 -1062 230 -1028
rect 264 -1062 320 -1028
rect 354 -1062 410 -1028
rect 444 -1062 500 -1028
rect 534 -1062 590 -1028
rect 624 -1062 680 -1028
rect 714 -1062 770 -1028
rect 804 -1062 934 -1028
rect -354 -1094 934 -1062
rect 1006 159 2294 194
rect 1006 136 1140 159
rect 1006 102 1039 136
rect 1073 125 1140 136
rect 1174 125 1230 159
rect 1264 125 1320 159
rect 1354 125 1410 159
rect 1444 125 1500 159
rect 1534 125 1590 159
rect 1624 125 1680 159
rect 1714 125 1770 159
rect 1804 125 1860 159
rect 1894 125 1950 159
rect 1984 125 2040 159
rect 2074 125 2130 159
rect 2164 136 2294 159
rect 2164 125 2226 136
rect 1073 102 2226 125
rect 2260 102 2294 136
rect 1006 93 2294 102
rect 1006 46 1107 93
rect 1006 12 1039 46
rect 1073 12 1107 46
rect 2193 46 2294 93
rect 1006 -44 1107 12
rect 1006 -78 1039 -44
rect 1073 -78 1107 -44
rect 1006 -134 1107 -78
rect 1006 -168 1039 -134
rect 1073 -168 1107 -134
rect 1006 -224 1107 -168
rect 1006 -258 1039 -224
rect 1073 -258 1107 -224
rect 1006 -314 1107 -258
rect 1006 -348 1039 -314
rect 1073 -348 1107 -314
rect 1006 -404 1107 -348
rect 1006 -438 1039 -404
rect 1073 -438 1107 -404
rect 1006 -494 1107 -438
rect 1006 -528 1039 -494
rect 1073 -528 1107 -494
rect 1006 -584 1107 -528
rect 1006 -618 1039 -584
rect 1073 -618 1107 -584
rect 1006 -674 1107 -618
rect 1006 -708 1039 -674
rect 1073 -708 1107 -674
rect 1006 -764 1107 -708
rect 1006 -798 1039 -764
rect 1073 -798 1107 -764
rect 1006 -854 1107 -798
rect 1006 -888 1039 -854
rect 1073 -888 1107 -854
rect 1006 -944 1107 -888
rect 2193 12 2226 46
rect 2260 12 2294 46
rect 2193 -44 2294 12
rect 2193 -78 2226 -44
rect 2260 -78 2294 -44
rect 2193 -134 2294 -78
rect 2193 -168 2226 -134
rect 2260 -168 2294 -134
rect 2193 -224 2294 -168
rect 2193 -258 2226 -224
rect 2260 -258 2294 -224
rect 2193 -314 2294 -258
rect 2193 -348 2226 -314
rect 2260 -348 2294 -314
rect 2193 -404 2294 -348
rect 2193 -438 2226 -404
rect 2260 -438 2294 -404
rect 2193 -494 2294 -438
rect 2193 -528 2226 -494
rect 2260 -528 2294 -494
rect 2193 -584 2294 -528
rect 2193 -618 2226 -584
rect 2260 -618 2294 -584
rect 2193 -674 2294 -618
rect 2193 -708 2226 -674
rect 2260 -708 2294 -674
rect 2193 -764 2294 -708
rect 2193 -798 2226 -764
rect 2260 -798 2294 -764
rect 2193 -854 2294 -798
rect 2193 -888 2226 -854
rect 2260 -888 2294 -854
rect 1006 -978 1039 -944
rect 1073 -978 1107 -944
rect 1006 -993 1107 -978
rect 2193 -944 2294 -888
rect 2193 -978 2226 -944
rect 2260 -978 2294 -944
rect 2193 -993 2294 -978
rect 1006 -1028 2294 -993
rect 1006 -1062 1140 -1028
rect 1174 -1062 1230 -1028
rect 1264 -1062 1320 -1028
rect 1354 -1062 1410 -1028
rect 1444 -1062 1500 -1028
rect 1534 -1062 1590 -1028
rect 1624 -1062 1680 -1028
rect 1714 -1062 1770 -1028
rect 1804 -1062 1860 -1028
rect 1894 -1062 1950 -1028
rect 1984 -1062 2040 -1028
rect 2074 -1062 2130 -1028
rect 2164 -1062 2294 -1028
rect 1006 -1094 2294 -1062
rect -1714 -1201 -426 -1166
rect -1714 -1224 -1580 -1201
rect -1714 -1258 -1681 -1224
rect -1647 -1235 -1580 -1224
rect -1546 -1235 -1490 -1201
rect -1456 -1235 -1400 -1201
rect -1366 -1235 -1310 -1201
rect -1276 -1235 -1220 -1201
rect -1186 -1235 -1130 -1201
rect -1096 -1235 -1040 -1201
rect -1006 -1235 -950 -1201
rect -916 -1235 -860 -1201
rect -826 -1235 -770 -1201
rect -736 -1235 -680 -1201
rect -646 -1235 -590 -1201
rect -556 -1224 -426 -1201
rect -556 -1235 -494 -1224
rect -1647 -1258 -494 -1235
rect -460 -1258 -426 -1224
rect -1714 -1267 -426 -1258
rect -1714 -1314 -1613 -1267
rect -1714 -1348 -1681 -1314
rect -1647 -1348 -1613 -1314
rect -527 -1314 -426 -1267
rect -1714 -1404 -1613 -1348
rect -1714 -1438 -1681 -1404
rect -1647 -1438 -1613 -1404
rect -1714 -1494 -1613 -1438
rect -1714 -1528 -1681 -1494
rect -1647 -1528 -1613 -1494
rect -1714 -1584 -1613 -1528
rect -1714 -1618 -1681 -1584
rect -1647 -1618 -1613 -1584
rect -1714 -1674 -1613 -1618
rect -1714 -1708 -1681 -1674
rect -1647 -1708 -1613 -1674
rect -1714 -1764 -1613 -1708
rect -1714 -1798 -1681 -1764
rect -1647 -1798 -1613 -1764
rect -1714 -1854 -1613 -1798
rect -1714 -1888 -1681 -1854
rect -1647 -1888 -1613 -1854
rect -1714 -1944 -1613 -1888
rect -1714 -1978 -1681 -1944
rect -1647 -1978 -1613 -1944
rect -1714 -2034 -1613 -1978
rect -1714 -2068 -1681 -2034
rect -1647 -2068 -1613 -2034
rect -1714 -2124 -1613 -2068
rect -1714 -2158 -1681 -2124
rect -1647 -2158 -1613 -2124
rect -1714 -2214 -1613 -2158
rect -1714 -2248 -1681 -2214
rect -1647 -2248 -1613 -2214
rect -1714 -2304 -1613 -2248
rect -527 -1348 -494 -1314
rect -460 -1348 -426 -1314
rect -527 -1404 -426 -1348
rect -527 -1438 -494 -1404
rect -460 -1438 -426 -1404
rect -527 -1494 -426 -1438
rect -527 -1528 -494 -1494
rect -460 -1528 -426 -1494
rect -527 -1584 -426 -1528
rect -527 -1618 -494 -1584
rect -460 -1618 -426 -1584
rect -527 -1674 -426 -1618
rect -527 -1708 -494 -1674
rect -460 -1708 -426 -1674
rect -527 -1764 -426 -1708
rect -527 -1798 -494 -1764
rect -460 -1798 -426 -1764
rect -527 -1854 -426 -1798
rect -527 -1888 -494 -1854
rect -460 -1888 -426 -1854
rect -527 -1944 -426 -1888
rect -527 -1978 -494 -1944
rect -460 -1978 -426 -1944
rect -527 -2034 -426 -1978
rect -527 -2068 -494 -2034
rect -460 -2068 -426 -2034
rect -527 -2124 -426 -2068
rect -527 -2158 -494 -2124
rect -460 -2158 -426 -2124
rect -527 -2214 -426 -2158
rect -527 -2248 -494 -2214
rect -460 -2248 -426 -2214
rect -1714 -2338 -1681 -2304
rect -1647 -2338 -1613 -2304
rect -1714 -2353 -1613 -2338
rect -527 -2304 -426 -2248
rect -527 -2338 -494 -2304
rect -460 -2338 -426 -2304
rect -527 -2353 -426 -2338
rect -1714 -2388 -426 -2353
rect -1714 -2422 -1580 -2388
rect -1546 -2422 -1490 -2388
rect -1456 -2422 -1400 -2388
rect -1366 -2422 -1310 -2388
rect -1276 -2422 -1220 -2388
rect -1186 -2422 -1130 -2388
rect -1096 -2422 -1040 -2388
rect -1006 -2422 -950 -2388
rect -916 -2422 -860 -2388
rect -826 -2422 -770 -2388
rect -736 -2422 -680 -2388
rect -646 -2422 -590 -2388
rect -556 -2422 -426 -2388
rect -1714 -2454 -426 -2422
rect -354 -1201 934 -1166
rect -354 -1224 -220 -1201
rect -354 -1258 -321 -1224
rect -287 -1235 -220 -1224
rect -186 -1235 -130 -1201
rect -96 -1235 -40 -1201
rect -6 -1235 50 -1201
rect 84 -1235 140 -1201
rect 174 -1235 230 -1201
rect 264 -1235 320 -1201
rect 354 -1235 410 -1201
rect 444 -1235 500 -1201
rect 534 -1235 590 -1201
rect 624 -1235 680 -1201
rect 714 -1235 770 -1201
rect 804 -1224 934 -1201
rect 804 -1235 866 -1224
rect -287 -1258 866 -1235
rect 900 -1258 934 -1224
rect -354 -1267 934 -1258
rect -354 -1314 -253 -1267
rect -354 -1348 -321 -1314
rect -287 -1348 -253 -1314
rect 833 -1314 934 -1267
rect -354 -1404 -253 -1348
rect -354 -1438 -321 -1404
rect -287 -1438 -253 -1404
rect -354 -1494 -253 -1438
rect -354 -1528 -321 -1494
rect -287 -1528 -253 -1494
rect -354 -1584 -253 -1528
rect -354 -1618 -321 -1584
rect -287 -1618 -253 -1584
rect -354 -1674 -253 -1618
rect -354 -1708 -321 -1674
rect -287 -1708 -253 -1674
rect -354 -1764 -253 -1708
rect -354 -1798 -321 -1764
rect -287 -1798 -253 -1764
rect -354 -1854 -253 -1798
rect -354 -1888 -321 -1854
rect -287 -1888 -253 -1854
rect -354 -1944 -253 -1888
rect -354 -1978 -321 -1944
rect -287 -1978 -253 -1944
rect -354 -2034 -253 -1978
rect -354 -2068 -321 -2034
rect -287 -2068 -253 -2034
rect -354 -2124 -253 -2068
rect -354 -2158 -321 -2124
rect -287 -2158 -253 -2124
rect -354 -2214 -253 -2158
rect -354 -2248 -321 -2214
rect -287 -2248 -253 -2214
rect -354 -2304 -253 -2248
rect 833 -1348 866 -1314
rect 900 -1348 934 -1314
rect 833 -1404 934 -1348
rect 833 -1438 866 -1404
rect 900 -1438 934 -1404
rect 833 -1494 934 -1438
rect 833 -1528 866 -1494
rect 900 -1528 934 -1494
rect 833 -1584 934 -1528
rect 833 -1618 866 -1584
rect 900 -1618 934 -1584
rect 833 -1674 934 -1618
rect 833 -1708 866 -1674
rect 900 -1708 934 -1674
rect 833 -1764 934 -1708
rect 833 -1798 866 -1764
rect 900 -1798 934 -1764
rect 833 -1854 934 -1798
rect 833 -1888 866 -1854
rect 900 -1888 934 -1854
rect 833 -1944 934 -1888
rect 833 -1978 866 -1944
rect 900 -1978 934 -1944
rect 833 -2034 934 -1978
rect 833 -2068 866 -2034
rect 900 -2068 934 -2034
rect 833 -2124 934 -2068
rect 833 -2158 866 -2124
rect 900 -2158 934 -2124
rect 833 -2214 934 -2158
rect 833 -2248 866 -2214
rect 900 -2248 934 -2214
rect -354 -2338 -321 -2304
rect -287 -2338 -253 -2304
rect -354 -2353 -253 -2338
rect 833 -2304 934 -2248
rect 833 -2338 866 -2304
rect 900 -2338 934 -2304
rect 833 -2353 934 -2338
rect -354 -2388 934 -2353
rect -354 -2422 -220 -2388
rect -186 -2422 -130 -2388
rect -96 -2422 -40 -2388
rect -6 -2422 50 -2388
rect 84 -2422 140 -2388
rect 174 -2422 230 -2388
rect 264 -2422 320 -2388
rect 354 -2422 410 -2388
rect 444 -2422 500 -2388
rect 534 -2422 590 -2388
rect 624 -2422 680 -2388
rect 714 -2422 770 -2388
rect 804 -2422 934 -2388
rect -354 -2454 934 -2422
rect 1006 -1201 2294 -1166
rect 1006 -1224 1140 -1201
rect 1006 -1258 1039 -1224
rect 1073 -1235 1140 -1224
rect 1174 -1235 1230 -1201
rect 1264 -1235 1320 -1201
rect 1354 -1235 1410 -1201
rect 1444 -1235 1500 -1201
rect 1534 -1235 1590 -1201
rect 1624 -1235 1680 -1201
rect 1714 -1235 1770 -1201
rect 1804 -1235 1860 -1201
rect 1894 -1235 1950 -1201
rect 1984 -1235 2040 -1201
rect 2074 -1235 2130 -1201
rect 2164 -1224 2294 -1201
rect 2164 -1235 2226 -1224
rect 1073 -1258 2226 -1235
rect 2260 -1258 2294 -1224
rect 1006 -1267 2294 -1258
rect 1006 -1314 1107 -1267
rect 1006 -1348 1039 -1314
rect 1073 -1348 1107 -1314
rect 2193 -1314 2294 -1267
rect 1006 -1404 1107 -1348
rect 1006 -1438 1039 -1404
rect 1073 -1438 1107 -1404
rect 1006 -1494 1107 -1438
rect 1006 -1528 1039 -1494
rect 1073 -1528 1107 -1494
rect 1006 -1584 1107 -1528
rect 1006 -1618 1039 -1584
rect 1073 -1618 1107 -1584
rect 1006 -1674 1107 -1618
rect 1006 -1708 1039 -1674
rect 1073 -1708 1107 -1674
rect 1006 -1764 1107 -1708
rect 1006 -1798 1039 -1764
rect 1073 -1798 1107 -1764
rect 1006 -1854 1107 -1798
rect 1006 -1888 1039 -1854
rect 1073 -1888 1107 -1854
rect 1006 -1944 1107 -1888
rect 1006 -1978 1039 -1944
rect 1073 -1978 1107 -1944
rect 1006 -2034 1107 -1978
rect 1006 -2068 1039 -2034
rect 1073 -2068 1107 -2034
rect 1006 -2124 1107 -2068
rect 1006 -2158 1039 -2124
rect 1073 -2158 1107 -2124
rect 1006 -2214 1107 -2158
rect 1006 -2248 1039 -2214
rect 1073 -2248 1107 -2214
rect 1006 -2304 1107 -2248
rect 2193 -1348 2226 -1314
rect 2260 -1348 2294 -1314
rect 2193 -1404 2294 -1348
rect 2193 -1438 2226 -1404
rect 2260 -1438 2294 -1404
rect 2193 -1494 2294 -1438
rect 2193 -1528 2226 -1494
rect 2260 -1528 2294 -1494
rect 2193 -1584 2294 -1528
rect 2193 -1618 2226 -1584
rect 2260 -1618 2294 -1584
rect 2193 -1674 2294 -1618
rect 2193 -1708 2226 -1674
rect 2260 -1708 2294 -1674
rect 2193 -1764 2294 -1708
rect 2193 -1798 2226 -1764
rect 2260 -1798 2294 -1764
rect 2193 -1854 2294 -1798
rect 2193 -1888 2226 -1854
rect 2260 -1888 2294 -1854
rect 2193 -1944 2294 -1888
rect 2193 -1978 2226 -1944
rect 2260 -1978 2294 -1944
rect 2193 -2034 2294 -1978
rect 2193 -2068 2226 -2034
rect 2260 -2068 2294 -2034
rect 2193 -2124 2294 -2068
rect 2193 -2158 2226 -2124
rect 2260 -2158 2294 -2124
rect 2990 -1450 3070 -1420
rect 2990 -1490 3010 -1450
rect 3050 -1490 3070 -1450
rect 2990 -1520 3070 -1490
rect 2193 -2214 2294 -2158
rect 2193 -2248 2226 -2214
rect 2260 -2248 2294 -2214
rect 1006 -2338 1039 -2304
rect 1073 -2338 1107 -2304
rect 1006 -2353 1107 -2338
rect 2193 -2304 2294 -2248
rect 2193 -2338 2226 -2304
rect 2260 -2338 2294 -2304
rect 2193 -2353 2294 -2338
rect 1006 -2388 2294 -2353
rect 1006 -2422 1140 -2388
rect 1174 -2422 1230 -2388
rect 1264 -2422 1320 -2388
rect 1354 -2422 1410 -2388
rect 1444 -2422 1500 -2388
rect 1534 -2422 1590 -2388
rect 1624 -2422 1680 -2388
rect 1714 -2422 1770 -2388
rect 1804 -2422 1860 -2388
rect 1894 -2422 1950 -2388
rect 1984 -2422 2040 -2388
rect 2074 -2422 2130 -2388
rect 2164 -2422 2294 -2388
rect 1006 -2454 2294 -2422
rect 240 -2540 340 -2510
rect 240 -2580 270 -2540
rect 310 -2580 340 -2540
rect 240 -2620 340 -2580
rect 240 -2660 270 -2620
rect 310 -2660 340 -2620
rect 240 -2700 340 -2660
rect 240 -2740 270 -2700
rect 310 -2740 340 -2700
rect 240 -2770 340 -2740
<< nsubdiff >>
rect -1110 12490 -1030 12520
rect -1110 12450 -1090 12490
rect -1050 12450 -1030 12490
rect -1110 12420 -1030 12450
rect 1260 12490 1340 12520
rect 1260 12450 1280 12490
rect 1320 12450 1340 12490
rect 1260 12420 1340 12450
rect 9200 12530 10210 12570
rect 10370 12530 11420 12570
rect 4130 12490 4210 12520
rect 4130 12450 4150 12490
rect 4190 12450 4210 12490
rect 4130 12420 4210 12450
rect 5430 12490 5510 12520
rect 5430 12450 5450 12490
rect 5490 12450 5510 12490
rect 5430 12420 5510 12450
rect 6730 12490 6810 12520
rect 6730 12450 6750 12490
rect 6790 12450 6810 12490
rect 6730 12420 6810 12450
rect 8030 12490 8110 12520
rect 8030 12450 8050 12490
rect 8090 12450 8110 12490
rect 8030 12420 8110 12450
rect 9200 11600 9240 12530
rect 11380 11600 11420 12530
rect 9200 10840 9240 11270
rect 11380 10840 11420 11270
rect 9200 10800 10210 10840
rect 10370 10800 11250 10840
rect 11320 10800 11420 10840
rect -720 9790 -640 9820
rect -720 9750 -700 9790
rect -660 9750 -640 9790
rect -720 9690 -640 9750
rect -720 9650 -700 9690
rect -660 9650 -640 9690
rect -720 9590 -640 9650
rect -720 9550 -700 9590
rect -660 9550 -640 9590
rect -720 9490 -640 9550
rect -720 9450 -700 9490
rect -660 9450 -640 9490
rect -720 9420 -640 9450
rect 180 9790 260 9820
rect 180 9750 200 9790
rect 240 9750 260 9790
rect 180 9690 260 9750
rect 180 9650 200 9690
rect 240 9650 260 9690
rect 180 9590 260 9650
rect 180 9550 200 9590
rect 240 9550 260 9590
rect 180 9490 260 9550
rect 180 9450 200 9490
rect 240 9450 260 9490
rect 180 9420 260 9450
rect 1080 9790 1160 9820
rect 1080 9750 1100 9790
rect 1140 9750 1160 9790
rect 1080 9690 1160 9750
rect 1080 9650 1100 9690
rect 1140 9650 1160 9690
rect 1080 9590 1160 9650
rect 1080 9550 1100 9590
rect 1140 9550 1160 9590
rect 1080 9490 1160 9550
rect 1080 9450 1100 9490
rect 1140 9450 1160 9490
rect 1080 9420 1160 9450
rect 1220 9790 1300 9820
rect 1220 9750 1240 9790
rect 1280 9750 1300 9790
rect 1220 9690 1300 9750
rect 1220 9650 1240 9690
rect 1280 9650 1300 9690
rect 1220 9590 1300 9650
rect 1220 9550 1240 9590
rect 1280 9550 1300 9590
rect 1220 9490 1300 9550
rect 1220 9450 1240 9490
rect 1280 9450 1300 9490
rect 1220 9430 1300 9450
rect 1220 9420 1280 9430
rect 1660 9790 1740 9820
rect 1660 9750 1680 9790
rect 1720 9750 1740 9790
rect 1660 9690 1740 9750
rect 1660 9650 1680 9690
rect 1720 9650 1740 9690
rect 1660 9590 1740 9650
rect 1660 9550 1680 9590
rect 1720 9550 1740 9590
rect 1660 9490 1740 9550
rect 1660 9450 1680 9490
rect 1720 9450 1740 9490
rect 1660 9420 1740 9450
rect 1990 9790 2070 9820
rect 1990 9750 2010 9790
rect 2050 9750 2070 9790
rect 1990 9690 2070 9750
rect 1990 9650 2010 9690
rect 2050 9650 2070 9690
rect 1990 9590 2070 9650
rect 1990 9550 2010 9590
rect 2050 9550 2070 9590
rect 1990 9490 2070 9550
rect 1990 9450 2010 9490
rect 2050 9450 2070 9490
rect 1990 9420 2070 9450
rect 2390 9790 2490 9820
rect 2390 9750 2420 9790
rect 2460 9750 2490 9790
rect 2390 9690 2490 9750
rect 2390 9650 2420 9690
rect 2460 9650 2490 9690
rect 2390 9590 2490 9650
rect 2390 9550 2420 9590
rect 2460 9550 2490 9590
rect 2390 9490 2490 9550
rect 2390 9450 2420 9490
rect 2460 9450 2490 9490
rect 2390 9420 2490 9450
rect 2780 9790 2880 9820
rect 2780 9750 2810 9790
rect 2850 9750 2880 9790
rect 2780 9690 2880 9750
rect 2780 9650 2810 9690
rect 2850 9650 2880 9690
rect 2780 9590 2880 9650
rect 2780 9550 2810 9590
rect 2850 9550 2880 9590
rect 2780 9490 2880 9550
rect 2780 9450 2810 9490
rect 2850 9450 2880 9490
rect 2780 9420 2880 9450
rect 3170 9790 3270 9820
rect 3170 9750 3200 9790
rect 3240 9750 3270 9790
rect 3170 9690 3270 9750
rect 3170 9650 3200 9690
rect 3240 9650 3270 9690
rect 3170 9590 3270 9650
rect 3170 9550 3200 9590
rect 3240 9550 3270 9590
rect 3170 9490 3270 9550
rect 3170 9450 3200 9490
rect 3240 9450 3270 9490
rect 3170 9420 3270 9450
rect 3850 9790 3950 9820
rect 3850 9750 3880 9790
rect 3920 9750 3950 9790
rect 3850 9690 3950 9750
rect 3850 9650 3880 9690
rect 3920 9650 3950 9690
rect 3850 9590 3950 9650
rect 3850 9550 3880 9590
rect 3920 9550 3950 9590
rect 3850 9490 3950 9550
rect 3850 9450 3880 9490
rect 3920 9450 3950 9490
rect 3850 9420 3950 9450
rect 5540 9760 5640 9790
rect 5540 9720 5570 9760
rect 5610 9720 5640 9760
rect 5540 9660 5640 9720
rect 5540 9620 5570 9660
rect 5610 9620 5640 9660
rect 5540 9560 5640 9620
rect 5540 9520 5570 9560
rect 5610 9520 5640 9560
rect 5540 9460 5640 9520
rect 5540 9420 5570 9460
rect 5610 9420 5640 9460
rect 5540 9390 5640 9420
rect 7060 9760 7160 9790
rect 7060 9720 7090 9760
rect 7130 9720 7160 9760
rect 7060 9660 7160 9720
rect 7060 9620 7090 9660
rect 7130 9620 7160 9660
rect 7060 9560 7160 9620
rect 7060 9520 7090 9560
rect 7130 9520 7160 9560
rect 7060 9460 7160 9520
rect 7060 9420 7090 9460
rect 7130 9420 7160 9460
rect 7060 9390 7160 9420
rect 8580 9760 8680 9790
rect 8580 9720 8610 9760
rect 8650 9720 8680 9760
rect 8580 9660 8680 9720
rect 8580 9620 8610 9660
rect 8650 9620 8680 9660
rect 8580 9560 8680 9620
rect 8580 9520 8610 9560
rect 8650 9520 8680 9560
rect 8580 9460 8680 9520
rect 8580 9420 8610 9460
rect 8650 9420 8680 9460
rect 8580 9390 8680 9420
rect -720 9030 -640 9060
rect -720 8990 -700 9030
rect -660 8990 -640 9030
rect -720 8930 -640 8990
rect -720 8890 -700 8930
rect -660 8890 -640 8930
rect -720 8830 -640 8890
rect -720 8790 -700 8830
rect -660 8790 -640 8830
rect -720 8730 -640 8790
rect -720 8690 -700 8730
rect -660 8690 -640 8730
rect -720 8660 -640 8690
rect 180 9030 260 9060
rect 180 8990 200 9030
rect 240 8990 260 9030
rect 180 8930 260 8990
rect 180 8890 200 8930
rect 240 8890 260 8930
rect 180 8830 260 8890
rect 180 8790 200 8830
rect 240 8790 260 8830
rect 180 8730 260 8790
rect 180 8690 200 8730
rect 240 8690 260 8730
rect 180 8660 260 8690
rect 1080 9030 1160 9060
rect 1080 8990 1100 9030
rect 1140 8990 1160 9030
rect 1080 8930 1160 8990
rect 1080 8890 1100 8930
rect 1140 8890 1160 8930
rect 1080 8830 1160 8890
rect 1080 8790 1100 8830
rect 1140 8790 1160 8830
rect 1080 8730 1160 8790
rect 1080 8690 1100 8730
rect 1140 8690 1160 8730
rect 1080 8660 1160 8690
rect 1480 9030 1560 9060
rect 1480 8990 1500 9030
rect 1540 8990 1560 9030
rect 1480 8930 1560 8990
rect 1480 8890 1500 8930
rect 1540 8890 1560 8930
rect 1480 8830 1560 8890
rect 1480 8790 1500 8830
rect 1540 8790 1560 8830
rect 1480 8730 1560 8790
rect 1480 8690 1500 8730
rect 1540 8690 1560 8730
rect 1480 8660 1560 8690
rect 1810 9030 1890 9060
rect 1810 8990 1830 9030
rect 1870 8990 1890 9030
rect 1810 8930 1890 8990
rect 1810 8890 1830 8930
rect 1870 8890 1890 8930
rect 1810 8830 1890 8890
rect 1810 8790 1830 8830
rect 1870 8790 1890 8830
rect 1810 8730 1890 8790
rect 1810 8690 1830 8730
rect 1870 8690 1890 8730
rect 1810 8660 1890 8690
rect 2140 9030 2220 9060
rect 2140 8990 2160 9030
rect 2200 8990 2220 9030
rect 2140 8930 2220 8990
rect 2140 8890 2160 8930
rect 2200 8890 2220 8930
rect 2140 8830 2220 8890
rect 2140 8790 2160 8830
rect 2200 8790 2220 8830
rect 2140 8730 2220 8790
rect 2140 8690 2160 8730
rect 2200 8690 2220 8730
rect 2140 8660 2220 8690
rect 2390 9030 2490 9060
rect 2390 8990 2420 9030
rect 2460 8990 2490 9030
rect 2390 8930 2490 8990
rect 2390 8890 2420 8930
rect 2460 8890 2490 8930
rect 2390 8830 2490 8890
rect 2390 8790 2420 8830
rect 2460 8790 2490 8830
rect 2390 8730 2490 8790
rect 2390 8690 2420 8730
rect 2460 8690 2490 8730
rect 2390 8660 2490 8690
rect 3170 9030 3270 9060
rect 3170 8990 3200 9030
rect 3240 8990 3270 9030
rect 3170 8930 3270 8990
rect 3170 8890 3200 8930
rect 3240 8890 3270 8930
rect 3170 8830 3270 8890
rect 3170 8790 3200 8830
rect 3240 8790 3270 8830
rect 3170 8730 3270 8790
rect 3170 8690 3200 8730
rect 3240 8690 3270 8730
rect 3170 8660 3270 8690
rect -1440 6840 -1360 6870
rect -1440 6800 -1420 6840
rect -1380 6800 -1360 6840
rect -1440 6740 -1360 6800
rect -1440 6700 -1420 6740
rect -1380 6700 -1360 6740
rect -1440 6670 -1360 6700
rect 40 6840 120 6870
rect 40 6800 60 6840
rect 100 6800 120 6840
rect 40 6740 120 6800
rect 40 6700 60 6740
rect 100 6700 120 6740
rect 40 6670 120 6700
rect 460 6840 540 6870
rect 460 6800 480 6840
rect 520 6800 540 6840
rect 460 6740 540 6800
rect 460 6700 480 6740
rect 520 6700 540 6740
rect 460 6670 540 6700
rect 1940 6840 2020 6870
rect 1940 6800 1960 6840
rect 2000 6800 2020 6840
rect 1940 6740 2020 6800
rect 1940 6700 1960 6740
rect 2000 6700 2020 6740
rect 1940 6670 2020 6700
rect -1450 6240 -1370 6270
rect -1450 6200 -1430 6240
rect -1390 6200 -1370 6240
rect -1450 6140 -1370 6200
rect -1450 6100 -1430 6140
rect -1390 6100 -1370 6140
rect -1450 6040 -1370 6100
rect -1450 6000 -1430 6040
rect -1390 6000 -1370 6040
rect -1450 5940 -1370 6000
rect -1450 5900 -1430 5940
rect -1390 5900 -1370 5940
rect -1450 5840 -1370 5900
rect -1450 5800 -1430 5840
rect -1390 5800 -1370 5840
rect -1450 5740 -1370 5800
rect -1450 5700 -1430 5740
rect -1390 5700 -1370 5740
rect -1450 5670 -1370 5700
rect 1950 6240 2030 6270
rect 1950 6200 1970 6240
rect 2010 6200 2030 6240
rect 1950 6140 2030 6200
rect 1950 6100 1970 6140
rect 2010 6100 2030 6140
rect 1950 6040 2030 6100
rect 1950 6000 1970 6040
rect 2010 6000 2030 6040
rect 1950 5940 2030 6000
rect 1950 5900 1970 5940
rect 2010 5900 2030 5940
rect 1950 5840 2030 5900
rect 2410 6040 2490 6070
rect 2410 6000 2430 6040
rect 2470 6000 2490 6040
rect 2410 5940 2490 6000
rect 2410 5900 2430 5940
rect 2470 5900 2490 5940
rect 2410 5870 2490 5900
rect 3020 6040 3100 6070
rect 3020 6000 3040 6040
rect 3080 6000 3100 6040
rect 3020 5940 3100 6000
rect 3020 5900 3040 5940
rect 3080 5900 3100 5940
rect 3020 5870 3100 5900
rect 1950 5800 1970 5840
rect 2010 5800 2030 5840
rect 1950 5740 2030 5800
rect 1950 5700 1970 5740
rect 2010 5700 2030 5740
rect 1950 5670 2030 5700
rect -2550 4680 -2470 4710
rect -2550 4640 -2530 4680
rect -2490 4640 -2470 4680
rect -2550 4580 -2470 4640
rect -2550 4540 -2530 4580
rect -2490 4540 -2470 4580
rect -2550 4510 -2470 4540
rect 10 4680 90 4710
rect 10 4640 30 4680
rect 70 4640 90 4680
rect 10 4580 90 4640
rect 10 4540 30 4580
rect 70 4540 90 4580
rect 10 4510 90 4540
rect 490 4680 570 4710
rect 490 4640 510 4680
rect 550 4640 570 4680
rect 490 4580 570 4640
rect 490 4540 510 4580
rect 550 4540 570 4580
rect 490 4510 570 4540
rect 3050 4680 3130 4710
rect 3050 4640 3070 4680
rect 3110 4640 3130 4680
rect 3050 4580 3130 4640
rect 6590 4760 6690 4790
rect 6590 4720 6620 4760
rect 6660 4720 6690 4760
rect 6590 4660 6690 4720
rect 6590 4620 6620 4660
rect 6660 4620 6690 4660
rect 6590 4590 6690 4620
rect 7570 4760 7670 4790
rect 7570 4720 7600 4760
rect 7640 4720 7670 4760
rect 7570 4660 7670 4720
rect 7570 4620 7600 4660
rect 7640 4620 7670 4660
rect 7570 4590 7670 4620
rect 7730 4760 7830 4790
rect 7730 4720 7760 4760
rect 7800 4720 7830 4760
rect 7730 4660 7830 4720
rect 7730 4620 7760 4660
rect 7800 4620 7830 4660
rect 7730 4590 7830 4620
rect 8710 4760 8810 4790
rect 8710 4720 8740 4760
rect 8780 4720 8810 4760
rect 8710 4660 8810 4720
rect 8710 4620 8740 4660
rect 8780 4620 8810 4660
rect 8710 4590 8810 4620
rect 3050 4540 3070 4580
rect 3110 4540 3130 4580
rect 3050 4510 3130 4540
rect 5520 4110 5620 4140
rect 5520 4070 5550 4110
rect 5590 4070 5620 4110
rect 5520 4010 5620 4070
rect 5520 3970 5550 4010
rect 5590 3970 5620 4010
rect 5520 3910 5620 3970
rect 5520 3870 5550 3910
rect 5590 3870 5620 3910
rect 5520 3810 5620 3870
rect 5520 3770 5550 3810
rect 5590 3770 5620 3810
rect 5520 3710 5620 3770
rect 5520 3670 5550 3710
rect 5590 3670 5620 3710
rect 5520 3640 5620 3670
rect 7720 4110 7820 4140
rect 7720 4070 7750 4110
rect 7790 4070 7820 4110
rect 7720 4010 7820 4070
rect 7720 3970 7750 4010
rect 7790 3970 7820 4010
rect 7720 3910 7820 3970
rect 7720 3870 7750 3910
rect 7790 3870 7820 3910
rect 7720 3810 7820 3870
rect 7720 3770 7750 3810
rect 7790 3770 7820 3810
rect 7720 3710 7820 3770
rect 7720 3670 7750 3710
rect 7790 3670 7820 3710
rect 7720 3640 7820 3670
rect -1551 1372 -589 1391
rect -1551 1338 -1474 1372
rect -1440 1338 -1384 1372
rect -1350 1338 -1294 1372
rect -1260 1338 -1204 1372
rect -1170 1338 -1114 1372
rect -1080 1338 -1024 1372
rect -990 1338 -934 1372
rect -900 1338 -844 1372
rect -810 1338 -754 1372
rect -720 1338 -589 1372
rect -1551 1319 -589 1338
rect -1551 1296 -1479 1319
rect -1551 1262 -1532 1296
rect -1498 1262 -1479 1296
rect -1551 1206 -1479 1262
rect -661 1315 -589 1319
rect -661 1281 -642 1315
rect -608 1281 -589 1315
rect -1551 1172 -1532 1206
rect -1498 1172 -1479 1206
rect -1551 1116 -1479 1172
rect -1551 1082 -1532 1116
rect -1498 1082 -1479 1116
rect -1551 1026 -1479 1082
rect -1551 992 -1532 1026
rect -1498 992 -1479 1026
rect -1551 936 -1479 992
rect -1551 902 -1532 936
rect -1498 902 -1479 936
rect -1551 846 -1479 902
rect -1551 812 -1532 846
rect -1498 812 -1479 846
rect -1551 756 -1479 812
rect -1551 722 -1532 756
rect -1498 722 -1479 756
rect -1551 666 -1479 722
rect -1551 632 -1532 666
rect -1498 632 -1479 666
rect -1551 576 -1479 632
rect -1551 542 -1532 576
rect -1498 542 -1479 576
rect -661 1225 -589 1281
rect -661 1191 -642 1225
rect -608 1191 -589 1225
rect -661 1135 -589 1191
rect -661 1101 -642 1135
rect -608 1101 -589 1135
rect -661 1045 -589 1101
rect -661 1011 -642 1045
rect -608 1011 -589 1045
rect -661 955 -589 1011
rect -661 921 -642 955
rect -608 921 -589 955
rect -661 865 -589 921
rect -661 831 -642 865
rect -608 831 -589 865
rect -661 775 -589 831
rect -661 741 -642 775
rect -608 741 -589 775
rect -661 685 -589 741
rect -661 651 -642 685
rect -608 651 -589 685
rect -661 595 -589 651
rect -1551 501 -1479 542
rect -661 561 -642 595
rect -608 561 -589 595
rect -661 501 -589 561
rect -1551 482 -589 501
rect -1551 448 -1440 482
rect -1406 448 -1350 482
rect -1316 448 -1260 482
rect -1226 448 -1170 482
rect -1136 448 -1080 482
rect -1046 448 -990 482
rect -956 448 -900 482
rect -866 448 -810 482
rect -776 448 -720 482
rect -686 448 -589 482
rect -1551 429 -589 448
rect -191 1372 771 1391
rect -191 1338 -114 1372
rect -80 1338 -24 1372
rect 10 1338 66 1372
rect 100 1338 156 1372
rect 190 1338 246 1372
rect 280 1338 336 1372
rect 370 1338 426 1372
rect 460 1338 516 1372
rect 550 1338 606 1372
rect 640 1338 771 1372
rect -191 1319 771 1338
rect -191 1296 -119 1319
rect -191 1262 -172 1296
rect -138 1262 -119 1296
rect -191 1206 -119 1262
rect 699 1315 771 1319
rect 699 1281 718 1315
rect 752 1281 771 1315
rect -191 1172 -172 1206
rect -138 1172 -119 1206
rect -191 1116 -119 1172
rect -191 1082 -172 1116
rect -138 1082 -119 1116
rect -191 1026 -119 1082
rect -191 992 -172 1026
rect -138 992 -119 1026
rect -191 936 -119 992
rect -191 902 -172 936
rect -138 902 -119 936
rect -191 846 -119 902
rect -191 812 -172 846
rect -138 812 -119 846
rect -191 756 -119 812
rect -191 722 -172 756
rect -138 722 -119 756
rect -191 666 -119 722
rect -191 632 -172 666
rect -138 632 -119 666
rect -191 576 -119 632
rect -191 542 -172 576
rect -138 542 -119 576
rect 699 1225 771 1281
rect 699 1191 718 1225
rect 752 1191 771 1225
rect 699 1135 771 1191
rect 699 1101 718 1135
rect 752 1101 771 1135
rect 699 1045 771 1101
rect 699 1011 718 1045
rect 752 1011 771 1045
rect 699 955 771 1011
rect 699 921 718 955
rect 752 921 771 955
rect 699 865 771 921
rect 699 831 718 865
rect 752 831 771 865
rect 699 775 771 831
rect 699 741 718 775
rect 752 741 771 775
rect 699 685 771 741
rect 699 651 718 685
rect 752 651 771 685
rect 699 595 771 651
rect -191 501 -119 542
rect 699 561 718 595
rect 752 561 771 595
rect 699 501 771 561
rect -191 482 771 501
rect -191 448 -80 482
rect -46 448 10 482
rect 44 448 100 482
rect 134 448 190 482
rect 224 448 280 482
rect 314 448 370 482
rect 404 448 460 482
rect 494 448 550 482
rect 584 448 640 482
rect 674 448 771 482
rect -191 429 771 448
rect 1169 1372 2131 1391
rect 1169 1338 1246 1372
rect 1280 1338 1336 1372
rect 1370 1338 1426 1372
rect 1460 1338 1516 1372
rect 1550 1338 1606 1372
rect 1640 1338 1696 1372
rect 1730 1338 1786 1372
rect 1820 1338 1876 1372
rect 1910 1338 1966 1372
rect 2000 1338 2131 1372
rect 1169 1319 2131 1338
rect 1169 1296 1241 1319
rect 1169 1262 1188 1296
rect 1222 1262 1241 1296
rect 1169 1206 1241 1262
rect 2059 1315 2131 1319
rect 2059 1281 2078 1315
rect 2112 1281 2131 1315
rect 1169 1172 1188 1206
rect 1222 1172 1241 1206
rect 1169 1116 1241 1172
rect 1169 1082 1188 1116
rect 1222 1082 1241 1116
rect 1169 1026 1241 1082
rect 1169 992 1188 1026
rect 1222 992 1241 1026
rect 1169 936 1241 992
rect 1169 902 1188 936
rect 1222 902 1241 936
rect 1169 846 1241 902
rect 1169 812 1188 846
rect 1222 812 1241 846
rect 1169 756 1241 812
rect 1169 722 1188 756
rect 1222 722 1241 756
rect 1169 666 1241 722
rect 1169 632 1188 666
rect 1222 632 1241 666
rect 1169 576 1241 632
rect 1169 542 1188 576
rect 1222 542 1241 576
rect 2059 1225 2131 1281
rect 2059 1191 2078 1225
rect 2112 1191 2131 1225
rect 2059 1135 2131 1191
rect 2059 1101 2078 1135
rect 2112 1101 2131 1135
rect 2059 1045 2131 1101
rect 2059 1011 2078 1045
rect 2112 1011 2131 1045
rect 2059 955 2131 1011
rect 2059 921 2078 955
rect 2112 921 2131 955
rect 2059 865 2131 921
rect 2059 831 2078 865
rect 2112 831 2131 865
rect 2059 775 2131 831
rect 2059 741 2078 775
rect 2112 741 2131 775
rect 2059 685 2131 741
rect 2059 651 2078 685
rect 2112 651 2131 685
rect 2059 595 2131 651
rect 1169 501 1241 542
rect 2059 561 2078 595
rect 2112 561 2131 595
rect 2059 501 2131 561
rect 1169 482 2131 501
rect 1169 448 1280 482
rect 1314 448 1370 482
rect 1404 448 1460 482
rect 1494 448 1550 482
rect 1584 448 1640 482
rect 1674 448 1730 482
rect 1764 448 1820 482
rect 1854 448 1910 482
rect 1944 448 2000 482
rect 2034 448 2131 482
rect 1169 429 2131 448
rect -1551 12 -589 31
rect -1551 -22 -1474 12
rect -1440 -22 -1384 12
rect -1350 -22 -1294 12
rect -1260 -22 -1204 12
rect -1170 -22 -1114 12
rect -1080 -22 -1024 12
rect -990 -22 -934 12
rect -900 -22 -844 12
rect -810 -22 -754 12
rect -720 -22 -589 12
rect -1551 -41 -589 -22
rect -1551 -64 -1479 -41
rect -1551 -98 -1532 -64
rect -1498 -98 -1479 -64
rect -1551 -154 -1479 -98
rect -661 -45 -589 -41
rect -661 -79 -642 -45
rect -608 -79 -589 -45
rect -1551 -188 -1532 -154
rect -1498 -188 -1479 -154
rect -1551 -244 -1479 -188
rect -1551 -278 -1532 -244
rect -1498 -278 -1479 -244
rect -1551 -334 -1479 -278
rect -1551 -368 -1532 -334
rect -1498 -368 -1479 -334
rect -1551 -424 -1479 -368
rect -1551 -458 -1532 -424
rect -1498 -458 -1479 -424
rect -1551 -514 -1479 -458
rect -1551 -548 -1532 -514
rect -1498 -548 -1479 -514
rect -1551 -604 -1479 -548
rect -1551 -638 -1532 -604
rect -1498 -638 -1479 -604
rect -1551 -694 -1479 -638
rect -1551 -728 -1532 -694
rect -1498 -728 -1479 -694
rect -1551 -784 -1479 -728
rect -1551 -818 -1532 -784
rect -1498 -818 -1479 -784
rect -661 -135 -589 -79
rect -661 -169 -642 -135
rect -608 -169 -589 -135
rect -661 -225 -589 -169
rect -661 -259 -642 -225
rect -608 -259 -589 -225
rect -661 -315 -589 -259
rect -661 -349 -642 -315
rect -608 -349 -589 -315
rect -661 -405 -589 -349
rect -661 -439 -642 -405
rect -608 -439 -589 -405
rect -661 -495 -589 -439
rect -661 -529 -642 -495
rect -608 -529 -589 -495
rect -661 -585 -589 -529
rect -661 -619 -642 -585
rect -608 -619 -589 -585
rect -661 -675 -589 -619
rect -661 -709 -642 -675
rect -608 -709 -589 -675
rect -661 -765 -589 -709
rect -1551 -859 -1479 -818
rect -661 -799 -642 -765
rect -608 -799 -589 -765
rect -661 -859 -589 -799
rect -1551 -878 -589 -859
rect -1551 -912 -1440 -878
rect -1406 -912 -1350 -878
rect -1316 -912 -1260 -878
rect -1226 -912 -1170 -878
rect -1136 -912 -1080 -878
rect -1046 -912 -990 -878
rect -956 -912 -900 -878
rect -866 -912 -810 -878
rect -776 -912 -720 -878
rect -686 -912 -589 -878
rect -1551 -931 -589 -912
rect -191 12 771 31
rect -191 -22 -114 12
rect -80 -22 -24 12
rect 10 -22 66 12
rect 100 -22 156 12
rect 190 -22 246 12
rect 280 -22 336 12
rect 370 -22 426 12
rect 460 -22 516 12
rect 550 -22 606 12
rect 640 -22 771 12
rect -191 -41 771 -22
rect -191 -64 -119 -41
rect -191 -98 -172 -64
rect -138 -98 -119 -64
rect -191 -154 -119 -98
rect 699 -45 771 -41
rect 699 -79 718 -45
rect 752 -79 771 -45
rect -191 -188 -172 -154
rect -138 -188 -119 -154
rect -191 -244 -119 -188
rect -191 -278 -172 -244
rect -138 -278 -119 -244
rect -191 -334 -119 -278
rect -191 -368 -172 -334
rect -138 -368 -119 -334
rect -191 -424 -119 -368
rect -191 -458 -172 -424
rect -138 -458 -119 -424
rect -191 -514 -119 -458
rect -191 -548 -172 -514
rect -138 -548 -119 -514
rect -191 -604 -119 -548
rect -191 -638 -172 -604
rect -138 -638 -119 -604
rect -191 -694 -119 -638
rect -191 -728 -172 -694
rect -138 -728 -119 -694
rect -191 -784 -119 -728
rect -191 -818 -172 -784
rect -138 -818 -119 -784
rect 699 -135 771 -79
rect 699 -169 718 -135
rect 752 -169 771 -135
rect 699 -225 771 -169
rect 699 -259 718 -225
rect 752 -259 771 -225
rect 699 -315 771 -259
rect 699 -349 718 -315
rect 752 -349 771 -315
rect 699 -405 771 -349
rect 699 -439 718 -405
rect 752 -439 771 -405
rect 699 -495 771 -439
rect 699 -529 718 -495
rect 752 -529 771 -495
rect 699 -585 771 -529
rect 699 -619 718 -585
rect 752 -619 771 -585
rect 699 -675 771 -619
rect 699 -709 718 -675
rect 752 -709 771 -675
rect 699 -765 771 -709
rect -191 -859 -119 -818
rect 699 -799 718 -765
rect 752 -799 771 -765
rect 699 -859 771 -799
rect -191 -878 771 -859
rect -191 -912 -80 -878
rect -46 -912 10 -878
rect 44 -912 100 -878
rect 134 -912 190 -878
rect 224 -912 280 -878
rect 314 -912 370 -878
rect 404 -912 460 -878
rect 494 -912 550 -878
rect 584 -912 640 -878
rect 674 -912 771 -878
rect -191 -931 771 -912
rect 1169 12 2131 31
rect 1169 -22 1246 12
rect 1280 -22 1336 12
rect 1370 -22 1426 12
rect 1460 -22 1516 12
rect 1550 -22 1606 12
rect 1640 -22 1696 12
rect 1730 -22 1786 12
rect 1820 -22 1876 12
rect 1910 -22 1966 12
rect 2000 -22 2131 12
rect 1169 -41 2131 -22
rect 1169 -64 1241 -41
rect 1169 -98 1188 -64
rect 1222 -98 1241 -64
rect 1169 -154 1241 -98
rect 2059 -45 2131 -41
rect 2059 -79 2078 -45
rect 2112 -79 2131 -45
rect 1169 -188 1188 -154
rect 1222 -188 1241 -154
rect 1169 -244 1241 -188
rect 1169 -278 1188 -244
rect 1222 -278 1241 -244
rect 1169 -334 1241 -278
rect 1169 -368 1188 -334
rect 1222 -368 1241 -334
rect 1169 -424 1241 -368
rect 1169 -458 1188 -424
rect 1222 -458 1241 -424
rect 1169 -514 1241 -458
rect 1169 -548 1188 -514
rect 1222 -548 1241 -514
rect 1169 -604 1241 -548
rect 1169 -638 1188 -604
rect 1222 -638 1241 -604
rect 1169 -694 1241 -638
rect 1169 -728 1188 -694
rect 1222 -728 1241 -694
rect 1169 -784 1241 -728
rect 1169 -818 1188 -784
rect 1222 -818 1241 -784
rect 2059 -135 2131 -79
rect 2059 -169 2078 -135
rect 2112 -169 2131 -135
rect 2059 -225 2131 -169
rect 2059 -259 2078 -225
rect 2112 -259 2131 -225
rect 2059 -315 2131 -259
rect 2059 -349 2078 -315
rect 2112 -349 2131 -315
rect 2059 -405 2131 -349
rect 2059 -439 2078 -405
rect 2112 -439 2131 -405
rect 2059 -495 2131 -439
rect 2059 -529 2078 -495
rect 2112 -529 2131 -495
rect 2059 -585 2131 -529
rect 2059 -619 2078 -585
rect 2112 -619 2131 -585
rect 2059 -675 2131 -619
rect 2059 -709 2078 -675
rect 2112 -709 2131 -675
rect 2059 -765 2131 -709
rect 1169 -859 1241 -818
rect 2059 -799 2078 -765
rect 2112 -799 2131 -765
rect 2059 -859 2131 -799
rect 1169 -878 2131 -859
rect 1169 -912 1280 -878
rect 1314 -912 1370 -878
rect 1404 -912 1460 -878
rect 1494 -912 1550 -878
rect 1584 -912 1640 -878
rect 1674 -912 1730 -878
rect 1764 -912 1820 -878
rect 1854 -912 1910 -878
rect 1944 -912 2000 -878
rect 2034 -912 2131 -878
rect 1169 -931 2131 -912
rect -1551 -1348 -589 -1329
rect -1551 -1382 -1474 -1348
rect -1440 -1382 -1384 -1348
rect -1350 -1382 -1294 -1348
rect -1260 -1382 -1204 -1348
rect -1170 -1382 -1114 -1348
rect -1080 -1382 -1024 -1348
rect -990 -1382 -934 -1348
rect -900 -1382 -844 -1348
rect -810 -1382 -754 -1348
rect -720 -1382 -589 -1348
rect -1551 -1401 -589 -1382
rect -1551 -1424 -1479 -1401
rect -1551 -1458 -1532 -1424
rect -1498 -1458 -1479 -1424
rect -1551 -1514 -1479 -1458
rect -661 -1405 -589 -1401
rect -661 -1439 -642 -1405
rect -608 -1439 -589 -1405
rect -1551 -1548 -1532 -1514
rect -1498 -1548 -1479 -1514
rect -1551 -1604 -1479 -1548
rect -1551 -1638 -1532 -1604
rect -1498 -1638 -1479 -1604
rect -1551 -1694 -1479 -1638
rect -1551 -1728 -1532 -1694
rect -1498 -1728 -1479 -1694
rect -1551 -1784 -1479 -1728
rect -1551 -1818 -1532 -1784
rect -1498 -1818 -1479 -1784
rect -1551 -1874 -1479 -1818
rect -1551 -1908 -1532 -1874
rect -1498 -1908 -1479 -1874
rect -1551 -1964 -1479 -1908
rect -1551 -1998 -1532 -1964
rect -1498 -1998 -1479 -1964
rect -1551 -2054 -1479 -1998
rect -1551 -2088 -1532 -2054
rect -1498 -2088 -1479 -2054
rect -1551 -2144 -1479 -2088
rect -1551 -2178 -1532 -2144
rect -1498 -2178 -1479 -2144
rect -661 -1495 -589 -1439
rect -661 -1529 -642 -1495
rect -608 -1529 -589 -1495
rect -661 -1585 -589 -1529
rect -661 -1619 -642 -1585
rect -608 -1619 -589 -1585
rect -661 -1675 -589 -1619
rect -661 -1709 -642 -1675
rect -608 -1709 -589 -1675
rect -661 -1765 -589 -1709
rect -661 -1799 -642 -1765
rect -608 -1799 -589 -1765
rect -661 -1855 -589 -1799
rect -661 -1889 -642 -1855
rect -608 -1889 -589 -1855
rect -661 -1945 -589 -1889
rect -661 -1979 -642 -1945
rect -608 -1979 -589 -1945
rect -661 -2035 -589 -1979
rect -661 -2069 -642 -2035
rect -608 -2069 -589 -2035
rect -661 -2125 -589 -2069
rect -1551 -2219 -1479 -2178
rect -661 -2159 -642 -2125
rect -608 -2159 -589 -2125
rect -661 -2219 -589 -2159
rect -1551 -2238 -589 -2219
rect -1551 -2272 -1440 -2238
rect -1406 -2272 -1350 -2238
rect -1316 -2272 -1260 -2238
rect -1226 -2272 -1170 -2238
rect -1136 -2272 -1080 -2238
rect -1046 -2272 -990 -2238
rect -956 -2272 -900 -2238
rect -866 -2272 -810 -2238
rect -776 -2272 -720 -2238
rect -686 -2272 -589 -2238
rect -1551 -2291 -589 -2272
rect -191 -1348 771 -1329
rect -191 -1382 -114 -1348
rect -80 -1382 -24 -1348
rect 10 -1382 66 -1348
rect 100 -1382 156 -1348
rect 190 -1382 246 -1348
rect 280 -1382 336 -1348
rect 370 -1382 426 -1348
rect 460 -1382 516 -1348
rect 550 -1382 606 -1348
rect 640 -1382 771 -1348
rect -191 -1401 771 -1382
rect -191 -1424 -119 -1401
rect -191 -1458 -172 -1424
rect -138 -1458 -119 -1424
rect -191 -1514 -119 -1458
rect 699 -1405 771 -1401
rect 699 -1439 718 -1405
rect 752 -1439 771 -1405
rect -191 -1548 -172 -1514
rect -138 -1548 -119 -1514
rect -191 -1604 -119 -1548
rect -191 -1638 -172 -1604
rect -138 -1638 -119 -1604
rect -191 -1694 -119 -1638
rect -191 -1728 -172 -1694
rect -138 -1728 -119 -1694
rect -191 -1784 -119 -1728
rect -191 -1818 -172 -1784
rect -138 -1818 -119 -1784
rect -191 -1874 -119 -1818
rect -191 -1908 -172 -1874
rect -138 -1908 -119 -1874
rect -191 -1964 -119 -1908
rect -191 -1998 -172 -1964
rect -138 -1998 -119 -1964
rect -191 -2054 -119 -1998
rect -191 -2088 -172 -2054
rect -138 -2088 -119 -2054
rect -191 -2144 -119 -2088
rect -191 -2178 -172 -2144
rect -138 -2178 -119 -2144
rect 699 -1495 771 -1439
rect 699 -1529 718 -1495
rect 752 -1529 771 -1495
rect 699 -1585 771 -1529
rect 699 -1619 718 -1585
rect 752 -1619 771 -1585
rect 699 -1675 771 -1619
rect 699 -1709 718 -1675
rect 752 -1709 771 -1675
rect 699 -1765 771 -1709
rect 699 -1799 718 -1765
rect 752 -1799 771 -1765
rect 699 -1855 771 -1799
rect 699 -1889 718 -1855
rect 752 -1889 771 -1855
rect 699 -1945 771 -1889
rect 699 -1979 718 -1945
rect 752 -1979 771 -1945
rect 699 -2035 771 -1979
rect 699 -2069 718 -2035
rect 752 -2069 771 -2035
rect 699 -2125 771 -2069
rect -191 -2219 -119 -2178
rect 699 -2159 718 -2125
rect 752 -2159 771 -2125
rect 699 -2219 771 -2159
rect -191 -2238 771 -2219
rect -191 -2272 -80 -2238
rect -46 -2272 10 -2238
rect 44 -2272 100 -2238
rect 134 -2272 190 -2238
rect 224 -2272 280 -2238
rect 314 -2272 370 -2238
rect 404 -2272 460 -2238
rect 494 -2272 550 -2238
rect 584 -2272 640 -2238
rect 674 -2272 771 -2238
rect -191 -2291 771 -2272
rect 1169 -1348 2131 -1329
rect 1169 -1382 1246 -1348
rect 1280 -1382 1336 -1348
rect 1370 -1382 1426 -1348
rect 1460 -1382 1516 -1348
rect 1550 -1382 1606 -1348
rect 1640 -1382 1696 -1348
rect 1730 -1382 1786 -1348
rect 1820 -1382 1876 -1348
rect 1910 -1382 1966 -1348
rect 2000 -1382 2131 -1348
rect 1169 -1401 2131 -1382
rect 1169 -1424 1241 -1401
rect 1169 -1458 1188 -1424
rect 1222 -1458 1241 -1424
rect 1169 -1514 1241 -1458
rect 2059 -1405 2131 -1401
rect 2059 -1439 2078 -1405
rect 2112 -1439 2131 -1405
rect 1169 -1548 1188 -1514
rect 1222 -1548 1241 -1514
rect 1169 -1604 1241 -1548
rect 1169 -1638 1188 -1604
rect 1222 -1638 1241 -1604
rect 1169 -1694 1241 -1638
rect 1169 -1728 1188 -1694
rect 1222 -1728 1241 -1694
rect 1169 -1784 1241 -1728
rect 1169 -1818 1188 -1784
rect 1222 -1818 1241 -1784
rect 1169 -1874 1241 -1818
rect 1169 -1908 1188 -1874
rect 1222 -1908 1241 -1874
rect 1169 -1964 1241 -1908
rect 1169 -1998 1188 -1964
rect 1222 -1998 1241 -1964
rect 1169 -2054 1241 -1998
rect 1169 -2088 1188 -2054
rect 1222 -2088 1241 -2054
rect 1169 -2144 1241 -2088
rect 1169 -2178 1188 -2144
rect 1222 -2178 1241 -2144
rect 2059 -1495 2131 -1439
rect 2059 -1529 2078 -1495
rect 2112 -1529 2131 -1495
rect 2059 -1585 2131 -1529
rect 2059 -1619 2078 -1585
rect 2112 -1619 2131 -1585
rect 2059 -1675 2131 -1619
rect 2059 -1709 2078 -1675
rect 2112 -1709 2131 -1675
rect 2059 -1765 2131 -1709
rect 2059 -1799 2078 -1765
rect 2112 -1799 2131 -1765
rect 2059 -1855 2131 -1799
rect 2059 -1889 2078 -1855
rect 2112 -1889 2131 -1855
rect 2059 -1945 2131 -1889
rect 2059 -1979 2078 -1945
rect 2112 -1979 2131 -1945
rect 2059 -2035 2131 -1979
rect 2059 -2069 2078 -2035
rect 2112 -2069 2131 -2035
rect 2059 -2125 2131 -2069
rect 1169 -2219 1241 -2178
rect 2059 -2159 2078 -2125
rect 2112 -2159 2131 -2125
rect 2059 -2219 2131 -2159
rect 1169 -2238 2131 -2219
rect 1169 -2272 1280 -2238
rect 1314 -2272 1370 -2238
rect 1404 -2272 1460 -2238
rect 1494 -2272 1550 -2238
rect 1584 -2272 1640 -2238
rect 1674 -2272 1730 -2238
rect 1764 -2272 1820 -2238
rect 1854 -2272 1910 -2238
rect 1944 -2272 2000 -2238
rect 2034 -2272 2131 -2238
rect 1169 -2291 2131 -2272
<< psubdiffcont >>
rect 10330 13850 10470 13890
rect 9200 13210 9240 13470
rect 11190 13210 11230 13470
rect 5050 12860 5090 12900
rect 1810 12770 1850 12810
rect 3260 12770 3300 12810
rect 6350 12860 6390 12900
rect 7650 12860 7690 12900
rect 10330 12730 10470 12770
rect -700 10170 -660 10210
rect -700 10070 -660 10110
rect 200 10170 240 10210
rect 200 10070 240 10110
rect 1100 10170 1140 10210
rect 1100 10070 1140 10110
rect 1240 10170 1280 10210
rect 1240 10070 1280 10110
rect 1680 10170 1720 10210
rect 1680 10070 1720 10110
rect 2010 10170 2050 10210
rect 2010 10070 2050 10110
rect 2430 10170 2470 10210
rect 2430 10070 2470 10110
rect 2820 10170 2860 10210
rect 2820 10070 2860 10110
rect 3210 10170 3250 10210
rect 3210 10070 3250 10110
rect 5370 8620 5410 8660
rect 5370 8520 5410 8560
rect -700 8370 -660 8410
rect -700 8270 -660 8310
rect 200 8370 240 8410
rect 200 8270 240 8310
rect 1100 8370 1140 8410
rect 1100 8270 1140 8310
rect 1500 8370 1540 8410
rect 1500 8270 1540 8310
rect 1830 8370 1870 8410
rect 1830 8270 1870 8310
rect 2160 8370 2200 8410
rect 2160 8270 2200 8310
rect 2420 8370 2460 8410
rect 2420 8270 2460 8310
rect 3200 8370 3240 8410
rect 3200 8270 3240 8310
rect 3880 8370 3920 8410
rect 3880 8270 3920 8310
rect 5370 8420 5410 8460
rect 5370 8320 5410 8360
rect 6450 8620 6490 8660
rect 6450 8520 6490 8560
rect 6450 8420 6490 8460
rect 6450 8320 6490 8360
rect 7530 8620 7570 8660
rect 7530 8520 7570 8560
rect 7530 8420 7570 8460
rect 7530 8320 7570 8360
rect 8610 8620 8650 8660
rect 8610 8520 8650 8560
rect 8610 8420 8650 8460
rect 8610 8320 8650 8360
rect 5430 5980 5470 6030
rect 5430 5840 5470 5890
rect 7630 5980 7670 6030
rect 7630 5840 7670 5890
rect 5480 5300 5520 5340
rect 6460 5300 6500 5340
rect 7760 5300 7800 5340
rect 8740 5300 8780 5340
rect -170 3770 -130 3810
rect -170 3690 -130 3730
rect -170 3610 -130 3650
rect 710 3770 750 3810
rect 710 3690 750 3730
rect 710 3610 750 3650
rect -1070 3090 -1030 3130
rect -1070 2990 -1030 3030
rect -1070 2890 -1030 2930
rect -1070 2790 -1030 2830
rect -1070 2690 -1030 2730
rect 1610 3090 1650 3130
rect 1610 2990 1650 3030
rect 1610 2890 1650 2930
rect 1610 2790 1650 2830
rect 1610 2690 1650 2730
rect 2430 2180 2470 2220
rect 2430 2080 2470 2120
rect -1681 1462 -1647 1496
rect -1580 1485 -1546 1519
rect -1490 1485 -1456 1519
rect -1400 1485 -1366 1519
rect -1310 1485 -1276 1519
rect -1220 1485 -1186 1519
rect -1130 1485 -1096 1519
rect -1040 1485 -1006 1519
rect -950 1485 -916 1519
rect -860 1485 -826 1519
rect -770 1485 -736 1519
rect -680 1485 -646 1519
rect -590 1485 -556 1519
rect -494 1462 -460 1496
rect -1681 1372 -1647 1406
rect -1681 1282 -1647 1316
rect -1681 1192 -1647 1226
rect -1681 1102 -1647 1136
rect -1681 1012 -1647 1046
rect -1681 922 -1647 956
rect -1681 832 -1647 866
rect -1681 742 -1647 776
rect -1681 652 -1647 686
rect -1681 562 -1647 596
rect -1681 472 -1647 506
rect -494 1372 -460 1406
rect -494 1282 -460 1316
rect -494 1192 -460 1226
rect -494 1102 -460 1136
rect -494 1012 -460 1046
rect -494 922 -460 956
rect -494 832 -460 866
rect -494 742 -460 776
rect -494 652 -460 686
rect -494 562 -460 596
rect -494 472 -460 506
rect -1681 382 -1647 416
rect -494 382 -460 416
rect -1580 298 -1546 332
rect -1490 298 -1456 332
rect -1400 298 -1366 332
rect -1310 298 -1276 332
rect -1220 298 -1186 332
rect -1130 298 -1096 332
rect -1040 298 -1006 332
rect -950 298 -916 332
rect -860 298 -826 332
rect -770 298 -736 332
rect -680 298 -646 332
rect -590 298 -556 332
rect -321 1462 -287 1496
rect -220 1485 -186 1519
rect -130 1485 -96 1519
rect -40 1485 -6 1519
rect 50 1485 84 1519
rect 140 1485 174 1519
rect 230 1485 264 1519
rect 320 1485 354 1519
rect 410 1485 444 1519
rect 500 1485 534 1519
rect 590 1485 624 1519
rect 680 1485 714 1519
rect 770 1485 804 1519
rect 866 1462 900 1496
rect -321 1372 -287 1406
rect -321 1282 -287 1316
rect -321 1192 -287 1226
rect -321 1102 -287 1136
rect -321 1012 -287 1046
rect -321 922 -287 956
rect -321 832 -287 866
rect -321 742 -287 776
rect -321 652 -287 686
rect -321 562 -287 596
rect -321 472 -287 506
rect 866 1372 900 1406
rect 866 1282 900 1316
rect 866 1192 900 1226
rect 866 1102 900 1136
rect 866 1012 900 1046
rect 866 922 900 956
rect 866 832 900 866
rect 866 742 900 776
rect 866 652 900 686
rect 866 562 900 596
rect 866 472 900 506
rect -321 382 -287 416
rect 866 382 900 416
rect -220 298 -186 332
rect -130 298 -96 332
rect -40 298 -6 332
rect 50 298 84 332
rect 140 298 174 332
rect 230 298 264 332
rect 320 298 354 332
rect 410 298 444 332
rect 500 298 534 332
rect 590 298 624 332
rect 680 298 714 332
rect 770 298 804 332
rect 1039 1462 1073 1496
rect 1140 1485 1174 1519
rect 1230 1485 1264 1519
rect 1320 1485 1354 1519
rect 1410 1485 1444 1519
rect 1500 1485 1534 1519
rect 1590 1485 1624 1519
rect 1680 1485 1714 1519
rect 1770 1485 1804 1519
rect 1860 1485 1894 1519
rect 1950 1485 1984 1519
rect 2040 1485 2074 1519
rect 2130 1485 2164 1519
rect 2226 1462 2260 1496
rect 1039 1372 1073 1406
rect 1039 1282 1073 1316
rect 1039 1192 1073 1226
rect 1039 1102 1073 1136
rect 1039 1012 1073 1046
rect 1039 922 1073 956
rect 1039 832 1073 866
rect 1039 742 1073 776
rect 1039 652 1073 686
rect 1039 562 1073 596
rect 1039 472 1073 506
rect 2226 1372 2260 1406
rect 2226 1282 2260 1316
rect 2226 1192 2260 1226
rect 2226 1102 2260 1136
rect 2226 1012 2260 1046
rect 2226 922 2260 956
rect 2226 832 2260 866
rect 2226 742 2260 776
rect 2226 652 2260 686
rect 2226 562 2260 596
rect 2226 472 2260 506
rect 1039 382 1073 416
rect 2226 382 2260 416
rect 1140 298 1174 332
rect 1230 298 1264 332
rect 1320 298 1354 332
rect 1410 298 1444 332
rect 1500 298 1534 332
rect 1590 298 1624 332
rect 1680 298 1714 332
rect 1770 298 1804 332
rect 1860 298 1894 332
rect 1950 298 1984 332
rect 2040 298 2074 332
rect 2130 298 2164 332
rect -1681 102 -1647 136
rect -1580 125 -1546 159
rect -1490 125 -1456 159
rect -1400 125 -1366 159
rect -1310 125 -1276 159
rect -1220 125 -1186 159
rect -1130 125 -1096 159
rect -1040 125 -1006 159
rect -950 125 -916 159
rect -860 125 -826 159
rect -770 125 -736 159
rect -680 125 -646 159
rect -590 125 -556 159
rect -494 102 -460 136
rect -1681 12 -1647 46
rect -1681 -78 -1647 -44
rect -3020 -1430 -2980 -1390
rect -1681 -168 -1647 -134
rect -1681 -258 -1647 -224
rect -1681 -348 -1647 -314
rect -1681 -438 -1647 -404
rect -1681 -528 -1647 -494
rect -1681 -618 -1647 -584
rect -1681 -708 -1647 -674
rect -1681 -798 -1647 -764
rect -1681 -888 -1647 -854
rect -494 12 -460 46
rect -494 -78 -460 -44
rect -494 -168 -460 -134
rect -494 -258 -460 -224
rect -494 -348 -460 -314
rect -494 -438 -460 -404
rect -494 -528 -460 -494
rect -494 -618 -460 -584
rect -494 -708 -460 -674
rect -494 -798 -460 -764
rect -494 -888 -460 -854
rect -1681 -978 -1647 -944
rect -494 -978 -460 -944
rect -1580 -1062 -1546 -1028
rect -1490 -1062 -1456 -1028
rect -1400 -1062 -1366 -1028
rect -1310 -1062 -1276 -1028
rect -1220 -1062 -1186 -1028
rect -1130 -1062 -1096 -1028
rect -1040 -1062 -1006 -1028
rect -950 -1062 -916 -1028
rect -860 -1062 -826 -1028
rect -770 -1062 -736 -1028
rect -680 -1062 -646 -1028
rect -590 -1062 -556 -1028
rect -321 102 -287 136
rect -220 125 -186 159
rect -130 125 -96 159
rect -40 125 -6 159
rect 50 125 84 159
rect 140 125 174 159
rect 230 125 264 159
rect 320 125 354 159
rect 410 125 444 159
rect 500 125 534 159
rect 590 125 624 159
rect 680 125 714 159
rect 770 125 804 159
rect 866 102 900 136
rect -321 12 -287 46
rect -321 -78 -287 -44
rect -321 -168 -287 -134
rect -321 -258 -287 -224
rect -321 -348 -287 -314
rect -321 -438 -287 -404
rect -321 -528 -287 -494
rect -321 -618 -287 -584
rect -321 -708 -287 -674
rect -321 -798 -287 -764
rect -321 -888 -287 -854
rect 866 12 900 46
rect 866 -78 900 -44
rect 866 -168 900 -134
rect 866 -258 900 -224
rect 866 -348 900 -314
rect 866 -438 900 -404
rect 866 -528 900 -494
rect 866 -618 900 -584
rect 866 -708 900 -674
rect 866 -798 900 -764
rect 866 -888 900 -854
rect -321 -978 -287 -944
rect 866 -978 900 -944
rect -220 -1062 -186 -1028
rect -130 -1062 -96 -1028
rect -40 -1062 -6 -1028
rect 50 -1062 84 -1028
rect 140 -1062 174 -1028
rect 230 -1062 264 -1028
rect 320 -1062 354 -1028
rect 410 -1062 444 -1028
rect 500 -1062 534 -1028
rect 590 -1062 624 -1028
rect 680 -1062 714 -1028
rect 770 -1062 804 -1028
rect 1039 102 1073 136
rect 1140 125 1174 159
rect 1230 125 1264 159
rect 1320 125 1354 159
rect 1410 125 1444 159
rect 1500 125 1534 159
rect 1590 125 1624 159
rect 1680 125 1714 159
rect 1770 125 1804 159
rect 1860 125 1894 159
rect 1950 125 1984 159
rect 2040 125 2074 159
rect 2130 125 2164 159
rect 2226 102 2260 136
rect 1039 12 1073 46
rect 1039 -78 1073 -44
rect 1039 -168 1073 -134
rect 1039 -258 1073 -224
rect 1039 -348 1073 -314
rect 1039 -438 1073 -404
rect 1039 -528 1073 -494
rect 1039 -618 1073 -584
rect 1039 -708 1073 -674
rect 1039 -798 1073 -764
rect 1039 -888 1073 -854
rect 2226 12 2260 46
rect 2226 -78 2260 -44
rect 2226 -168 2260 -134
rect 2226 -258 2260 -224
rect 2226 -348 2260 -314
rect 2226 -438 2260 -404
rect 2226 -528 2260 -494
rect 2226 -618 2260 -584
rect 2226 -708 2260 -674
rect 2226 -798 2260 -764
rect 2226 -888 2260 -854
rect 1039 -978 1073 -944
rect 2226 -978 2260 -944
rect 1140 -1062 1174 -1028
rect 1230 -1062 1264 -1028
rect 1320 -1062 1354 -1028
rect 1410 -1062 1444 -1028
rect 1500 -1062 1534 -1028
rect 1590 -1062 1624 -1028
rect 1680 -1062 1714 -1028
rect 1770 -1062 1804 -1028
rect 1860 -1062 1894 -1028
rect 1950 -1062 1984 -1028
rect 2040 -1062 2074 -1028
rect 2130 -1062 2164 -1028
rect -1681 -1258 -1647 -1224
rect -1580 -1235 -1546 -1201
rect -1490 -1235 -1456 -1201
rect -1400 -1235 -1366 -1201
rect -1310 -1235 -1276 -1201
rect -1220 -1235 -1186 -1201
rect -1130 -1235 -1096 -1201
rect -1040 -1235 -1006 -1201
rect -950 -1235 -916 -1201
rect -860 -1235 -826 -1201
rect -770 -1235 -736 -1201
rect -680 -1235 -646 -1201
rect -590 -1235 -556 -1201
rect -494 -1258 -460 -1224
rect -1681 -1348 -1647 -1314
rect -1681 -1438 -1647 -1404
rect -1681 -1528 -1647 -1494
rect -1681 -1618 -1647 -1584
rect -1681 -1708 -1647 -1674
rect -1681 -1798 -1647 -1764
rect -1681 -1888 -1647 -1854
rect -1681 -1978 -1647 -1944
rect -1681 -2068 -1647 -2034
rect -1681 -2158 -1647 -2124
rect -1681 -2248 -1647 -2214
rect -494 -1348 -460 -1314
rect -494 -1438 -460 -1404
rect -494 -1528 -460 -1494
rect -494 -1618 -460 -1584
rect -494 -1708 -460 -1674
rect -494 -1798 -460 -1764
rect -494 -1888 -460 -1854
rect -494 -1978 -460 -1944
rect -494 -2068 -460 -2034
rect -494 -2158 -460 -2124
rect -494 -2248 -460 -2214
rect -1681 -2338 -1647 -2304
rect -494 -2338 -460 -2304
rect -1580 -2422 -1546 -2388
rect -1490 -2422 -1456 -2388
rect -1400 -2422 -1366 -2388
rect -1310 -2422 -1276 -2388
rect -1220 -2422 -1186 -2388
rect -1130 -2422 -1096 -2388
rect -1040 -2422 -1006 -2388
rect -950 -2422 -916 -2388
rect -860 -2422 -826 -2388
rect -770 -2422 -736 -2388
rect -680 -2422 -646 -2388
rect -590 -2422 -556 -2388
rect -321 -1258 -287 -1224
rect -220 -1235 -186 -1201
rect -130 -1235 -96 -1201
rect -40 -1235 -6 -1201
rect 50 -1235 84 -1201
rect 140 -1235 174 -1201
rect 230 -1235 264 -1201
rect 320 -1235 354 -1201
rect 410 -1235 444 -1201
rect 500 -1235 534 -1201
rect 590 -1235 624 -1201
rect 680 -1235 714 -1201
rect 770 -1235 804 -1201
rect 866 -1258 900 -1224
rect -321 -1348 -287 -1314
rect -321 -1438 -287 -1404
rect -321 -1528 -287 -1494
rect -321 -1618 -287 -1584
rect -321 -1708 -287 -1674
rect -321 -1798 -287 -1764
rect -321 -1888 -287 -1854
rect -321 -1978 -287 -1944
rect -321 -2068 -287 -2034
rect -321 -2158 -287 -2124
rect -321 -2248 -287 -2214
rect 866 -1348 900 -1314
rect 866 -1438 900 -1404
rect 866 -1528 900 -1494
rect 866 -1618 900 -1584
rect 866 -1708 900 -1674
rect 866 -1798 900 -1764
rect 866 -1888 900 -1854
rect 866 -1978 900 -1944
rect 866 -2068 900 -2034
rect 866 -2158 900 -2124
rect 866 -2248 900 -2214
rect -321 -2338 -287 -2304
rect 866 -2338 900 -2304
rect -220 -2422 -186 -2388
rect -130 -2422 -96 -2388
rect -40 -2422 -6 -2388
rect 50 -2422 84 -2388
rect 140 -2422 174 -2388
rect 230 -2422 264 -2388
rect 320 -2422 354 -2388
rect 410 -2422 444 -2388
rect 500 -2422 534 -2388
rect 590 -2422 624 -2388
rect 680 -2422 714 -2388
rect 770 -2422 804 -2388
rect 1039 -1258 1073 -1224
rect 1140 -1235 1174 -1201
rect 1230 -1235 1264 -1201
rect 1320 -1235 1354 -1201
rect 1410 -1235 1444 -1201
rect 1500 -1235 1534 -1201
rect 1590 -1235 1624 -1201
rect 1680 -1235 1714 -1201
rect 1770 -1235 1804 -1201
rect 1860 -1235 1894 -1201
rect 1950 -1235 1984 -1201
rect 2040 -1235 2074 -1201
rect 2130 -1235 2164 -1201
rect 2226 -1258 2260 -1224
rect 1039 -1348 1073 -1314
rect 1039 -1438 1073 -1404
rect 1039 -1528 1073 -1494
rect 1039 -1618 1073 -1584
rect 1039 -1708 1073 -1674
rect 1039 -1798 1073 -1764
rect 1039 -1888 1073 -1854
rect 1039 -1978 1073 -1944
rect 1039 -2068 1073 -2034
rect 1039 -2158 1073 -2124
rect 1039 -2248 1073 -2214
rect 2226 -1348 2260 -1314
rect 2226 -1438 2260 -1404
rect 2226 -1528 2260 -1494
rect 2226 -1618 2260 -1584
rect 2226 -1708 2260 -1674
rect 2226 -1798 2260 -1764
rect 2226 -1888 2260 -1854
rect 2226 -1978 2260 -1944
rect 2226 -2068 2260 -2034
rect 2226 -2158 2260 -2124
rect 3010 -1490 3050 -1450
rect 2226 -2248 2260 -2214
rect 1039 -2338 1073 -2304
rect 2226 -2338 2260 -2304
rect 1140 -2422 1174 -2388
rect 1230 -2422 1264 -2388
rect 1320 -2422 1354 -2388
rect 1410 -2422 1444 -2388
rect 1500 -2422 1534 -2388
rect 1590 -2422 1624 -2388
rect 1680 -2422 1714 -2388
rect 1770 -2422 1804 -2388
rect 1860 -2422 1894 -2388
rect 1950 -2422 1984 -2388
rect 2040 -2422 2074 -2388
rect 2130 -2422 2164 -2388
rect 270 -2580 310 -2540
rect 270 -2660 310 -2620
rect 270 -2740 310 -2700
<< nsubdiffcont >>
rect -1090 12450 -1050 12490
rect 1280 12450 1320 12490
rect 10210 12530 10370 12570
rect 4150 12450 4190 12490
rect 5450 12450 5490 12490
rect 6750 12450 6790 12490
rect 8050 12450 8090 12490
rect 9200 11270 9240 11600
rect 11380 11270 11420 11600
rect 10210 10800 10370 10840
rect 11250 10800 11320 10840
rect -700 9750 -660 9790
rect -700 9650 -660 9690
rect -700 9550 -660 9590
rect -700 9450 -660 9490
rect 200 9750 240 9790
rect 200 9650 240 9690
rect 200 9550 240 9590
rect 200 9450 240 9490
rect 1100 9750 1140 9790
rect 1100 9650 1140 9690
rect 1100 9550 1140 9590
rect 1100 9450 1140 9490
rect 1240 9750 1280 9790
rect 1240 9650 1280 9690
rect 1240 9550 1280 9590
rect 1240 9450 1280 9490
rect 1680 9750 1720 9790
rect 1680 9650 1720 9690
rect 1680 9550 1720 9590
rect 1680 9450 1720 9490
rect 2010 9750 2050 9790
rect 2010 9650 2050 9690
rect 2010 9550 2050 9590
rect 2010 9450 2050 9490
rect 2420 9750 2460 9790
rect 2420 9650 2460 9690
rect 2420 9550 2460 9590
rect 2420 9450 2460 9490
rect 2810 9750 2850 9790
rect 2810 9650 2850 9690
rect 2810 9550 2850 9590
rect 2810 9450 2850 9490
rect 3200 9750 3240 9790
rect 3200 9650 3240 9690
rect 3200 9550 3240 9590
rect 3200 9450 3240 9490
rect 3880 9750 3920 9790
rect 3880 9650 3920 9690
rect 3880 9550 3920 9590
rect 3880 9450 3920 9490
rect 5570 9720 5610 9760
rect 5570 9620 5610 9660
rect 5570 9520 5610 9560
rect 5570 9420 5610 9460
rect 7090 9720 7130 9760
rect 7090 9620 7130 9660
rect 7090 9520 7130 9560
rect 7090 9420 7130 9460
rect 8610 9720 8650 9760
rect 8610 9620 8650 9660
rect 8610 9520 8650 9560
rect 8610 9420 8650 9460
rect -700 8990 -660 9030
rect -700 8890 -660 8930
rect -700 8790 -660 8830
rect -700 8690 -660 8730
rect 200 8990 240 9030
rect 200 8890 240 8930
rect 200 8790 240 8830
rect 200 8690 240 8730
rect 1100 8990 1140 9030
rect 1100 8890 1140 8930
rect 1100 8790 1140 8830
rect 1100 8690 1140 8730
rect 1500 8990 1540 9030
rect 1500 8890 1540 8930
rect 1500 8790 1540 8830
rect 1500 8690 1540 8730
rect 1830 8990 1870 9030
rect 1830 8890 1870 8930
rect 1830 8790 1870 8830
rect 1830 8690 1870 8730
rect 2160 8990 2200 9030
rect 2160 8890 2200 8930
rect 2160 8790 2200 8830
rect 2160 8690 2200 8730
rect 2420 8990 2460 9030
rect 2420 8890 2460 8930
rect 2420 8790 2460 8830
rect 2420 8690 2460 8730
rect 3200 8990 3240 9030
rect 3200 8890 3240 8930
rect 3200 8790 3240 8830
rect 3200 8690 3240 8730
rect -1420 6800 -1380 6840
rect -1420 6700 -1380 6740
rect 60 6800 100 6840
rect 60 6700 100 6740
rect 480 6800 520 6840
rect 480 6700 520 6740
rect 1960 6800 2000 6840
rect 1960 6700 2000 6740
rect -1430 6200 -1390 6240
rect -1430 6100 -1390 6140
rect -1430 6000 -1390 6040
rect -1430 5900 -1390 5940
rect -1430 5800 -1390 5840
rect -1430 5700 -1390 5740
rect 1970 6200 2010 6240
rect 1970 6100 2010 6140
rect 1970 6000 2010 6040
rect 1970 5900 2010 5940
rect 2430 6000 2470 6040
rect 2430 5900 2470 5940
rect 3040 6000 3080 6040
rect 3040 5900 3080 5940
rect 1970 5800 2010 5840
rect 1970 5700 2010 5740
rect -2530 4640 -2490 4680
rect -2530 4540 -2490 4580
rect 30 4640 70 4680
rect 30 4540 70 4580
rect 510 4640 550 4680
rect 510 4540 550 4580
rect 3070 4640 3110 4680
rect 6620 4720 6660 4760
rect 6620 4620 6660 4660
rect 7600 4720 7640 4760
rect 7600 4620 7640 4660
rect 7760 4720 7800 4760
rect 7760 4620 7800 4660
rect 8740 4720 8780 4760
rect 8740 4620 8780 4660
rect 3070 4540 3110 4580
rect 5550 4070 5590 4110
rect 5550 3970 5590 4010
rect 5550 3870 5590 3910
rect 5550 3770 5590 3810
rect 5550 3670 5590 3710
rect 7750 4070 7790 4110
rect 7750 3970 7790 4010
rect 7750 3870 7790 3910
rect 7750 3770 7790 3810
rect 7750 3670 7790 3710
rect -1474 1338 -1440 1372
rect -1384 1338 -1350 1372
rect -1294 1338 -1260 1372
rect -1204 1338 -1170 1372
rect -1114 1338 -1080 1372
rect -1024 1338 -990 1372
rect -934 1338 -900 1372
rect -844 1338 -810 1372
rect -754 1338 -720 1372
rect -1532 1262 -1498 1296
rect -642 1281 -608 1315
rect -1532 1172 -1498 1206
rect -1532 1082 -1498 1116
rect -1532 992 -1498 1026
rect -1532 902 -1498 936
rect -1532 812 -1498 846
rect -1532 722 -1498 756
rect -1532 632 -1498 666
rect -1532 542 -1498 576
rect -642 1191 -608 1225
rect -642 1101 -608 1135
rect -642 1011 -608 1045
rect -642 921 -608 955
rect -642 831 -608 865
rect -642 741 -608 775
rect -642 651 -608 685
rect -642 561 -608 595
rect -1440 448 -1406 482
rect -1350 448 -1316 482
rect -1260 448 -1226 482
rect -1170 448 -1136 482
rect -1080 448 -1046 482
rect -990 448 -956 482
rect -900 448 -866 482
rect -810 448 -776 482
rect -720 448 -686 482
rect -114 1338 -80 1372
rect -24 1338 10 1372
rect 66 1338 100 1372
rect 156 1338 190 1372
rect 246 1338 280 1372
rect 336 1338 370 1372
rect 426 1338 460 1372
rect 516 1338 550 1372
rect 606 1338 640 1372
rect -172 1262 -138 1296
rect 718 1281 752 1315
rect -172 1172 -138 1206
rect -172 1082 -138 1116
rect -172 992 -138 1026
rect -172 902 -138 936
rect -172 812 -138 846
rect -172 722 -138 756
rect -172 632 -138 666
rect -172 542 -138 576
rect 718 1191 752 1225
rect 718 1101 752 1135
rect 718 1011 752 1045
rect 718 921 752 955
rect 718 831 752 865
rect 718 741 752 775
rect 718 651 752 685
rect 718 561 752 595
rect -80 448 -46 482
rect 10 448 44 482
rect 100 448 134 482
rect 190 448 224 482
rect 280 448 314 482
rect 370 448 404 482
rect 460 448 494 482
rect 550 448 584 482
rect 640 448 674 482
rect 1246 1338 1280 1372
rect 1336 1338 1370 1372
rect 1426 1338 1460 1372
rect 1516 1338 1550 1372
rect 1606 1338 1640 1372
rect 1696 1338 1730 1372
rect 1786 1338 1820 1372
rect 1876 1338 1910 1372
rect 1966 1338 2000 1372
rect 1188 1262 1222 1296
rect 2078 1281 2112 1315
rect 1188 1172 1222 1206
rect 1188 1082 1222 1116
rect 1188 992 1222 1026
rect 1188 902 1222 936
rect 1188 812 1222 846
rect 1188 722 1222 756
rect 1188 632 1222 666
rect 1188 542 1222 576
rect 2078 1191 2112 1225
rect 2078 1101 2112 1135
rect 2078 1011 2112 1045
rect 2078 921 2112 955
rect 2078 831 2112 865
rect 2078 741 2112 775
rect 2078 651 2112 685
rect 2078 561 2112 595
rect 1280 448 1314 482
rect 1370 448 1404 482
rect 1460 448 1494 482
rect 1550 448 1584 482
rect 1640 448 1674 482
rect 1730 448 1764 482
rect 1820 448 1854 482
rect 1910 448 1944 482
rect 2000 448 2034 482
rect -1474 -22 -1440 12
rect -1384 -22 -1350 12
rect -1294 -22 -1260 12
rect -1204 -22 -1170 12
rect -1114 -22 -1080 12
rect -1024 -22 -990 12
rect -934 -22 -900 12
rect -844 -22 -810 12
rect -754 -22 -720 12
rect -1532 -98 -1498 -64
rect -642 -79 -608 -45
rect -1532 -188 -1498 -154
rect -1532 -278 -1498 -244
rect -1532 -368 -1498 -334
rect -1532 -458 -1498 -424
rect -1532 -548 -1498 -514
rect -1532 -638 -1498 -604
rect -1532 -728 -1498 -694
rect -1532 -818 -1498 -784
rect -642 -169 -608 -135
rect -642 -259 -608 -225
rect -642 -349 -608 -315
rect -642 -439 -608 -405
rect -642 -529 -608 -495
rect -642 -619 -608 -585
rect -642 -709 -608 -675
rect -642 -799 -608 -765
rect -1440 -912 -1406 -878
rect -1350 -912 -1316 -878
rect -1260 -912 -1226 -878
rect -1170 -912 -1136 -878
rect -1080 -912 -1046 -878
rect -990 -912 -956 -878
rect -900 -912 -866 -878
rect -810 -912 -776 -878
rect -720 -912 -686 -878
rect -114 -22 -80 12
rect -24 -22 10 12
rect 66 -22 100 12
rect 156 -22 190 12
rect 246 -22 280 12
rect 336 -22 370 12
rect 426 -22 460 12
rect 516 -22 550 12
rect 606 -22 640 12
rect -172 -98 -138 -64
rect 718 -79 752 -45
rect -172 -188 -138 -154
rect -172 -278 -138 -244
rect -172 -368 -138 -334
rect -172 -458 -138 -424
rect -172 -548 -138 -514
rect -172 -638 -138 -604
rect -172 -728 -138 -694
rect -172 -818 -138 -784
rect 718 -169 752 -135
rect 718 -259 752 -225
rect 718 -349 752 -315
rect 718 -439 752 -405
rect 718 -529 752 -495
rect 718 -619 752 -585
rect 718 -709 752 -675
rect 718 -799 752 -765
rect -80 -912 -46 -878
rect 10 -912 44 -878
rect 100 -912 134 -878
rect 190 -912 224 -878
rect 280 -912 314 -878
rect 370 -912 404 -878
rect 460 -912 494 -878
rect 550 -912 584 -878
rect 640 -912 674 -878
rect 1246 -22 1280 12
rect 1336 -22 1370 12
rect 1426 -22 1460 12
rect 1516 -22 1550 12
rect 1606 -22 1640 12
rect 1696 -22 1730 12
rect 1786 -22 1820 12
rect 1876 -22 1910 12
rect 1966 -22 2000 12
rect 1188 -98 1222 -64
rect 2078 -79 2112 -45
rect 1188 -188 1222 -154
rect 1188 -278 1222 -244
rect 1188 -368 1222 -334
rect 1188 -458 1222 -424
rect 1188 -548 1222 -514
rect 1188 -638 1222 -604
rect 1188 -728 1222 -694
rect 1188 -818 1222 -784
rect 2078 -169 2112 -135
rect 2078 -259 2112 -225
rect 2078 -349 2112 -315
rect 2078 -439 2112 -405
rect 2078 -529 2112 -495
rect 2078 -619 2112 -585
rect 2078 -709 2112 -675
rect 2078 -799 2112 -765
rect 1280 -912 1314 -878
rect 1370 -912 1404 -878
rect 1460 -912 1494 -878
rect 1550 -912 1584 -878
rect 1640 -912 1674 -878
rect 1730 -912 1764 -878
rect 1820 -912 1854 -878
rect 1910 -912 1944 -878
rect 2000 -912 2034 -878
rect -1474 -1382 -1440 -1348
rect -1384 -1382 -1350 -1348
rect -1294 -1382 -1260 -1348
rect -1204 -1382 -1170 -1348
rect -1114 -1382 -1080 -1348
rect -1024 -1382 -990 -1348
rect -934 -1382 -900 -1348
rect -844 -1382 -810 -1348
rect -754 -1382 -720 -1348
rect -1532 -1458 -1498 -1424
rect -642 -1439 -608 -1405
rect -1532 -1548 -1498 -1514
rect -1532 -1638 -1498 -1604
rect -1532 -1728 -1498 -1694
rect -1532 -1818 -1498 -1784
rect -1532 -1908 -1498 -1874
rect -1532 -1998 -1498 -1964
rect -1532 -2088 -1498 -2054
rect -1532 -2178 -1498 -2144
rect -642 -1529 -608 -1495
rect -642 -1619 -608 -1585
rect -642 -1709 -608 -1675
rect -642 -1799 -608 -1765
rect -642 -1889 -608 -1855
rect -642 -1979 -608 -1945
rect -642 -2069 -608 -2035
rect -642 -2159 -608 -2125
rect -1440 -2272 -1406 -2238
rect -1350 -2272 -1316 -2238
rect -1260 -2272 -1226 -2238
rect -1170 -2272 -1136 -2238
rect -1080 -2272 -1046 -2238
rect -990 -2272 -956 -2238
rect -900 -2272 -866 -2238
rect -810 -2272 -776 -2238
rect -720 -2272 -686 -2238
rect -114 -1382 -80 -1348
rect -24 -1382 10 -1348
rect 66 -1382 100 -1348
rect 156 -1382 190 -1348
rect 246 -1382 280 -1348
rect 336 -1382 370 -1348
rect 426 -1382 460 -1348
rect 516 -1382 550 -1348
rect 606 -1382 640 -1348
rect -172 -1458 -138 -1424
rect 718 -1439 752 -1405
rect -172 -1548 -138 -1514
rect -172 -1638 -138 -1604
rect -172 -1728 -138 -1694
rect -172 -1818 -138 -1784
rect -172 -1908 -138 -1874
rect -172 -1998 -138 -1964
rect -172 -2088 -138 -2054
rect -172 -2178 -138 -2144
rect 718 -1529 752 -1495
rect 718 -1619 752 -1585
rect 718 -1709 752 -1675
rect 718 -1799 752 -1765
rect 718 -1889 752 -1855
rect 718 -1979 752 -1945
rect 718 -2069 752 -2035
rect 718 -2159 752 -2125
rect -80 -2272 -46 -2238
rect 10 -2272 44 -2238
rect 100 -2272 134 -2238
rect 190 -2272 224 -2238
rect 280 -2272 314 -2238
rect 370 -2272 404 -2238
rect 460 -2272 494 -2238
rect 550 -2272 584 -2238
rect 640 -2272 674 -2238
rect 1246 -1382 1280 -1348
rect 1336 -1382 1370 -1348
rect 1426 -1382 1460 -1348
rect 1516 -1382 1550 -1348
rect 1606 -1382 1640 -1348
rect 1696 -1382 1730 -1348
rect 1786 -1382 1820 -1348
rect 1876 -1382 1910 -1348
rect 1966 -1382 2000 -1348
rect 1188 -1458 1222 -1424
rect 2078 -1439 2112 -1405
rect 1188 -1548 1222 -1514
rect 1188 -1638 1222 -1604
rect 1188 -1728 1222 -1694
rect 1188 -1818 1222 -1784
rect 1188 -1908 1222 -1874
rect 1188 -1998 1222 -1964
rect 1188 -2088 1222 -2054
rect 1188 -2178 1222 -2144
rect 2078 -1529 2112 -1495
rect 2078 -1619 2112 -1585
rect 2078 -1709 2112 -1675
rect 2078 -1799 2112 -1765
rect 2078 -1889 2112 -1855
rect 2078 -1979 2112 -1945
rect 2078 -2069 2112 -2035
rect 2078 -2159 2112 -2125
rect 1280 -2272 1314 -2238
rect 1370 -2272 1404 -2238
rect 1460 -2272 1494 -2238
rect 1550 -2272 1584 -2238
rect 1640 -2272 1674 -2238
rect 1730 -2272 1764 -2238
rect 1820 -2272 1854 -2238
rect 1910 -2272 1944 -2238
rect 2000 -2272 2034 -2238
<< poly >>
rect 9380 13790 9410 13820
rect 9900 13790 9930 13820
rect 10420 13790 10450 13820
rect 11020 13790 11050 13820
rect 9380 13560 9410 13590
rect 9900 13560 9930 13590
rect 10420 13560 10450 13590
rect 11020 13560 11050 13590
rect 9366 13542 9424 13560
rect 9366 13508 9378 13542
rect 9412 13508 9424 13542
rect 9366 13490 9424 13508
rect 9886 13542 9944 13560
rect 9886 13508 9898 13542
rect 9932 13508 9944 13542
rect 9886 13490 9944 13508
rect 10406 13542 10464 13560
rect 10406 13508 10418 13542
rect 10452 13508 10464 13542
rect 10406 13490 10464 13508
rect 10974 13542 11050 13560
rect 10974 13508 10986 13542
rect 11020 13508 11050 13542
rect 10974 13490 11050 13508
rect 9380 13410 9410 13440
rect 9900 13410 9930 13440
rect 10420 13410 10450 13440
rect -1510 12930 -1430 12950
rect -1510 12890 -1490 12930
rect -1450 12890 -1430 12930
rect -1510 12870 -1430 12890
rect -560 12910 -480 12930
rect -560 12870 -540 12910
rect -500 12870 -480 12910
rect 510 12920 590 12940
rect 510 12880 530 12920
rect 570 12880 590 12920
rect 510 12870 590 12880
rect 2070 12920 2160 12940
rect 2070 12880 2090 12920
rect 2130 12880 2160 12920
rect 2070 12870 2160 12880
rect 4684 12930 4750 12950
rect 5250 12930 5280 12960
rect 5360 12930 5390 12960
rect 5470 12930 5500 12960
rect 5580 12930 5610 12960
rect 5910 12930 5940 12960
rect 6020 12930 6050 12960
rect 6130 12930 6160 12960
rect 6550 12930 6580 12960
rect 6660 12930 6690 12960
rect 6770 12930 6800 12960
rect 6880 12930 6910 12960
rect 7210 12930 7240 12960
rect 7320 12930 7350 12960
rect 7430 12930 7460 12960
rect 7850 12930 7880 12960
rect 7960 12930 7990 12960
rect 8070 12930 8100 12960
rect 8180 12930 8210 12960
rect 8510 12930 8540 12960
rect 8620 12930 8650 12960
rect 8730 12930 8760 12960
rect 4684 12890 4694 12930
rect 4734 12890 4750 12930
rect 4684 12870 4750 12890
rect -1380 12840 -1350 12870
rect -1270 12840 -1240 12870
rect -1160 12840 -1130 12870
rect -1050 12840 -1020 12870
rect -800 12840 -770 12870
rect -690 12840 -660 12870
rect -560 12850 -480 12870
rect -1380 12710 -1350 12740
rect -1270 12720 -1240 12740
rect -1160 12720 -1130 12740
rect -1050 12720 -1020 12740
rect -800 12720 -770 12740
rect -1270 12710 -770 12720
rect -1400 12690 -1320 12710
rect -1270 12690 -740 12710
rect -1400 12650 -1380 12690
rect -1340 12650 -1320 12690
rect -1400 12630 -1320 12650
rect -1220 12520 -1190 12690
rect -820 12650 -800 12690
rect -760 12650 -740 12690
rect -820 12630 -740 12650
rect -690 12610 -660 12740
rect -560 12610 -530 12850
rect -350 12840 -320 12870
rect -240 12840 -210 12870
rect -130 12840 -100 12870
rect -20 12840 10 12870
rect 310 12840 340 12870
rect 420 12840 450 12870
rect 530 12840 560 12870
rect 640 12840 670 12870
rect 990 12840 1020 12870
rect 1100 12840 1130 12870
rect 1210 12840 1240 12870
rect 1320 12840 1350 12870
rect 1570 12840 1600 12870
rect 1680 12840 1710 12870
rect 2130 12840 2160 12870
rect 2490 12840 2520 12870
rect 2740 12840 2770 12870
rect 2850 12840 2880 12870
rect 2960 12840 2990 12870
rect 3070 12840 3100 12870
rect 3400 12840 3430 12870
rect 3510 12840 3540 12870
rect 3620 12840 3650 12870
rect 3950 12840 3980 12870
rect 4060 12840 4090 12870
rect 4170 12840 4200 12870
rect 4280 12840 4310 12870
rect 4610 12840 4640 12870
rect 4720 12840 4750 12870
rect 4830 12840 4860 12870
rect 5250 12800 5280 12830
rect 5360 12810 5390 12830
rect 5470 12810 5500 12830
rect 5580 12810 5610 12830
rect 5910 12810 5940 12830
rect 5230 12780 5310 12800
rect 5230 12740 5250 12780
rect 5290 12740 5310 12780
rect -480 12690 -400 12710
rect -480 12650 -460 12690
rect -420 12650 -400 12690
rect -480 12630 -400 12650
rect -350 12630 -320 12740
rect -240 12710 -210 12740
rect -130 12710 -100 12740
rect -20 12710 10 12740
rect -240 12690 180 12710
rect -240 12680 120 12690
rect -690 12580 -530 12610
rect -350 12610 -200 12630
rect -350 12600 -260 12610
rect -800 12520 -770 12550
rect -690 12520 -660 12580
rect -1530 12490 -1450 12510
rect -1530 12450 -1510 12490
rect -1470 12450 -1450 12490
rect -1530 12430 -1450 12450
rect -1220 12390 -1190 12420
rect -800 12390 -770 12420
rect -690 12390 -660 12420
rect -560 12410 -530 12580
rect -280 12570 -260 12600
rect -220 12570 -200 12610
rect -280 12550 -200 12570
rect -130 12520 -100 12680
rect 100 12650 120 12680
rect 160 12650 180 12690
rect 100 12640 180 12650
rect 120 12580 200 12590
rect -20 12570 200 12580
rect -20 12550 140 12570
rect -20 12520 10 12550
rect 120 12530 140 12550
rect 180 12530 200 12570
rect 120 12510 200 12530
rect 310 12520 340 12740
rect 420 12520 450 12740
rect 530 12520 560 12740
rect 640 12710 670 12740
rect 990 12710 1020 12740
rect 1100 12720 1130 12740
rect 1210 12720 1240 12740
rect 1320 12720 1350 12740
rect 1570 12720 1600 12740
rect 1100 12710 1600 12720
rect 620 12690 850 12710
rect 620 12650 640 12690
rect 680 12680 850 12690
rect 680 12650 700 12680
rect 620 12640 700 12650
rect 820 12590 850 12680
rect 970 12690 1050 12710
rect 1100 12690 1630 12710
rect 970 12650 990 12690
rect 1030 12650 1050 12690
rect 970 12640 1050 12650
rect 1150 12590 1180 12690
rect 1550 12650 1570 12690
rect 1610 12650 1630 12690
rect 1550 12630 1630 12650
rect 820 12560 1180 12590
rect 1150 12520 1180 12560
rect 1680 12590 1710 12740
rect 1760 12690 1840 12710
rect 1760 12650 1780 12690
rect 1820 12680 1840 12690
rect 2000 12690 2080 12710
rect 2000 12680 2020 12690
rect 1820 12650 2020 12680
rect 2060 12650 2080 12690
rect 1760 12640 1840 12650
rect 2000 12630 2080 12650
rect 1680 12570 1900 12590
rect 2130 12570 2160 12740
rect 2340 12680 2420 12700
rect 2340 12640 2360 12680
rect 2400 12640 2420 12680
rect 2340 12620 2420 12640
rect 2490 12640 2520 12740
rect 2610 12640 2690 12660
rect 2490 12610 2630 12640
rect 2490 12570 2520 12610
rect 2610 12600 2630 12610
rect 2670 12600 2690 12640
rect 2740 12630 2770 12740
rect 2850 12710 2880 12740
rect 2960 12710 2990 12740
rect 3070 12710 3100 12740
rect 2850 12690 3320 12710
rect 2850 12680 3260 12690
rect 2740 12610 2890 12630
rect 2740 12600 2830 12610
rect 2610 12580 2690 12600
rect 1680 12560 1840 12570
rect 1570 12520 1600 12550
rect 1680 12520 1710 12560
rect 1820 12530 1840 12560
rect 1880 12530 1900 12570
rect 1820 12510 1900 12530
rect 2020 12540 2160 12570
rect 2020 12520 2050 12540
rect 2130 12520 2160 12540
rect 2380 12540 2520 12570
rect 2810 12570 2830 12600
rect 2870 12570 2890 12610
rect 2810 12550 2890 12570
rect 2380 12520 2410 12540
rect 2490 12520 2520 12540
rect 2960 12520 2990 12680
rect 3240 12650 3260 12680
rect 3300 12650 3320 12690
rect 3240 12640 3320 12650
rect 3210 12580 3290 12590
rect 3070 12570 3290 12580
rect 3070 12550 3230 12570
rect 3070 12520 3100 12550
rect 3210 12530 3230 12550
rect 3270 12530 3290 12570
rect 3210 12510 3290 12530
rect 3400 12520 3430 12740
rect 3510 12590 3540 12740
rect 3620 12710 3650 12740
rect 3950 12710 3980 12740
rect 4060 12720 4090 12740
rect 4170 12720 4200 12740
rect 4280 12720 4310 12740
rect 4610 12720 4640 12740
rect 3600 12690 3810 12710
rect 3600 12650 3620 12690
rect 3660 12680 3810 12690
rect 3660 12650 3680 12680
rect 3600 12640 3680 12650
rect 3780 12590 3810 12680
rect 3930 12690 4010 12710
rect 3930 12650 3950 12690
rect 3990 12650 4010 12690
rect 3930 12640 4010 12650
rect 4060 12690 4640 12720
rect 4060 12590 4090 12690
rect 4510 12650 4530 12690
rect 4570 12650 4590 12690
rect 4510 12630 4590 12650
rect 4720 12630 4750 12740
rect 3510 12560 3670 12590
rect 3780 12560 4090 12590
rect 4340 12610 4420 12630
rect 4340 12570 4360 12610
rect 4400 12570 4420 12610
rect 4640 12600 4750 12630
rect 4830 12660 4860 12740
rect 5230 12720 5310 12740
rect 5360 12780 5940 12810
rect 4980 12670 5060 12690
rect 4980 12660 5000 12670
rect 4830 12630 5000 12660
rect 5040 12630 5060 12670
rect 4640 12570 4670 12600
rect 3510 12520 3540 12560
rect 3640 12510 3670 12560
rect 4020 12520 4050 12560
rect 4340 12550 4420 12570
rect 4360 12520 4390 12550
rect 4470 12540 4670 12570
rect 4470 12520 4500 12540
rect 4720 12520 4750 12550
rect 4830 12520 4860 12630
rect 4980 12610 5060 12630
rect 5360 12580 5390 12780
rect 5810 12740 5830 12780
rect 5870 12740 5890 12780
rect 5810 12720 5890 12740
rect 6020 12660 6050 12830
rect 5770 12630 6050 12660
rect 6130 12660 6160 12830
rect 6550 12800 6580 12830
rect 6660 12810 6690 12830
rect 6770 12810 6800 12830
rect 6880 12810 6910 12830
rect 7210 12810 7240 12830
rect 6530 12780 6610 12800
rect 6530 12740 6550 12780
rect 6590 12740 6610 12780
rect 6530 12720 6610 12740
rect 6660 12780 7240 12810
rect 6280 12670 6360 12690
rect 6280 12660 6300 12670
rect 6130 12630 6300 12660
rect 6340 12630 6360 12670
rect 5320 12550 5390 12580
rect 5640 12610 5720 12630
rect 5640 12570 5660 12610
rect 5700 12570 5720 12610
rect 5640 12550 5720 12570
rect 5320 12520 5350 12550
rect 5660 12520 5690 12550
rect 5770 12520 5800 12630
rect 6020 12520 6050 12550
rect 6130 12520 6160 12630
rect 6280 12610 6360 12630
rect 6660 12580 6690 12780
rect 7110 12740 7130 12780
rect 7170 12740 7190 12780
rect 7110 12720 7190 12740
rect 7320 12660 7350 12830
rect 7070 12630 7350 12660
rect 7430 12660 7460 12830
rect 7850 12800 7880 12830
rect 7960 12810 7990 12830
rect 8070 12810 8100 12830
rect 8180 12810 8210 12830
rect 8510 12810 8540 12830
rect 7830 12780 7910 12800
rect 7830 12740 7850 12780
rect 7890 12740 7910 12780
rect 7830 12720 7910 12740
rect 7960 12780 8540 12810
rect 7580 12670 7660 12690
rect 7580 12660 7600 12670
rect 7430 12630 7600 12660
rect 7640 12630 7660 12670
rect 6620 12550 6690 12580
rect 6940 12610 7020 12630
rect 6940 12570 6960 12610
rect 7000 12570 7020 12610
rect 6940 12550 7020 12570
rect 6620 12520 6650 12550
rect 6960 12520 6990 12550
rect 7070 12520 7100 12630
rect 7320 12520 7350 12550
rect 7430 12520 7460 12630
rect 7580 12610 7660 12630
rect 7960 12580 7990 12780
rect 8410 12740 8430 12780
rect 8470 12740 8490 12780
rect 8410 12720 8490 12740
rect 8620 12660 8650 12830
rect 8370 12630 8650 12660
rect 8730 12660 8760 12830
rect 9380 13180 9410 13210
rect 9900 13180 9930 13210
rect 10420 13180 10450 13210
rect 9380 13162 9438 13180
rect 9380 13128 9392 13162
rect 9426 13128 9438 13162
rect 9380 13110 9438 13128
rect 9900 13162 9958 13180
rect 9900 13128 9912 13162
rect 9946 13128 9958 13162
rect 9900 13110 9958 13128
rect 10420 13162 10478 13180
rect 10420 13128 10432 13162
rect 10466 13128 10478 13162
rect 10420 13110 10478 13128
rect 9380 13030 9410 13060
rect 9900 13030 9930 13060
rect 10420 13030 10450 13060
rect 9380 12900 9410 12930
rect 9900 12900 9930 12930
rect 10420 12900 10450 12930
rect 9352 12882 9410 12900
rect 9352 12848 9364 12882
rect 9398 12848 9410 12882
rect 9352 12830 9410 12848
rect 9872 12882 9930 12900
rect 9872 12848 9884 12882
rect 9918 12848 9930 12882
rect 9872 12830 9930 12848
rect 10392 12882 10450 12900
rect 10392 12848 10404 12882
rect 10438 12848 10450 12882
rect 10392 12830 10450 12848
rect 8862 12662 8920 12690
rect 8862 12660 8874 12662
rect 8730 12630 8874 12660
rect 7920 12550 7990 12580
rect 8240 12610 8320 12630
rect 8240 12570 8260 12610
rect 8300 12570 8320 12610
rect 8240 12550 8320 12570
rect 7920 12520 7950 12550
rect 8260 12520 8290 12550
rect 8370 12520 8400 12630
rect 8620 12520 8650 12550
rect 8730 12520 8760 12630
rect 8862 12628 8874 12630
rect 8908 12628 8920 12662
rect 8862 12610 8920 12628
rect 3640 12490 3880 12510
rect 3640 12480 3820 12490
rect 3800 12450 3820 12480
rect 3860 12450 3880 12490
rect 3800 12430 3880 12450
rect -560 12390 -480 12410
rect -130 12390 -100 12420
rect -20 12390 10 12420
rect 310 12390 340 12420
rect 420 12390 450 12420
rect 530 12390 560 12420
rect 1150 12390 1180 12420
rect 1570 12390 1600 12420
rect 1680 12390 1710 12420
rect 2020 12390 2050 12420
rect 2130 12390 2160 12420
rect 2380 12390 2410 12420
rect 2490 12390 2520 12420
rect 2960 12390 2990 12420
rect 3070 12390 3100 12420
rect -870 12370 -770 12390
rect -870 12330 -850 12370
rect -810 12330 -770 12370
rect -560 12350 -540 12390
rect -500 12350 -480 12390
rect -560 12330 -480 12350
rect 250 12370 340 12390
rect 250 12330 270 12370
rect 310 12330 340 12370
rect -870 12310 -770 12330
rect 250 12310 340 12330
rect 390 12370 450 12390
rect 390 12330 400 12370
rect 440 12330 450 12370
rect 390 12310 450 12330
rect 1510 12370 1600 12390
rect 3400 12380 3430 12420
rect 3510 12390 3540 12420
rect 4020 12390 4050 12420
rect 4360 12390 4390 12420
rect 4470 12390 4500 12420
rect 4720 12400 4750 12420
rect 4830 12400 4860 12420
rect 1510 12330 1530 12370
rect 1570 12330 1600 12370
rect 1510 12310 1600 12330
rect 3270 12360 3430 12380
rect 4720 12370 4860 12400
rect 5320 12390 5350 12420
rect 5660 12390 5690 12420
rect 5770 12390 5800 12420
rect 6020 12400 6050 12420
rect 6130 12400 6160 12420
rect 5770 12370 5880 12390
rect 6020 12370 6160 12400
rect 6620 12390 6650 12420
rect 6960 12390 6990 12420
rect 7070 12390 7100 12420
rect 7320 12400 7350 12420
rect 7430 12400 7460 12420
rect 7070 12370 7180 12390
rect 7320 12370 7460 12400
rect 7920 12390 7950 12420
rect 8260 12390 8290 12420
rect 8370 12390 8400 12420
rect 8620 12400 8650 12420
rect 8730 12400 8760 12420
rect 8370 12370 8480 12390
rect 8620 12370 8760 12400
rect 3270 12320 3290 12360
rect 3330 12350 3430 12360
rect 3330 12320 3350 12350
rect 3270 12310 3350 12320
rect 5770 12330 5820 12370
rect 5860 12330 5880 12370
rect 5770 12310 5880 12330
rect 7070 12330 7120 12370
rect 7160 12330 7180 12370
rect 7070 12310 7180 12330
rect 8370 12330 8420 12370
rect 8460 12330 8480 12370
rect 8370 12310 8480 12330
rect 9352 12452 9410 12470
rect 9352 12418 9364 12452
rect 9398 12418 9410 12452
rect 9352 12400 9410 12418
rect 9872 12452 9930 12470
rect 9872 12418 9884 12452
rect 9918 12418 9930 12452
rect 9872 12400 9930 12418
rect 10392 12452 10450 12470
rect 10392 12418 10404 12452
rect 10438 12418 10450 12452
rect 10392 12400 10450 12418
rect 9380 12370 9410 12400
rect 9900 12370 9930 12400
rect 10420 12370 10450 12400
rect 9380 12140 9410 12170
rect 9900 12140 9930 12170
rect 10420 12140 10450 12170
rect 9380 12072 9438 12090
rect 9380 12038 9392 12072
rect 9426 12038 9438 12072
rect 9380 12020 9438 12038
rect 9900 12072 9958 12090
rect 9900 12038 9912 12072
rect 9946 12038 9958 12072
rect 9900 12020 9958 12038
rect 10420 12072 10478 12090
rect 10420 12038 10432 12072
rect 10466 12038 10478 12072
rect 10420 12020 10478 12038
rect 9380 11990 9410 12020
rect 9900 11990 9930 12020
rect 10420 11990 10450 12020
rect 9380 11560 9410 11590
rect 9900 11560 9930 11590
rect 10420 11560 10450 11590
rect 9490 11390 9570 11410
rect 9490 11350 9510 11390
rect 9550 11350 9570 11390
rect 9490 11330 9570 11350
rect 10010 11390 10090 11410
rect 10010 11350 10030 11390
rect 10070 11350 10090 11390
rect 10010 11330 10090 11350
rect 10530 11390 10610 11410
rect 10530 11350 10550 11390
rect 10590 11350 10610 11390
rect 10530 11330 10610 11350
rect 11060 11390 11120 11410
rect 11060 11350 11070 11390
rect 11110 11350 11120 11390
rect 11060 11330 11120 11350
rect 9380 11300 9680 11330
rect 9900 11300 10200 11330
rect 10420 11300 10720 11330
rect 10940 11300 11240 11330
rect 9380 10870 9680 10900
rect 9900 10870 10200 10900
rect 10420 10870 10720 10900
rect 10940 10870 11240 10900
rect -40 10320 370 10350
rect -560 10240 -530 10270
rect -450 10240 -420 10270
rect -40 10240 -10 10320
rect 70 10240 100 10270
rect 340 10240 370 10320
rect 1490 10330 1570 10350
rect 1490 10290 1510 10330
rect 1550 10290 1570 10330
rect 1490 10270 1570 10290
rect 450 10240 480 10270
rect 860 10240 890 10270
rect 970 10240 1000 10270
rect 1380 10240 1410 10270
rect 1490 10240 1520 10270
rect 1820 10240 1850 10270
rect 2150 10240 2180 10270
rect 2590 10240 2620 10270
rect 2980 10240 3010 10270
rect 3370 10240 3400 10270
rect 3660 10240 3690 10270
rect -560 9970 -530 10040
rect -760 9950 -530 9970
rect -760 9910 -740 9950
rect -700 9940 -530 9950
rect -700 9910 -680 9940
rect -760 9890 -680 9910
rect -560 9820 -530 9940
rect -450 10010 -420 10040
rect -450 9990 -350 10010
rect -40 10000 -10 10040
rect -450 9950 -410 9990
rect -370 9950 -350 9990
rect -450 9930 -350 9950
rect -260 9970 -10 10000
rect -450 9820 -420 9930
rect -260 9510 -230 9970
rect -40 9820 -10 9970
rect 70 9930 100 10040
rect 70 9910 170 9930
rect 70 9870 110 9910
rect 150 9870 170 9910
rect 70 9850 170 9870
rect 70 9820 100 9850
rect 340 9820 370 10040
rect 450 10010 480 10040
rect 450 9990 550 10010
rect 860 10000 890 10040
rect 450 9950 490 9990
rect 530 9950 550 9990
rect 450 9930 550 9950
rect 640 9970 890 10000
rect 450 9820 480 9930
rect -310 9490 -230 9510
rect -310 9450 -290 9490
rect -250 9450 -230 9490
rect -310 9430 -230 9450
rect 640 9510 670 9970
rect 860 9820 890 9970
rect 970 10000 1000 10040
rect 970 9980 1220 10000
rect 970 9970 1160 9980
rect 970 9820 1000 9970
rect 1140 9940 1160 9970
rect 1200 9940 1220 9980
rect 1140 9920 1220 9940
rect 1380 9820 1410 10040
rect 1490 9820 1520 10040
rect 1570 9940 1650 9960
rect 1820 9940 1850 10040
rect 1570 9900 1590 9940
rect 1630 9910 1850 9940
rect 1630 9900 1650 9910
rect 1570 9880 1650 9900
rect 1820 9820 1850 9910
rect 1900 9940 1980 9960
rect 2150 9940 2180 10040
rect 2360 9970 2440 9990
rect 1900 9900 1920 9940
rect 1960 9910 2180 9940
rect 1960 9900 1980 9910
rect 1900 9880 1980 9900
rect 2150 9820 2180 9910
rect 2230 9940 2310 9960
rect 2230 9900 2250 9940
rect 2290 9900 2310 9940
rect 2360 9930 2380 9970
rect 2420 9940 2440 9970
rect 2590 9940 2620 10040
rect 2980 9960 3010 10040
rect 3370 10010 3400 10040
rect 3660 10010 3690 10040
rect 2420 9930 2620 9940
rect 2360 9910 2620 9930
rect 2230 9880 2310 9900
rect 2590 9820 2620 9910
rect 2930 9940 3010 9960
rect 2930 9900 2950 9940
rect 2990 9900 3010 9940
rect 3320 9990 4080 10010
rect 3320 9950 3340 9990
rect 3380 9980 4080 9990
rect 3380 9950 3400 9980
rect 3320 9930 3400 9950
rect 2930 9880 3010 9900
rect 2980 9820 3010 9880
rect 3370 9820 3400 9930
rect 3450 9910 3530 9930
rect 3450 9870 3470 9910
rect 3510 9880 3530 9910
rect 3800 9910 3880 9930
rect 3800 9880 3820 9910
rect 3510 9870 3820 9880
rect 3860 9870 3880 9910
rect 3450 9850 3880 9870
rect 3660 9820 3690 9850
rect 4050 9820 4080 9980
rect 5650 9880 5730 9900
rect 5650 9840 5670 9880
rect 5710 9850 5730 9880
rect 8490 9880 8570 9900
rect 8490 9850 8510 9880
rect 5710 9840 5860 9850
rect 5650 9820 5860 9840
rect 590 9490 670 9510
rect 590 9450 610 9490
rect 650 9450 670 9490
rect 590 9430 670 9450
rect 5740 9790 5860 9820
rect 5960 9810 6740 9850
rect 5960 9790 6080 9810
rect 6180 9790 6300 9810
rect 6400 9790 6520 9810
rect 6620 9790 6740 9810
rect 6840 9790 6960 9820
rect 7260 9790 7380 9820
rect 7480 9810 8260 9850
rect 7480 9790 7600 9810
rect 7700 9790 7820 9810
rect 7920 9790 8040 9810
rect 8140 9790 8260 9810
rect 8360 9840 8510 9850
rect 8550 9840 8570 9880
rect 8360 9820 8570 9840
rect 8360 9790 8480 9820
rect -560 9390 -530 9420
rect -450 9390 -420 9420
rect -40 9390 -10 9420
rect 70 9390 100 9420
rect 340 9390 370 9420
rect 450 9390 480 9420
rect 860 9390 890 9420
rect 970 9390 1000 9420
rect 1380 9390 1410 9420
rect 1490 9390 1520 9420
rect 1820 9390 1850 9420
rect 2150 9390 2180 9420
rect 2590 9390 2620 9420
rect 2980 9390 3010 9420
rect 3370 9390 3400 9420
rect 3660 9390 3690 9420
rect 4050 9390 4080 9420
rect 1360 9370 1440 9390
rect 1360 9330 1380 9370
rect 1420 9330 1440 9370
rect 5740 9360 5860 9390
rect 5960 9370 6080 9390
rect 6180 9370 6300 9390
rect 6400 9370 6520 9390
rect 6620 9370 6740 9390
rect 5960 9340 6740 9370
rect 6840 9370 6960 9390
rect 7260 9370 7380 9390
rect 6840 9340 7380 9370
rect 7480 9360 7600 9390
rect 7700 9360 7820 9390
rect 7920 9360 8040 9390
rect 8140 9360 8260 9390
rect 8360 9360 8480 9390
rect 5960 9330 6330 9340
rect 1360 9320 1440 9330
rect 6310 9300 6330 9330
rect 6370 9330 6740 9340
rect 6370 9300 6390 9330
rect 6310 9280 6390 9300
rect 7070 9300 7090 9340
rect 7130 9300 7150 9340
rect 7070 9280 7150 9300
rect 7480 9330 8260 9360
rect 7480 9310 7560 9330
rect 7480 9270 7500 9310
rect 7540 9270 7560 9310
rect 7480 9250 7560 9270
rect 8180 9310 8260 9330
rect 8180 9270 8200 9310
rect 8240 9270 8260 9310
rect 8180 9250 8260 9270
rect -190 9150 -110 9170
rect -190 9110 -170 9150
rect -130 9110 -110 9150
rect -190 9090 -110 9110
rect 2930 9150 3010 9160
rect 2930 9110 2950 9150
rect 2990 9110 3010 9150
rect 2930 9090 3010 9110
rect -560 9060 -530 9090
rect -450 9060 -420 9090
rect -40 9060 -10 9090
rect 70 9060 100 9090
rect 340 9060 370 9090
rect 450 9060 480 9090
rect 860 9060 890 9090
rect 970 9060 1000 9090
rect 1370 9060 1400 9090
rect 1700 9060 1730 9090
rect 2030 9060 2060 9090
rect 2590 9060 2620 9090
rect 2980 9060 3010 9090
rect 3370 9060 3400 9090
rect 3660 9060 3690 9090
rect -310 9030 -230 9050
rect -310 8990 -290 9030
rect -250 8990 -230 9030
rect -310 8970 -230 8990
rect -760 8570 -680 8590
rect -760 8530 -740 8570
rect -700 8540 -680 8570
rect -560 8540 -530 8660
rect -700 8530 -530 8540
rect -760 8510 -530 8530
rect -560 8440 -530 8510
rect -450 8550 -420 8660
rect -450 8530 -350 8550
rect -450 8490 -410 8530
rect -370 8490 -350 8530
rect -450 8470 -350 8490
rect -260 8510 -230 8970
rect 590 9030 670 9050
rect 590 8990 610 9030
rect 650 8990 670 9030
rect 590 8970 670 8990
rect -40 8510 -10 8660
rect -260 8480 -10 8510
rect -450 8440 -420 8470
rect -40 8440 -10 8480
rect 70 8630 100 8660
rect 70 8610 170 8630
rect 70 8570 110 8610
rect 150 8570 170 8610
rect 70 8550 170 8570
rect 70 8440 100 8550
rect 340 8440 370 8660
rect 450 8550 480 8660
rect 450 8530 550 8550
rect 450 8490 490 8530
rect 530 8490 550 8530
rect 450 8470 550 8490
rect 640 8510 670 8970
rect 7920 8810 8000 8830
rect 5890 8770 5970 8790
rect 5890 8740 5910 8770
rect 5760 8730 5910 8740
rect 5950 8740 5970 8770
rect 6430 8780 6510 8800
rect 6430 8740 6450 8780
rect 6490 8740 6510 8780
rect 7510 8780 7590 8800
rect 7510 8740 7530 8780
rect 7570 8740 7590 8780
rect 7920 8770 7940 8810
rect 7980 8770 8000 8810
rect 7920 8750 8000 8770
rect 8180 8810 8260 8830
rect 8180 8770 8200 8810
rect 8240 8770 8260 8810
rect 8180 8750 8260 8770
rect 5950 8730 6100 8740
rect 5540 8690 5660 8720
rect 5760 8710 6100 8730
rect 5760 8690 5880 8710
rect 5980 8690 6100 8710
rect 6200 8710 6740 8740
rect 6200 8690 6320 8710
rect 6620 8690 6740 8710
rect 6840 8710 7180 8740
rect 6840 8690 6960 8710
rect 7060 8690 7180 8710
rect 7280 8710 7820 8740
rect 7280 8690 7400 8710
rect 7700 8690 7820 8710
rect 7920 8720 8260 8750
rect 7920 8690 8040 8720
rect 8140 8690 8260 8720
rect 8360 8690 8480 8720
rect 860 8510 890 8660
rect 640 8480 890 8510
rect 450 8440 480 8470
rect 860 8440 890 8480
rect 970 8600 1000 8660
rect 970 8580 1320 8600
rect 970 8570 1180 8580
rect 970 8440 1000 8570
rect 1160 8540 1180 8570
rect 1220 8540 1260 8580
rect 1300 8540 1320 8580
rect 1160 8520 1320 8540
rect 1370 8570 1400 8660
rect 1570 8580 1650 8600
rect 1570 8570 1590 8580
rect 1370 8540 1590 8570
rect 1630 8540 1650 8580
rect 1370 8440 1400 8540
rect 1570 8520 1650 8540
rect 1700 8570 1730 8660
rect 1900 8580 1980 8600
rect 1900 8570 1920 8580
rect 1700 8540 1920 8570
rect 1960 8540 1980 8580
rect 1700 8440 1730 8540
rect 1900 8520 1980 8540
rect 2030 8570 2060 8660
rect 2190 8580 2270 8600
rect 2190 8570 2210 8580
rect 2030 8540 2210 8570
rect 2250 8540 2270 8580
rect 2030 8440 2060 8540
rect 2190 8520 2270 8540
rect 2340 8570 2420 8590
rect 2340 8530 2360 8570
rect 2400 8540 2420 8570
rect 2590 8540 2620 8660
rect 2980 8630 3010 8660
rect 3370 8620 3400 8660
rect 3660 8620 3690 8660
rect 3060 8600 4080 8620
rect 3060 8560 3080 8600
rect 3120 8590 4080 8600
rect 3120 8560 3140 8590
rect 3060 8540 3140 8560
rect 2400 8530 2620 8540
rect 2340 8510 2620 8530
rect 2590 8440 2620 8510
rect 2980 8440 3010 8470
rect 3370 8440 3400 8590
rect 3450 8520 3530 8530
rect 3450 8480 3470 8520
rect 3510 8490 3530 8520
rect 3510 8480 3690 8490
rect 3450 8460 3690 8480
rect 3660 8440 3690 8460
rect 4050 8440 4080 8590
rect 5540 8260 5660 8290
rect 5450 8240 5660 8260
rect -560 8210 -530 8240
rect -450 8210 -420 8240
rect -40 8160 -10 8240
rect 70 8210 100 8240
rect 340 8160 370 8240
rect 450 8210 480 8240
rect 860 8210 890 8240
rect 970 8210 1000 8240
rect 1370 8210 1400 8240
rect 1700 8210 1730 8240
rect 2030 8210 2060 8240
rect 2590 8210 2620 8240
rect 2980 8210 3010 8240
rect 3370 8210 3400 8240
rect 3660 8210 3690 8240
rect 4050 8210 4080 8240
rect -40 8130 370 8160
rect 2980 8190 3090 8210
rect 2980 8150 3030 8190
rect 3070 8150 3090 8190
rect 2980 8130 3090 8150
rect 3640 8190 3720 8210
rect 3640 8150 3660 8190
rect 3700 8150 3720 8190
rect 5450 8200 5470 8240
rect 5510 8230 5660 8240
rect 5760 8270 5880 8290
rect 5980 8270 6100 8290
rect 5760 8230 6100 8270
rect 6200 8260 6320 8290
rect 6620 8260 6740 8290
rect 6840 8270 6960 8290
rect 7060 8270 7180 8290
rect 5510 8200 5530 8230
rect 5450 8180 5530 8200
rect 5980 8210 6100 8230
rect 6840 8230 7180 8270
rect 7280 8260 7400 8290
rect 7700 8260 7820 8290
rect 7920 8270 8040 8290
rect 8140 8270 8260 8290
rect 7920 8230 8260 8270
rect 8360 8260 8480 8290
rect 8360 8240 8570 8260
rect 8360 8230 8510 8240
rect 6840 8210 6960 8230
rect 5980 8180 6960 8210
rect 8490 8200 8510 8230
rect 8550 8200 8570 8240
rect 8490 8180 8570 8200
rect 3640 8130 3720 8150
rect -1360 6960 -1280 6980
rect -1360 6920 -1340 6960
rect -1300 6930 -1280 6960
rect -40 6960 40 6980
rect -40 6930 -20 6960
rect -1300 6920 -1250 6930
rect -1360 6900 -1250 6920
rect -70 6920 -20 6930
rect 20 6920 40 6960
rect -70 6900 40 6920
rect 540 6960 620 6980
rect 540 6920 560 6960
rect 600 6930 620 6960
rect 1860 6960 1940 6980
rect 1860 6930 1880 6960
rect 600 6920 650 6930
rect 540 6900 650 6920
rect 1830 6920 1880 6930
rect 1920 6920 1940 6960
rect 1830 6900 1940 6920
rect -1280 6870 -1250 6900
rect -1170 6870 -1140 6900
rect -1060 6870 -1030 6900
rect -950 6870 -920 6900
rect -840 6870 -810 6900
rect -730 6870 -700 6900
rect -620 6870 -590 6900
rect -510 6870 -480 6900
rect -400 6870 -370 6900
rect -290 6870 -260 6900
rect -180 6870 -150 6900
rect -70 6870 -40 6900
rect 620 6870 650 6900
rect 730 6870 760 6900
rect 840 6870 870 6900
rect 950 6870 980 6900
rect 1060 6870 1090 6900
rect 1170 6870 1200 6900
rect 1280 6870 1310 6900
rect 1390 6870 1420 6900
rect 1500 6870 1530 6900
rect 1610 6870 1640 6900
rect 1720 6870 1750 6900
rect 1830 6870 1860 6900
rect -1280 6640 -1250 6670
rect -1170 6640 -1140 6670
rect -1060 6640 -1030 6670
rect -950 6640 -920 6670
rect -840 6640 -810 6670
rect -730 6640 -700 6670
rect -620 6640 -590 6670
rect -510 6640 -480 6670
rect -400 6640 -370 6670
rect -290 6640 -260 6670
rect -180 6640 -150 6670
rect -70 6640 -40 6670
rect 620 6640 650 6670
rect 730 6640 760 6670
rect 840 6640 870 6670
rect 950 6640 980 6670
rect 1060 6640 1090 6670
rect 1170 6640 1200 6670
rect 1280 6640 1310 6670
rect 1390 6640 1420 6670
rect 1500 6640 1530 6670
rect 1610 6640 1640 6670
rect 1720 6640 1750 6670
rect 1830 6640 1860 6670
rect -1184 6622 -1126 6640
rect -1184 6588 -1172 6622
rect -1138 6588 -1126 6622
rect -1184 6570 -1126 6588
rect -1074 6622 -1016 6640
rect -1074 6588 -1062 6622
rect -1028 6588 -1016 6622
rect -1074 6570 -1016 6588
rect -964 6622 -906 6640
rect -964 6588 -952 6622
rect -918 6588 -906 6622
rect -964 6570 -906 6588
rect -854 6622 -796 6640
rect -854 6588 -842 6622
rect -808 6588 -796 6622
rect -854 6570 -796 6588
rect -744 6622 -686 6640
rect -744 6588 -732 6622
rect -698 6588 -686 6622
rect -744 6570 -686 6588
rect -634 6622 -576 6640
rect -634 6588 -622 6622
rect -588 6588 -576 6622
rect -634 6570 -576 6588
rect -524 6622 -466 6640
rect -524 6588 -512 6622
rect -478 6588 -466 6622
rect -524 6570 -466 6588
rect -414 6622 -356 6640
rect -414 6588 -402 6622
rect -368 6588 -356 6622
rect -414 6570 -356 6588
rect -304 6622 -246 6640
rect -304 6588 -292 6622
rect -258 6588 -246 6622
rect -304 6570 -246 6588
rect -194 6622 -136 6640
rect -194 6588 -182 6622
rect -148 6588 -136 6622
rect -194 6570 -136 6588
rect 716 6622 774 6640
rect 716 6588 728 6622
rect 762 6588 774 6622
rect 716 6570 774 6588
rect 826 6622 884 6640
rect 826 6588 838 6622
rect 872 6588 884 6622
rect 826 6570 884 6588
rect 936 6622 994 6640
rect 936 6588 948 6622
rect 982 6588 994 6622
rect 936 6570 994 6588
rect 1046 6622 1104 6640
rect 1046 6588 1058 6622
rect 1092 6588 1104 6622
rect 1046 6570 1104 6588
rect 1156 6622 1214 6640
rect 1156 6588 1168 6622
rect 1202 6588 1214 6622
rect 1156 6570 1214 6588
rect 1266 6622 1324 6640
rect 1266 6588 1278 6622
rect 1312 6588 1324 6622
rect 1266 6570 1324 6588
rect 1376 6622 1434 6640
rect 1376 6588 1388 6622
rect 1422 6588 1434 6622
rect 1376 6570 1434 6588
rect 1486 6622 1544 6640
rect 1486 6588 1498 6622
rect 1532 6588 1544 6622
rect 1486 6570 1544 6588
rect 1596 6622 1654 6640
rect 1596 6588 1608 6622
rect 1642 6588 1654 6622
rect 1596 6570 1654 6588
rect 1706 6622 1764 6640
rect 1706 6588 1718 6622
rect 1752 6588 1764 6622
rect 1706 6570 1764 6588
rect -1370 6360 -1290 6380
rect -1370 6320 -1350 6360
rect -1310 6330 -1290 6360
rect 1870 6360 1950 6380
rect 1870 6330 1890 6360
rect -1310 6320 -1190 6330
rect -1370 6300 -1190 6320
rect 1770 6320 1890 6330
rect 1930 6320 1950 6360
rect 1770 6300 1950 6320
rect 5354 6340 5784 6356
rect 5354 6306 5370 6340
rect 5404 6306 5784 6340
rect -1290 6270 -1190 6300
rect -1110 6270 -1010 6300
rect -930 6270 -830 6300
rect -750 6270 -650 6300
rect -570 6270 -470 6300
rect -390 6270 -290 6300
rect -210 6270 -110 6300
rect -30 6270 70 6300
rect 150 6270 250 6300
rect 330 6270 430 6300
rect 510 6270 610 6300
rect 690 6270 790 6300
rect 870 6270 970 6300
rect 1050 6270 1150 6300
rect 1230 6270 1330 6300
rect 1410 6270 1510 6300
rect 1590 6270 1690 6300
rect 1770 6270 1870 6300
rect 5354 6290 5784 6306
rect 6264 6340 6694 6356
rect 6264 6306 6644 6340
rect 6678 6306 6694 6340
rect 6264 6290 6694 6306
rect 2510 6160 2570 6180
rect 2510 6120 2520 6160
rect 2560 6120 2570 6160
rect 2950 6160 3010 6180
rect 2950 6120 2960 6160
rect 3000 6120 3010 6160
rect 2510 6090 2610 6120
rect 2580 6070 2610 6090
rect 2690 6070 2720 6100
rect 2800 6070 2830 6100
rect 2910 6090 3010 6120
rect 6310 6150 6390 6170
rect 6310 6110 6330 6150
rect 6370 6110 6390 6150
rect 6710 6150 6790 6170
rect 6710 6110 6730 6150
rect 6770 6110 6790 6150
rect 2910 6070 2940 6090
rect 5600 6060 5700 6090
rect 5800 6080 7300 6110
rect 5800 6060 5900 6080
rect 6000 6060 6100 6080
rect 6200 6060 6300 6080
rect 6400 6060 6500 6080
rect 6600 6060 6700 6080
rect 6800 6060 6900 6080
rect 7000 6060 7100 6080
rect 7200 6060 7300 6080
rect 7400 6060 7500 6090
rect 2580 5840 2610 5870
rect 2690 5850 2720 5870
rect 2800 5850 2830 5870
rect 2690 5820 2830 5850
rect 2910 5840 2940 5870
rect 2720 5780 2740 5820
rect 2780 5780 2800 5820
rect 5600 5780 5700 5810
rect 5800 5780 5900 5810
rect 6000 5780 6100 5810
rect 6200 5780 6300 5810
rect 6400 5780 6500 5810
rect 6600 5780 6700 5810
rect 6800 5780 6900 5810
rect 7000 5780 7100 5810
rect 7200 5780 7300 5810
rect 7400 5780 7500 5810
rect 2720 5760 2800 5780
rect 5510 5760 5700 5780
rect 5510 5720 5530 5760
rect 5570 5750 5700 5760
rect 7400 5760 7590 5780
rect 7400 5750 7530 5760
rect 5570 5720 5590 5750
rect 5510 5700 5590 5720
rect 7510 5720 7530 5750
rect 7570 5720 7590 5760
rect 7510 5700 7590 5720
rect -1290 5640 -1190 5670
rect -1110 5640 -1010 5670
rect -930 5640 -830 5670
rect -750 5640 -650 5670
rect -570 5640 -470 5670
rect -390 5640 -290 5670
rect -210 5640 -110 5670
rect -30 5640 70 5670
rect 150 5640 250 5670
rect 330 5640 430 5670
rect 510 5640 610 5670
rect 690 5640 790 5670
rect 870 5640 970 5670
rect 1050 5640 1150 5670
rect 1230 5640 1330 5670
rect 1410 5640 1510 5670
rect -1090 5620 -1020 5640
rect -1090 5580 -1080 5620
rect -1040 5580 -1020 5620
rect -1090 5560 -1020 5580
rect -920 5620 -840 5640
rect -920 5580 -900 5620
rect -860 5580 -840 5620
rect -920 5560 -840 5580
rect -740 5620 -660 5640
rect -740 5580 -720 5620
rect -680 5580 -660 5620
rect -740 5560 -660 5580
rect -560 5620 -480 5640
rect -560 5580 -540 5620
rect -500 5580 -480 5620
rect -560 5560 -480 5580
rect -380 5620 -300 5640
rect -380 5580 -360 5620
rect -320 5580 -300 5620
rect -380 5560 -300 5580
rect -200 5620 -120 5640
rect -200 5580 -180 5620
rect -140 5580 -120 5620
rect -200 5560 -120 5580
rect -20 5620 60 5640
rect -20 5580 0 5620
rect 40 5580 60 5620
rect -20 5560 60 5580
rect 160 5620 230 5640
rect 160 5580 180 5620
rect 220 5580 230 5620
rect 160 5560 230 5580
rect 350 5620 420 5640
rect 350 5580 360 5620
rect 400 5580 420 5620
rect 350 5560 420 5580
rect 520 5620 600 5640
rect 520 5580 540 5620
rect 580 5580 600 5620
rect 520 5560 600 5580
rect 700 5620 780 5640
rect 700 5580 720 5620
rect 760 5580 780 5620
rect 700 5560 780 5580
rect 880 5620 960 5640
rect 880 5580 900 5620
rect 940 5580 960 5620
rect 880 5560 960 5580
rect 1060 5620 1140 5640
rect 1060 5580 1080 5620
rect 1120 5580 1140 5620
rect 1060 5560 1140 5580
rect 1240 5620 1320 5640
rect 1240 5580 1260 5620
rect 1300 5580 1320 5620
rect 1240 5560 1320 5580
rect 1420 5620 1500 5640
rect 1590 5630 1690 5670
rect 1770 5640 1870 5670
rect 1420 5580 1440 5620
rect 1480 5580 1500 5620
rect 1420 5560 1500 5580
rect 1600 5620 1670 5630
rect 1600 5580 1620 5620
rect 1660 5580 1670 5620
rect 1600 5560 1670 5580
rect 5620 5470 5710 5490
rect 5620 5420 5640 5470
rect 5690 5420 5710 5470
rect 5620 5400 5710 5420
rect 6270 5470 6360 5490
rect 6270 5420 6290 5470
rect 6340 5420 6360 5470
rect 6270 5400 6360 5420
rect 6760 5460 6840 5480
rect 6760 5420 6780 5460
rect 6820 5420 6840 5460
rect 6760 5400 6840 5420
rect 7420 5460 7500 5480
rect 7420 5420 7440 5460
rect 7480 5420 7500 5460
rect 7420 5400 7500 5420
rect 7900 5460 7980 5480
rect 7900 5420 7920 5460
rect 7960 5420 7980 5460
rect 7900 5400 7980 5420
rect 8560 5460 8640 5480
rect 8560 5420 8580 5460
rect 8620 5420 8640 5460
rect 8560 5400 8640 5420
rect 5650 5370 5680 5400
rect 5780 5370 5810 5400
rect 5910 5370 5940 5400
rect 6040 5370 6070 5400
rect 6170 5370 6200 5400
rect 6300 5370 6330 5400
rect 6790 5370 6820 5400
rect 6920 5370 6950 5400
rect 7050 5370 7080 5400
rect 7180 5370 7210 5400
rect 7310 5370 7340 5400
rect 7440 5370 7470 5400
rect 7930 5370 7960 5400
rect 8060 5370 8090 5400
rect 8190 5370 8220 5400
rect 8320 5370 8350 5400
rect 8450 5370 8480 5400
rect 8580 5370 8610 5400
rect 5650 5240 5680 5270
rect 5780 5250 5810 5270
rect 5910 5250 5940 5270
rect 6040 5250 6070 5270
rect 6170 5250 6200 5270
rect 5780 5220 6200 5250
rect 6300 5240 6330 5270
rect 6790 5240 6820 5270
rect 6920 5250 6950 5270
rect 7050 5250 7080 5270
rect 6920 5240 7080 5250
rect 6870 5220 7080 5240
rect 7180 5250 7210 5270
rect 7310 5250 7340 5270
rect 7180 5240 7340 5250
rect 7440 5240 7470 5270
rect 7930 5240 7960 5270
rect 7180 5220 7390 5240
rect 5820 5180 5840 5220
rect 5880 5180 5900 5220
rect 5820 5160 5900 5180
rect 6870 5180 6890 5220
rect 6930 5180 6950 5220
rect 6870 5160 6950 5180
rect 7310 5180 7330 5220
rect 7370 5180 7390 5220
rect 7310 5160 7390 5180
rect 8060 5190 8090 5270
rect 8190 5190 8220 5270
rect 8320 5190 8350 5270
rect 8450 5190 8480 5270
rect 8580 5240 8610 5270
rect 8850 5220 8930 5240
rect 8850 5190 8870 5220
rect 8060 5180 8870 5190
rect 8910 5180 8930 5220
rect 8060 5160 8930 5180
rect 8060 5120 8090 5160
rect 8010 5100 8090 5120
rect 8010 5060 8030 5100
rect 8070 5060 8090 5100
rect 8010 5040 8090 5060
rect 5730 4880 5810 4900
rect 5730 4840 5750 4880
rect 5790 4840 5810 4880
rect 6170 4880 6250 4900
rect 6170 4840 6190 4880
rect 6230 4840 6250 4880
rect 6960 4890 7040 4910
rect 6960 4850 6980 4890
rect 7020 4850 7040 4890
rect 6960 4840 7040 4850
rect 8010 4880 8930 4900
rect 8010 4840 8030 4880
rect 8070 4870 8870 4880
rect 8070 4840 8090 4870
rect 5730 4820 5940 4840
rect -2460 4800 -2400 4820
rect -2460 4760 -2450 4800
rect -2410 4770 -2400 4800
rect -60 4800 0 4820
rect -60 4770 -50 4800
rect -2410 4760 -2350 4770
rect -2460 4740 -2350 4760
rect -110 4760 -50 4770
rect -10 4760 0 4800
rect -110 4740 0 4760
rect 580 4800 640 4820
rect 580 4760 590 4800
rect 630 4770 640 4800
rect 2980 4800 3040 4820
rect 2980 4770 2990 4800
rect 630 4760 690 4770
rect 580 4740 690 4760
rect 2930 4760 2990 4770
rect 3030 4760 3040 4800
rect 5650 4790 5680 4820
rect 5780 4810 5940 4820
rect 5780 4790 5810 4810
rect 5910 4790 5940 4810
rect 6040 4820 6250 4840
rect 6040 4810 6200 4820
rect 6040 4790 6070 4810
rect 6170 4790 6200 4810
rect 6300 4790 6330 4820
rect 6790 4790 6820 4820
rect 6920 4810 7340 4840
rect 8010 4820 8090 4840
rect 6920 4790 6950 4810
rect 7050 4790 7080 4810
rect 7180 4790 7210 4810
rect 7310 4790 7340 4810
rect 7440 4790 7470 4820
rect 7930 4790 7960 4820
rect 8060 4790 8090 4820
rect 8190 4790 8220 4870
rect 8320 4790 8350 4870
rect 8450 4790 8480 4870
rect 8850 4840 8870 4870
rect 8910 4840 8930 4880
rect 8850 4820 8930 4840
rect 8580 4790 8610 4820
rect 2930 4740 3040 4760
rect -2390 4710 -2350 4740
rect -2270 4710 -2230 4740
rect -2150 4710 -2110 4740
rect -2030 4710 -1990 4740
rect -1910 4710 -1870 4740
rect -1790 4710 -1750 4740
rect -1670 4710 -1630 4740
rect -1550 4710 -1510 4740
rect -1430 4710 -1390 4740
rect -1310 4710 -1270 4740
rect -1190 4710 -1150 4740
rect -1070 4710 -1030 4740
rect -950 4710 -910 4740
rect -830 4710 -790 4740
rect -710 4710 -670 4740
rect -590 4710 -550 4740
rect -470 4710 -430 4740
rect -350 4710 -310 4740
rect -230 4710 -190 4740
rect -110 4710 -70 4740
rect 650 4710 690 4740
rect 770 4710 810 4740
rect 890 4710 930 4740
rect 1010 4710 1050 4740
rect 1130 4710 1170 4740
rect 1250 4710 1290 4740
rect 1370 4710 1410 4740
rect 1490 4710 1530 4740
rect 1610 4710 1650 4740
rect 1730 4710 1770 4740
rect 1850 4710 1890 4740
rect 1970 4710 2010 4740
rect 2090 4710 2130 4740
rect 2210 4710 2250 4740
rect 2330 4710 2370 4740
rect 2450 4710 2490 4740
rect 2570 4710 2610 4740
rect 2690 4710 2730 4740
rect 2810 4710 2850 4740
rect 2930 4710 2970 4740
rect 5650 4560 5680 4590
rect 5780 4560 5810 4590
rect 5910 4560 5940 4590
rect 6040 4560 6070 4590
rect 6170 4560 6200 4590
rect 6300 4560 6330 4590
rect 6790 4560 6820 4590
rect 6920 4560 6950 4590
rect 7050 4560 7080 4590
rect 7180 4560 7210 4590
rect 7310 4560 7340 4590
rect 7440 4560 7470 4590
rect 7930 4560 7960 4590
rect 8060 4560 8090 4590
rect 8190 4560 8220 4590
rect 8320 4560 8350 4590
rect 8450 4560 8480 4590
rect 8580 4560 8610 4590
rect 5620 4540 5700 4560
rect -2390 4480 -2350 4510
rect -2270 4470 -2230 4510
rect -2150 4490 -2110 4510
rect -2030 4490 -1990 4510
rect -1910 4490 -1870 4510
rect -1790 4490 -1750 4510
rect -2280 4450 -2220 4470
rect -2150 4460 -1750 4490
rect -1670 4490 -1630 4510
rect -1550 4490 -1510 4510
rect -1670 4460 -1510 4490
rect -1430 4490 -1390 4510
rect -1310 4490 -1270 4510
rect -1190 4490 -1150 4510
rect -1070 4490 -1030 4510
rect -1430 4460 -1030 4490
rect -950 4490 -910 4510
rect -830 4490 -790 4510
rect -950 4460 -790 4490
rect -710 4490 -670 4510
rect -590 4490 -550 4510
rect -470 4490 -430 4510
rect -350 4490 -310 4510
rect -710 4460 -310 4490
rect -230 4480 -190 4510
rect -110 4480 -70 4510
rect 650 4480 690 4510
rect 770 4480 810 4510
rect 890 4490 930 4510
rect 1010 4490 1050 4510
rect 1130 4490 1170 4510
rect 1250 4490 1290 4510
rect -240 4460 -180 4480
rect -2280 4410 -2270 4450
rect -2230 4410 -2220 4450
rect -2280 4390 -2220 4410
rect -2110 4420 -2090 4460
rect -2050 4420 -2030 4460
rect -2110 4400 -2030 4420
rect -1620 4420 -1610 4460
rect -1570 4420 -1560 4460
rect -1620 4400 -1560 4420
rect -1390 4420 -1370 4460
rect -1330 4420 -1310 4460
rect -1390 4400 -1310 4420
rect -900 4420 -890 4460
rect -850 4420 -840 4460
rect -900 4400 -840 4420
rect -670 4420 -650 4460
rect -610 4420 -590 4460
rect -670 4400 -590 4420
rect -240 4420 -230 4460
rect -190 4420 -180 4460
rect -240 4400 -180 4420
rect 760 4460 820 4480
rect 890 4460 1290 4490
rect 1370 4490 1410 4510
rect 1490 4490 1530 4510
rect 1370 4460 1530 4490
rect 1610 4490 1650 4510
rect 1730 4490 1770 4510
rect 1850 4490 1890 4510
rect 1970 4490 2010 4510
rect 1610 4460 2010 4490
rect 2090 4490 2130 4510
rect 2210 4490 2250 4510
rect 2090 4460 2250 4490
rect 2330 4490 2370 4510
rect 2450 4490 2490 4510
rect 2570 4490 2610 4510
rect 2690 4490 2730 4510
rect 2330 4460 2730 4490
rect 2810 4470 2850 4510
rect 2930 4480 2970 4510
rect 5620 4500 5640 4540
rect 5680 4500 5700 4540
rect 5620 4480 5700 4500
rect 6280 4540 6360 4560
rect 6280 4500 6300 4540
rect 6340 4500 6360 4540
rect 6280 4480 6360 4500
rect 6760 4540 6840 4560
rect 6760 4500 6780 4540
rect 6820 4500 6840 4540
rect 6760 4480 6840 4500
rect 7420 4540 7500 4560
rect 7420 4500 7440 4540
rect 7480 4500 7500 4540
rect 7420 4480 7500 4500
rect 7900 4540 7980 4560
rect 7900 4500 7920 4540
rect 7960 4500 7980 4540
rect 7900 4480 7980 4500
rect 8560 4540 8640 4560
rect 8560 4500 8580 4540
rect 8620 4500 8640 4540
rect 8560 4480 8640 4500
rect 760 4420 770 4460
rect 810 4420 820 4460
rect 760 4400 820 4420
rect 1170 4420 1190 4460
rect 1230 4420 1250 4460
rect 1170 4400 1250 4420
rect 1420 4420 1430 4460
rect 1470 4420 1480 4460
rect 1420 4400 1480 4420
rect 1890 4420 1910 4460
rect 1950 4420 1970 4460
rect 1890 4400 1970 4420
rect 2140 4420 2150 4460
rect 2190 4420 2200 4460
rect 2140 4400 2200 4420
rect 2610 4420 2630 4460
rect 2670 4420 2690 4460
rect 2610 4400 2690 4420
rect 2800 4450 2860 4470
rect 2800 4410 2810 4450
rect 2850 4410 2860 4450
rect 2800 4390 2860 4410
rect 5630 4230 5710 4250
rect 5630 4190 5650 4230
rect 5690 4200 5710 4230
rect 7630 4230 7710 4250
rect 7630 4200 7650 4230
rect 5690 4190 5820 4200
rect 5630 4170 5820 4190
rect 7520 4190 7650 4200
rect 7690 4190 7710 4230
rect 7520 4170 7710 4190
rect 5720 4140 5820 4170
rect 5920 4140 6020 4170
rect 6120 4140 6220 4170
rect 6320 4140 6420 4170
rect 6520 4140 6620 4170
rect 6720 4140 6820 4170
rect 6920 4140 7020 4170
rect 7120 4140 7220 4170
rect 7320 4140 7420 4170
rect 7520 4140 7620 4170
rect -1458 3852 -1390 3870
rect -1458 3818 -1446 3852
rect -1412 3818 -1390 3852
rect -1458 3800 -1390 3818
rect -1550 3770 -1510 3800
rect -1430 3770 -1390 3800
rect -1310 3852 -1242 3870
rect -1310 3818 -1288 3852
rect -1254 3818 -1242 3852
rect -1310 3800 -1242 3818
rect -976 3852 -910 3870
rect -976 3818 -964 3852
rect -930 3818 -910 3852
rect -976 3800 -910 3818
rect -1310 3770 -1270 3800
rect -1190 3770 -1150 3800
rect -1070 3770 -1030 3800
rect -950 3770 -910 3800
rect -830 3852 -764 3870
rect -830 3818 -810 3852
rect -776 3818 -764 3852
rect -830 3800 -764 3818
rect -498 3852 -430 3870
rect -498 3818 -486 3852
rect -452 3818 -430 3852
rect 1010 3852 1078 3870
rect -498 3800 -430 3818
rect -830 3770 -790 3800
rect -710 3770 -670 3800
rect -590 3770 -550 3800
rect -470 3770 -430 3800
rect -1550 3640 -1510 3670
rect -1430 3640 -1390 3670
rect -1310 3640 -1270 3670
rect -1190 3640 -1150 3670
rect -1070 3640 -1030 3670
rect -950 3640 -910 3670
rect -830 3640 -790 3670
rect -710 3640 -670 3670
rect -590 3640 -550 3670
rect -470 3640 -430 3670
rect -1559 3622 -1501 3640
rect -1559 3588 -1547 3622
rect -1513 3588 -1501 3622
rect -1559 3570 -1501 3588
rect -1199 3622 -1141 3640
rect -1199 3588 -1187 3622
rect -1153 3588 -1141 3622
rect -1199 3570 -1141 3588
rect -1079 3622 -1021 3640
rect -1079 3588 -1067 3622
rect -1033 3588 -1021 3622
rect -1079 3570 -1021 3588
rect -719 3622 -661 3640
rect -719 3588 -707 3622
rect -673 3588 -661 3622
rect -719 3570 -661 3588
rect -599 3622 -541 3640
rect -599 3588 -587 3622
rect -553 3588 -541 3622
rect -599 3570 -541 3588
rect 1010 3818 1032 3852
rect 1066 3818 1078 3852
rect 1010 3800 1078 3818
rect 1344 3852 1410 3870
rect 1344 3818 1356 3852
rect 1390 3818 1410 3852
rect 1344 3800 1410 3818
rect 1010 3770 1050 3800
rect 1130 3770 1170 3800
rect 1250 3770 1290 3800
rect 1370 3770 1410 3800
rect 1490 3852 1556 3870
rect 1490 3818 1510 3852
rect 1544 3818 1556 3852
rect 1490 3800 1556 3818
rect 1822 3852 1890 3870
rect 1822 3818 1834 3852
rect 1868 3818 1890 3852
rect 1822 3800 1890 3818
rect 1490 3770 1530 3800
rect 1610 3770 1650 3800
rect 1730 3770 1770 3800
rect 1850 3770 1890 3800
rect 1970 3852 2038 3870
rect 1970 3818 1992 3852
rect 2026 3818 2038 3852
rect 1970 3800 2038 3818
rect 1970 3770 2010 3800
rect 2090 3770 2130 3800
rect 1010 3640 1050 3670
rect 1130 3640 1170 3670
rect 1250 3640 1290 3670
rect 1370 3640 1410 3670
rect 1490 3640 1530 3670
rect 1610 3640 1650 3670
rect 1730 3640 1770 3670
rect 1850 3640 1890 3670
rect 1970 3640 2010 3670
rect 2090 3640 2130 3670
rect 1121 3622 1179 3640
rect 1121 3588 1133 3622
rect 1167 3588 1179 3622
rect 1121 3570 1179 3588
rect 1241 3622 1299 3640
rect 1241 3588 1253 3622
rect 1287 3588 1299 3622
rect 1241 3570 1299 3588
rect 1601 3622 1659 3640
rect 1601 3588 1613 3622
rect 1647 3588 1659 3622
rect 1601 3570 1659 3588
rect 1721 3622 1779 3640
rect 1721 3588 1733 3622
rect 1767 3588 1779 3622
rect 1721 3570 1779 3588
rect 2081 3622 2139 3640
rect 2081 3588 2093 3622
rect 2127 3588 2139 3622
rect 5720 3610 5820 3640
rect 5920 3620 6020 3640
rect 6120 3620 6220 3640
rect 6320 3620 6420 3640
rect 6520 3620 6620 3640
rect 6720 3620 6820 3640
rect 6920 3620 7020 3640
rect 7120 3620 7220 3640
rect 7320 3620 7420 3640
rect 5920 3590 7420 3620
rect 7520 3610 7620 3640
rect 2081 3570 2139 3588
rect 6430 3550 6450 3590
rect 6490 3550 6510 3590
rect 6430 3530 6510 3550
rect 6830 3550 6850 3590
rect 6890 3550 6910 3590
rect 6830 3530 6910 3550
rect -2070 3250 -1990 3270
rect -2070 3210 -2050 3250
rect -2010 3210 -1990 3250
rect -2070 3190 -1990 3210
rect -1830 3250 -1750 3270
rect -1830 3210 -1810 3250
rect -1770 3210 -1750 3250
rect -1830 3190 -1750 3210
rect -1590 3250 -1510 3270
rect -1590 3210 -1570 3250
rect -1530 3210 -1510 3250
rect -1590 3190 -1510 3210
rect -1350 3250 -1270 3270
rect -1350 3210 -1330 3250
rect -1290 3210 -1270 3250
rect -1350 3190 -1270 3210
rect -710 3250 -630 3270
rect -710 3210 -690 3250
rect -650 3210 -630 3250
rect -710 3190 -630 3210
rect -470 3250 -390 3270
rect -470 3210 -450 3250
rect -410 3210 -390 3250
rect -470 3190 -390 3210
rect -230 3250 -150 3270
rect -230 3210 -210 3250
rect -170 3210 -150 3250
rect -230 3190 -150 3210
rect 730 3250 810 3270
rect 730 3210 750 3250
rect 790 3210 810 3250
rect 730 3190 810 3210
rect 970 3250 1050 3270
rect 970 3210 990 3250
rect 1030 3210 1050 3250
rect 970 3190 1050 3210
rect 1210 3250 1290 3270
rect 1210 3210 1230 3250
rect 1270 3210 1290 3250
rect 1210 3190 1290 3210
rect 1850 3250 1930 3270
rect 1850 3210 1870 3250
rect 1910 3210 1930 3250
rect 1850 3190 1930 3210
rect 2090 3250 2170 3270
rect 2090 3210 2110 3250
rect 2150 3210 2170 3250
rect 2090 3190 2170 3210
rect 2330 3250 2410 3270
rect 2330 3210 2350 3250
rect 2390 3210 2410 3250
rect 2330 3190 2410 3210
rect 2570 3250 2650 3270
rect 2570 3210 2590 3250
rect 2630 3210 2650 3250
rect 2570 3190 2650 3210
rect -2170 3160 -1170 3190
rect -930 3160 70 3190
rect 510 3160 1510 3190
rect 1750 3160 2750 3190
rect -2170 2630 -1170 2660
rect -930 2630 70 2660
rect 510 2630 1510 2660
rect 1750 2630 2750 2660
rect -1670 2340 -1590 2360
rect -1670 2300 -1650 2340
rect -1610 2300 -1590 2340
rect -1670 2280 -1590 2300
rect -1510 2340 -1430 2360
rect -1510 2300 -1490 2340
rect -1450 2300 -1430 2340
rect -1510 2280 -1430 2300
rect -1350 2340 -1270 2360
rect -1350 2300 -1330 2340
rect -1290 2300 -1270 2340
rect -1350 2280 -1270 2300
rect -1190 2340 -1110 2360
rect -1190 2300 -1170 2340
rect -1130 2300 -1110 2340
rect -1190 2280 -1110 2300
rect -1030 2340 -950 2360
rect -1030 2300 -1010 2340
rect -970 2300 -950 2340
rect -1030 2280 -950 2300
rect -870 2340 -790 2360
rect -870 2300 -850 2340
rect -810 2300 -790 2340
rect -870 2280 -790 2300
rect -710 2340 -630 2360
rect -710 2300 -690 2340
rect -650 2300 -630 2340
rect -710 2280 -630 2300
rect -550 2340 -470 2360
rect -550 2300 -530 2340
rect -490 2300 -470 2340
rect -550 2280 -470 2300
rect -390 2340 -310 2360
rect -390 2300 -370 2340
rect -330 2300 -310 2340
rect -390 2280 -310 2300
rect -230 2340 -150 2360
rect -230 2300 -210 2340
rect -170 2300 -150 2340
rect -230 2280 -150 2300
rect -70 2340 10 2360
rect -70 2300 -50 2340
rect -10 2300 10 2340
rect -70 2280 10 2300
rect 90 2340 170 2360
rect 90 2300 110 2340
rect 150 2300 170 2340
rect 90 2280 170 2300
rect 410 2340 490 2360
rect 410 2300 430 2340
rect 470 2300 490 2340
rect 410 2280 490 2300
rect 570 2340 650 2360
rect 570 2300 590 2340
rect 630 2300 650 2340
rect 570 2280 650 2300
rect 730 2340 810 2360
rect 730 2300 750 2340
rect 790 2300 810 2340
rect 730 2280 810 2300
rect 890 2340 970 2360
rect 890 2300 910 2340
rect 950 2300 970 2340
rect 890 2280 970 2300
rect 1050 2340 1130 2360
rect 1050 2300 1070 2340
rect 1110 2300 1130 2340
rect 1050 2280 1130 2300
rect 1210 2340 1290 2360
rect 1210 2300 1230 2340
rect 1270 2300 1290 2340
rect 1210 2280 1290 2300
rect 1370 2340 1450 2360
rect 1370 2300 1390 2340
rect 1430 2300 1450 2340
rect 1370 2280 1450 2300
rect 1530 2340 1610 2360
rect 1530 2300 1550 2340
rect 1590 2300 1610 2340
rect 1530 2280 1610 2300
rect 1690 2340 1770 2360
rect 1690 2300 1710 2340
rect 1750 2300 1770 2340
rect 1690 2280 1770 2300
rect 1850 2340 1930 2360
rect 1850 2300 1870 2340
rect 1910 2300 1930 2340
rect 1850 2280 1930 2300
rect 2010 2340 2090 2360
rect 2010 2300 2030 2340
rect 2070 2300 2090 2340
rect 2010 2280 2090 2300
rect 2170 2340 2250 2360
rect 2170 2300 2190 2340
rect 2230 2300 2250 2340
rect 2170 2280 2250 2300
rect -1750 2250 250 2280
rect 330 2250 2330 2280
rect -1750 2020 250 2050
rect 330 2020 2330 2050
<< polycont >>
rect 9378 13508 9412 13542
rect 9898 13508 9932 13542
rect 10418 13508 10452 13542
rect 10986 13508 11020 13542
rect -1490 12890 -1450 12930
rect -540 12870 -500 12910
rect 530 12880 570 12920
rect 2090 12880 2130 12920
rect 4694 12890 4734 12930
rect -1380 12650 -1340 12690
rect -800 12650 -760 12690
rect 5250 12740 5290 12780
rect -460 12650 -420 12690
rect -1510 12450 -1470 12490
rect -260 12570 -220 12610
rect 120 12650 160 12690
rect 140 12530 180 12570
rect 640 12650 680 12690
rect 990 12650 1030 12690
rect 1570 12650 1610 12690
rect 1780 12650 1820 12690
rect 2020 12650 2060 12690
rect 2360 12640 2400 12680
rect 2630 12600 2670 12640
rect 1840 12530 1880 12570
rect 2830 12570 2870 12610
rect 3260 12650 3300 12690
rect 3230 12530 3270 12570
rect 3620 12650 3660 12690
rect 3950 12650 3990 12690
rect 4530 12650 4570 12690
rect 4360 12570 4400 12610
rect 5000 12630 5040 12670
rect 5830 12740 5870 12780
rect 6550 12740 6590 12780
rect 6300 12630 6340 12670
rect 5660 12570 5700 12610
rect 7130 12740 7170 12780
rect 7850 12740 7890 12780
rect 7600 12630 7640 12670
rect 6960 12570 7000 12610
rect 8430 12740 8470 12780
rect 9392 13128 9426 13162
rect 9912 13128 9946 13162
rect 10432 13128 10466 13162
rect 9364 12848 9398 12882
rect 9884 12848 9918 12882
rect 10404 12848 10438 12882
rect 8260 12570 8300 12610
rect 8874 12628 8908 12662
rect 3820 12450 3860 12490
rect -850 12330 -810 12370
rect -540 12350 -500 12390
rect 270 12330 310 12370
rect 400 12330 440 12370
rect 1530 12330 1570 12370
rect 3290 12320 3330 12360
rect 5820 12330 5860 12370
rect 7120 12330 7160 12370
rect 8420 12330 8460 12370
rect 9364 12418 9398 12452
rect 9884 12418 9918 12452
rect 10404 12418 10438 12452
rect 9392 12038 9426 12072
rect 9912 12038 9946 12072
rect 10432 12038 10466 12072
rect 9510 11350 9550 11390
rect 10030 11350 10070 11390
rect 10550 11350 10590 11390
rect 11070 11350 11110 11390
rect 1510 10290 1550 10330
rect -740 9910 -700 9950
rect -410 9950 -370 9990
rect 110 9870 150 9910
rect 490 9950 530 9990
rect -290 9450 -250 9490
rect 1160 9940 1200 9980
rect 1590 9900 1630 9940
rect 1920 9900 1960 9940
rect 2250 9900 2290 9940
rect 2380 9930 2420 9970
rect 2950 9900 2990 9940
rect 3340 9950 3380 9990
rect 3470 9870 3510 9910
rect 3820 9870 3860 9910
rect 5670 9840 5710 9880
rect 610 9450 650 9490
rect 8510 9840 8550 9880
rect 1380 9330 1420 9370
rect 6330 9300 6370 9340
rect 7090 9300 7130 9340
rect 7500 9270 7540 9310
rect 8200 9270 8240 9310
rect -170 9110 -130 9150
rect 2950 9110 2990 9150
rect -290 8990 -250 9030
rect -740 8530 -700 8570
rect -410 8490 -370 8530
rect 610 8990 650 9030
rect 110 8570 150 8610
rect 490 8490 530 8530
rect 5910 8730 5950 8770
rect 6450 8740 6490 8780
rect 7530 8740 7570 8780
rect 7940 8770 7980 8810
rect 8200 8770 8240 8810
rect 1180 8540 1220 8580
rect 1260 8540 1300 8580
rect 1590 8540 1630 8580
rect 1920 8540 1960 8580
rect 2210 8540 2250 8580
rect 2360 8530 2400 8570
rect 3080 8560 3120 8600
rect 3470 8480 3510 8520
rect 3030 8150 3070 8190
rect 3660 8150 3700 8190
rect 5470 8200 5510 8240
rect 8510 8200 8550 8240
rect -1340 6920 -1300 6960
rect -20 6920 20 6960
rect 560 6920 600 6960
rect 1880 6920 1920 6960
rect -1172 6588 -1138 6622
rect -1062 6588 -1028 6622
rect -952 6588 -918 6622
rect -842 6588 -808 6622
rect -732 6588 -698 6622
rect -622 6588 -588 6622
rect -512 6588 -478 6622
rect -402 6588 -368 6622
rect -292 6588 -258 6622
rect -182 6588 -148 6622
rect 728 6588 762 6622
rect 838 6588 872 6622
rect 948 6588 982 6622
rect 1058 6588 1092 6622
rect 1168 6588 1202 6622
rect 1278 6588 1312 6622
rect 1388 6588 1422 6622
rect 1498 6588 1532 6622
rect 1608 6588 1642 6622
rect 1718 6588 1752 6622
rect -1350 6320 -1310 6360
rect 1890 6320 1930 6360
rect 5370 6306 5404 6340
rect 6644 6306 6678 6340
rect 2520 6120 2560 6160
rect 2960 6120 3000 6160
rect 6330 6110 6370 6150
rect 6730 6110 6770 6150
rect 2740 5780 2780 5820
rect 5530 5720 5570 5760
rect 7530 5720 7570 5760
rect -1080 5580 -1040 5620
rect -900 5580 -860 5620
rect -720 5580 -680 5620
rect -540 5580 -500 5620
rect -360 5580 -320 5620
rect -180 5580 -140 5620
rect 0 5580 40 5620
rect 180 5580 220 5620
rect 360 5580 400 5620
rect 540 5580 580 5620
rect 720 5580 760 5620
rect 900 5580 940 5620
rect 1080 5580 1120 5620
rect 1260 5580 1300 5620
rect 1440 5580 1480 5620
rect 1620 5580 1660 5620
rect 5640 5420 5690 5470
rect 6290 5420 6340 5470
rect 6780 5420 6820 5460
rect 7440 5420 7480 5460
rect 7920 5420 7960 5460
rect 8580 5420 8620 5460
rect 5840 5180 5880 5220
rect 6890 5180 6930 5220
rect 7330 5180 7370 5220
rect 8870 5180 8910 5220
rect 8030 5060 8070 5100
rect 5750 4840 5790 4880
rect 6190 4840 6230 4880
rect 6980 4850 7020 4890
rect 8030 4840 8070 4880
rect -2450 4760 -2410 4800
rect -50 4760 -10 4800
rect 590 4760 630 4800
rect 2990 4760 3030 4800
rect 8870 4840 8910 4880
rect -2270 4410 -2230 4450
rect -2090 4420 -2050 4460
rect -1610 4420 -1570 4460
rect -1370 4420 -1330 4460
rect -890 4420 -850 4460
rect -650 4420 -610 4460
rect -230 4420 -190 4460
rect 5640 4500 5680 4540
rect 6300 4500 6340 4540
rect 6780 4500 6820 4540
rect 7440 4500 7480 4540
rect 7920 4500 7960 4540
rect 8580 4500 8620 4540
rect 770 4420 810 4460
rect 1190 4420 1230 4460
rect 1430 4420 1470 4460
rect 1910 4420 1950 4460
rect 2150 4420 2190 4460
rect 2630 4420 2670 4460
rect 2810 4410 2850 4450
rect 5650 4190 5690 4230
rect 7650 4190 7690 4230
rect -1446 3818 -1412 3852
rect -1288 3818 -1254 3852
rect -964 3818 -930 3852
rect -810 3818 -776 3852
rect -486 3818 -452 3852
rect -1547 3588 -1513 3622
rect -1187 3588 -1153 3622
rect -1067 3588 -1033 3622
rect -707 3588 -673 3622
rect -587 3588 -553 3622
rect 1032 3818 1066 3852
rect 1356 3818 1390 3852
rect 1510 3818 1544 3852
rect 1834 3818 1868 3852
rect 1992 3818 2026 3852
rect 1133 3588 1167 3622
rect 1253 3588 1287 3622
rect 1613 3588 1647 3622
rect 1733 3588 1767 3622
rect 2093 3588 2127 3622
rect 6450 3550 6490 3590
rect 6850 3550 6890 3590
rect -2050 3210 -2010 3250
rect -1810 3210 -1770 3250
rect -1570 3210 -1530 3250
rect -1330 3210 -1290 3250
rect -690 3210 -650 3250
rect -450 3210 -410 3250
rect -210 3210 -170 3250
rect 750 3210 790 3250
rect 990 3210 1030 3250
rect 1230 3210 1270 3250
rect 1870 3210 1910 3250
rect 2110 3210 2150 3250
rect 2350 3210 2390 3250
rect 2590 3210 2630 3250
rect -1650 2300 -1610 2340
rect -1490 2300 -1450 2340
rect -1330 2300 -1290 2340
rect -1170 2300 -1130 2340
rect -1010 2300 -970 2340
rect -850 2300 -810 2340
rect -690 2300 -650 2340
rect -530 2300 -490 2340
rect -370 2300 -330 2340
rect -210 2300 -170 2340
rect -50 2300 -10 2340
rect 110 2300 150 2340
rect 430 2300 470 2340
rect 590 2300 630 2340
rect 750 2300 790 2340
rect 910 2300 950 2340
rect 1070 2300 1110 2340
rect 1230 2300 1270 2340
rect 1390 2300 1430 2340
rect 1550 2300 1590 2340
rect 1710 2300 1750 2340
rect 1870 2300 1910 2340
rect 2030 2300 2070 2340
rect 2190 2300 2230 2340
<< xpolycontact >>
rect -358 1720 82 1790
rect 510 1720 950 1790
rect -2860 -962 -2790 -522
rect -2860 -1778 -2790 -1340
rect -2740 -910 -2670 -470
rect -2740 -1988 -2670 -1548
rect -2620 -910 -2550 -470
rect -2620 -1988 -2550 -1548
rect -2500 -910 -2430 -470
rect -2500 -1988 -2430 -1548
rect -2310 -530 -2240 -90
rect -2310 -2138 -2240 -1698
rect -2190 -530 -2120 -90
rect -2190 -2138 -2120 -1698
rect -2070 -530 -2000 -90
rect 2460 -530 2530 -90
rect -2070 -2138 -2000 -1698
rect 2460 -2138 2530 -1698
rect 2580 -530 2650 -90
rect 2580 -2138 2650 -1698
rect 2700 -530 2770 -90
rect 2700 -2138 2770 -1698
rect 2820 -1380 2890 -940
rect 3480 -1172 3550 -732
rect 2820 -1988 2890 -1548
rect 3480 -1988 3550 -1550
rect 2978 -2980 3418 -2910
rect 4890 -2980 5330 -2910
<< npolyres >>
rect 5784 6290 6264 6356
<< ppolyres >>
rect -2860 -1340 -2790 -962
rect 3480 -1550 3550 -1172
<< xpolyres >>
rect 82 1720 510 1790
rect -2740 -1548 -2670 -910
rect -2620 -1548 -2550 -910
rect -2500 -1548 -2430 -910
rect -2310 -1698 -2240 -530
rect -2190 -1698 -2120 -530
rect -2070 -1698 -2000 -530
rect 2460 -1698 2530 -530
rect 2580 -1698 2650 -530
rect 2700 -1698 2770 -530
rect 2820 -1548 2890 -1380
rect 3418 -2980 4890 -2910
<< locali >>
rect 9410 13890 9490 13910
rect 9930 13890 10010 13910
rect 10450 13890 10530 13910
rect 10940 13890 11020 13910
rect 9200 13850 9430 13890
rect 9470 13850 9950 13890
rect 9990 13850 10330 13890
rect 10510 13850 10960 13890
rect 11000 13850 11230 13890
rect 9200 13470 9240 13850
rect 9410 13830 9490 13850
rect 9930 13830 10010 13850
rect 10450 13830 10530 13850
rect 10940 13830 11020 13850
rect 9310 13760 9370 13780
rect 9310 13720 9320 13760
rect 9360 13720 9370 13760
rect 9310 13660 9370 13720
rect 9310 13620 9320 13660
rect 9360 13620 9370 13660
rect 9310 13600 9370 13620
rect 9420 13760 9480 13780
rect 9420 13720 9430 13760
rect 9470 13720 9480 13760
rect 9420 13660 9480 13720
rect 9420 13620 9430 13660
rect 9470 13620 9480 13660
rect 9420 13600 9480 13620
rect 9830 13760 9890 13780
rect 9830 13720 9840 13760
rect 9880 13720 9890 13760
rect 9830 13660 9890 13720
rect 9830 13620 9840 13660
rect 9880 13620 9890 13660
rect 9830 13600 9890 13620
rect 9940 13760 10000 13780
rect 9940 13720 9950 13760
rect 9990 13720 10000 13760
rect 9940 13660 10000 13720
rect 9940 13620 9950 13660
rect 9990 13620 10000 13660
rect 9940 13600 10000 13620
rect 10350 13760 10410 13780
rect 10350 13720 10360 13760
rect 10400 13720 10410 13760
rect 10350 13660 10410 13720
rect 10350 13620 10360 13660
rect 10400 13620 10410 13660
rect 10350 13600 10410 13620
rect 10460 13760 10520 13780
rect 10460 13720 10470 13760
rect 10510 13720 10520 13760
rect 10460 13660 10520 13720
rect 10460 13620 10470 13660
rect 10510 13620 10520 13660
rect 10460 13600 10520 13620
rect 10950 13760 11010 13780
rect 10950 13720 10960 13760
rect 11000 13720 11010 13760
rect 10950 13660 11010 13720
rect 10950 13620 10960 13660
rect 11000 13620 11010 13660
rect 10950 13600 11010 13620
rect 11060 13760 11120 13780
rect 11060 13720 11070 13760
rect 11110 13720 11120 13760
rect 11060 13660 11120 13720
rect 11060 13620 11070 13660
rect 11110 13620 11120 13660
rect 11060 13600 11120 13620
rect 9366 13542 9424 13560
rect 9366 13508 9378 13542
rect 9412 13508 9424 13542
rect 9366 13490 9424 13508
rect 9886 13542 9944 13560
rect 9886 13508 9898 13542
rect 9932 13508 9944 13542
rect 9886 13490 9944 13508
rect 10406 13542 10464 13560
rect 10406 13508 10418 13542
rect 10452 13508 10464 13542
rect 10406 13490 10464 13508
rect 10974 13542 11032 13560
rect 10974 13508 10986 13542
rect 11020 13508 11032 13542
rect 10974 13490 11032 13508
rect 11190 13470 11230 13850
rect 9310 13380 9370 13400
rect 9310 13340 9320 13380
rect 9360 13340 9370 13380
rect 9310 13280 9370 13340
rect 9310 13240 9320 13280
rect 9360 13240 9370 13280
rect 9310 13220 9370 13240
rect 9420 13380 9480 13400
rect 9420 13340 9430 13380
rect 9470 13340 9480 13380
rect 9420 13280 9480 13340
rect 9420 13240 9430 13280
rect 9470 13240 9480 13280
rect 9420 13220 9480 13240
rect 9830 13380 9890 13400
rect 9830 13340 9840 13380
rect 9880 13340 9890 13380
rect 9830 13280 9890 13340
rect 9830 13240 9840 13280
rect 9880 13240 9890 13280
rect 9830 13220 9890 13240
rect 9940 13380 10000 13400
rect 9940 13340 9950 13380
rect 9990 13340 10000 13380
rect 9940 13280 10000 13340
rect 9940 13240 9950 13280
rect 9990 13240 10000 13280
rect 9940 13220 10000 13240
rect 10350 13380 10410 13400
rect 10350 13340 10360 13380
rect 10400 13340 10410 13380
rect 10350 13280 10410 13340
rect 10350 13240 10360 13280
rect 10400 13240 10410 13280
rect 10350 13220 10410 13240
rect 10460 13380 10520 13400
rect 10460 13340 10470 13380
rect 10510 13340 10520 13380
rect 10460 13280 10520 13340
rect 10460 13240 10470 13280
rect 10510 13240 10520 13280
rect 10460 13220 10520 13240
rect -1350 13040 -1270 13060
rect -1350 13000 -1330 13040
rect -1290 13000 -1270 13040
rect -1350 12980 -1270 13000
rect -1130 13040 -1050 13060
rect -1130 13000 -1110 13040
rect -1070 13000 -1050 13040
rect -1130 12980 -1050 13000
rect -660 13040 -580 13060
rect -660 13000 -640 13040
rect -600 13000 -580 13040
rect -660 12980 -580 13000
rect -320 13040 -240 13060
rect -320 13000 -300 13040
rect -260 13000 -240 13040
rect -320 12980 -240 13000
rect -100 13040 -20 13060
rect -100 13000 -80 13040
rect -40 13000 -20 13040
rect -100 12980 -20 13000
rect 340 13040 420 13060
rect 340 13000 360 13040
rect 400 13000 420 13040
rect 340 12980 420 13000
rect 1020 13040 1100 13060
rect 1020 13000 1040 13040
rect 1080 13000 1100 13040
rect 1020 12980 1100 13000
rect 1240 13040 1320 13060
rect 1240 13000 1260 13040
rect 1300 13000 1320 13040
rect 1240 12980 1320 13000
rect 1710 13040 1790 13060
rect 1710 13000 1730 13040
rect 1770 13000 1790 13040
rect 1710 12980 1790 13000
rect 2170 13040 2250 13060
rect 2170 13000 2190 13040
rect 2230 13000 2250 13040
rect 2170 12980 2250 13000
rect 2520 13040 2600 13060
rect 2520 13000 2540 13040
rect 2580 13000 2600 13040
rect 2520 12980 2600 13000
rect 2770 13040 2850 13060
rect 2770 13000 2790 13040
rect 2830 13000 2850 13040
rect 2770 12980 2850 13000
rect 2990 13040 3070 13060
rect 2990 13000 3010 13040
rect 3050 13000 3070 13040
rect 2990 12980 3070 13000
rect 3320 13040 3400 13060
rect 3320 13000 3340 13040
rect 3380 13000 3400 13040
rect 3320 12980 3400 13000
rect 3980 13040 4060 13060
rect 3980 13000 4000 13040
rect 4040 13000 4060 13040
rect 3980 12980 4060 13000
rect 4200 13040 4280 13060
rect 4200 13000 4220 13040
rect 4260 13000 4280 13040
rect 4200 12980 4280 13000
rect 4770 13040 4850 13060
rect 4770 13000 4790 13040
rect 4830 13000 4850 13040
rect 4770 12980 4850 13000
rect 5030 13040 5110 13060
rect 5030 13000 5050 13040
rect 5090 13000 5110 13040
rect 5030 12980 5110 13000
rect 5280 13040 5360 13060
rect 5280 13000 5300 13040
rect 5340 13000 5360 13040
rect 5280 12980 5360 13000
rect 5500 13040 5580 13060
rect 5500 13000 5520 13040
rect 5560 13000 5580 13040
rect 5500 12980 5580 13000
rect 6050 13040 6130 13060
rect 6050 13000 6070 13040
rect 6110 13000 6130 13040
rect 6050 12980 6130 13000
rect 6330 13040 6410 13060
rect 6330 13000 6350 13040
rect 6390 13000 6410 13040
rect 6330 12980 6410 13000
rect 6580 13040 6660 13060
rect 6580 13000 6600 13040
rect 6640 13000 6660 13040
rect 6580 12980 6660 13000
rect 6800 13040 6880 13060
rect 6800 13000 6820 13040
rect 6860 13000 6880 13040
rect 6800 12980 6880 13000
rect 7350 13040 7430 13060
rect 7350 13000 7370 13040
rect 7410 13000 7430 13040
rect 7350 12980 7430 13000
rect 7630 13040 7710 13060
rect 7630 13000 7650 13040
rect 7690 13000 7710 13040
rect 7630 12980 7710 13000
rect 7880 13040 7960 13060
rect 7880 13000 7900 13040
rect 7940 13000 7960 13040
rect 7880 12980 7960 13000
rect 8100 13040 8180 13060
rect 8100 13000 8120 13040
rect 8160 13000 8180 13040
rect 8100 12980 8180 13000
rect 8650 13040 8730 13060
rect 8650 13000 8670 13040
rect 8710 13000 8730 13040
rect 8650 12980 8730 13000
rect -1510 12930 -1430 12950
rect -1510 12890 -1490 12930
rect -1450 12890 -1430 12930
rect -1510 12870 -1430 12890
rect -1490 12830 -1450 12870
rect -1330 12830 -1290 12980
rect -1110 12830 -1070 12980
rect -640 12830 -600 12980
rect -560 12910 -480 12930
rect -560 12870 -540 12910
rect -500 12870 -480 12910
rect -430 12920 -350 12940
rect -430 12880 -410 12920
rect -370 12880 -350 12920
rect -430 12870 -350 12880
rect -560 12850 -480 12870
rect -410 12830 -370 12870
rect -300 12830 -260 12980
rect -80 12830 -40 12980
rect 360 12830 400 12980
rect 510 12920 590 12940
rect 510 12880 530 12920
rect 570 12880 590 12920
rect 510 12870 590 12880
rect 1040 12830 1080 12980
rect 1260 12830 1300 12980
rect 1730 12830 1770 12980
rect 2070 12920 2150 12940
rect 2070 12880 2090 12920
rect 2130 12880 2150 12920
rect 2070 12870 2150 12880
rect 2190 12830 2230 12980
rect 2540 12830 2580 12980
rect 2790 12830 2830 12980
rect 3010 12830 3050 12980
rect 3340 12830 3380 12980
rect 4000 12830 4040 12980
rect 4220 12830 4260 12980
rect 4684 12930 4750 12950
rect 4684 12890 4694 12930
rect 4734 12890 4750 12930
rect 4684 12870 4750 12890
rect 4790 12830 4830 12980
rect 5050 12920 5090 12980
rect 5300 12920 5340 12980
rect 5520 12920 5560 12980
rect 6070 12920 6110 12980
rect 6350 12920 6390 12980
rect 6600 12920 6640 12980
rect 6820 12920 6860 12980
rect 7370 12920 7410 12980
rect 7650 12920 7690 12980
rect 7900 12920 7940 12980
rect 8120 12920 8160 12980
rect 8670 12920 8710 12980
rect 5040 12900 5100 12920
rect 5180 12900 5240 12920
rect 5040 12860 5050 12900
rect 5090 12860 5100 12900
rect 5040 12840 5100 12860
rect 5140 12860 5190 12900
rect 5230 12860 5240 12900
rect 5140 12840 5240 12860
rect 5290 12900 5350 12920
rect 5290 12860 5300 12900
rect 5340 12860 5350 12900
rect 5290 12840 5350 12860
rect 5400 12900 5460 12920
rect 5400 12860 5410 12900
rect 5450 12860 5460 12900
rect 5400 12840 5460 12860
rect 5510 12900 5570 12920
rect 5510 12860 5520 12900
rect 5560 12860 5570 12900
rect 5510 12840 5570 12860
rect 5620 12900 5680 12920
rect 5620 12860 5630 12900
rect 5670 12860 5680 12900
rect 5840 12900 5900 12920
rect 5840 12880 5850 12900
rect 5620 12840 5680 12860
rect 5720 12860 5850 12880
rect 5890 12860 5900 12900
rect 5720 12840 5900 12860
rect 5950 12900 6010 12920
rect 5950 12860 5960 12900
rect 6000 12860 6010 12900
rect 5950 12840 6010 12860
rect 6060 12900 6120 12920
rect 6060 12860 6070 12900
rect 6110 12860 6120 12900
rect 6060 12840 6120 12860
rect 6170 12900 6230 12920
rect 6170 12860 6180 12900
rect 6220 12860 6230 12900
rect 6170 12840 6230 12860
rect 6340 12900 6400 12920
rect 6480 12900 6540 12920
rect 6340 12860 6350 12900
rect 6390 12860 6400 12900
rect 6340 12840 6400 12860
rect 6440 12860 6490 12900
rect 6530 12860 6540 12900
rect 6440 12840 6540 12860
rect 6590 12900 6650 12920
rect 6590 12860 6600 12900
rect 6640 12860 6650 12900
rect 6590 12840 6650 12860
rect 6700 12900 6760 12920
rect 6700 12860 6710 12900
rect 6750 12860 6760 12900
rect 6700 12840 6760 12860
rect 6810 12900 6870 12920
rect 6810 12860 6820 12900
rect 6860 12860 6870 12900
rect 6810 12840 6870 12860
rect 6920 12900 6980 12920
rect 6920 12860 6930 12900
rect 6970 12860 6980 12900
rect 7140 12900 7200 12920
rect 7140 12880 7150 12900
rect 6920 12840 6980 12860
rect 7020 12860 7150 12880
rect 7190 12860 7200 12900
rect 7020 12840 7200 12860
rect 7250 12900 7310 12920
rect 7250 12860 7260 12900
rect 7300 12860 7310 12900
rect 7250 12840 7310 12860
rect 7360 12900 7420 12920
rect 7360 12860 7370 12900
rect 7410 12860 7420 12900
rect 7360 12840 7420 12860
rect 7470 12900 7530 12920
rect 7470 12860 7480 12900
rect 7520 12860 7530 12900
rect 7470 12840 7530 12860
rect 7640 12900 7700 12920
rect 7780 12900 7840 12920
rect 7640 12860 7650 12900
rect 7690 12860 7700 12900
rect 7640 12840 7700 12860
rect 7740 12860 7790 12900
rect 7830 12860 7840 12900
rect 7740 12840 7840 12860
rect 7890 12900 7950 12920
rect 7890 12860 7900 12900
rect 7940 12860 7950 12900
rect 7890 12840 7950 12860
rect 8000 12900 8060 12920
rect 8000 12860 8010 12900
rect 8050 12860 8060 12900
rect 8000 12840 8060 12860
rect 8110 12900 8170 12920
rect 8110 12860 8120 12900
rect 8160 12860 8170 12900
rect 8110 12840 8170 12860
rect 8220 12900 8280 12920
rect 8220 12860 8230 12900
rect 8270 12860 8280 12900
rect 8440 12900 8500 12920
rect 8440 12880 8450 12900
rect 8220 12840 8280 12860
rect 8320 12860 8450 12880
rect 8490 12860 8500 12900
rect 8320 12840 8500 12860
rect 8550 12900 8610 12920
rect 8550 12860 8560 12900
rect 8600 12860 8610 12900
rect 8550 12840 8610 12860
rect 8660 12900 8720 12920
rect 8660 12860 8670 12900
rect 8710 12860 8720 12900
rect 8660 12840 8720 12860
rect 8770 12900 8830 12920
rect 8770 12860 8780 12900
rect 8820 12860 8830 12900
rect 8770 12840 8830 12860
rect -1490 12810 -1390 12830
rect -1490 12770 -1440 12810
rect -1400 12770 -1390 12810
rect -1490 12750 -1390 12770
rect -1340 12810 -1280 12830
rect -1340 12770 -1330 12810
rect -1290 12770 -1280 12810
rect -1340 12750 -1280 12770
rect -1230 12810 -1170 12830
rect -1230 12770 -1220 12810
rect -1180 12770 -1170 12810
rect -1230 12750 -1170 12770
rect -1120 12810 -1060 12830
rect -1120 12770 -1110 12810
rect -1070 12770 -1060 12810
rect -1120 12750 -1060 12770
rect -1010 12810 -950 12830
rect -870 12810 -810 12830
rect -1010 12770 -1000 12810
rect -960 12770 -950 12810
rect -1010 12750 -950 12770
rect -910 12770 -860 12810
rect -820 12770 -810 12810
rect -910 12750 -810 12770
rect -760 12810 -700 12830
rect -760 12770 -750 12810
rect -710 12770 -700 12810
rect -760 12750 -700 12770
rect -650 12810 -590 12830
rect -650 12770 -640 12810
rect -600 12770 -590 12810
rect -650 12750 -590 12770
rect -420 12810 -360 12830
rect -420 12770 -410 12810
rect -370 12770 -360 12810
rect -420 12750 -360 12770
rect -310 12810 -250 12830
rect -310 12770 -300 12810
rect -260 12770 -250 12810
rect -310 12750 -250 12770
rect -200 12810 -140 12830
rect -200 12770 -190 12810
rect -150 12770 -140 12810
rect -200 12750 -140 12770
rect -90 12810 -30 12830
rect -90 12770 -80 12810
rect -40 12770 -30 12810
rect -90 12750 -30 12770
rect 20 12810 80 12830
rect 20 12770 30 12810
rect 70 12770 80 12810
rect 20 12750 80 12770
rect 240 12810 300 12830
rect 240 12770 250 12810
rect 290 12770 300 12810
rect 240 12750 300 12770
rect 350 12810 410 12830
rect 350 12770 360 12810
rect 400 12770 410 12810
rect 350 12750 410 12770
rect 460 12810 520 12830
rect 460 12770 470 12810
rect 510 12770 520 12810
rect 460 12750 520 12770
rect 570 12810 630 12830
rect 570 12770 580 12810
rect 620 12770 630 12810
rect 570 12750 630 12770
rect 680 12810 740 12830
rect 920 12810 980 12830
rect 680 12770 690 12810
rect 730 12770 780 12810
rect 680 12750 780 12770
rect -1490 12680 -1450 12750
rect -1220 12710 -1180 12750
rect -1000 12710 -960 12750
rect -1570 12660 -1450 12680
rect -1570 12620 -1550 12660
rect -1510 12620 -1450 12660
rect -1400 12690 -960 12710
rect -1400 12650 -1380 12690
rect -1340 12670 -960 12690
rect -1340 12650 -1320 12670
rect -1400 12630 -1320 12650
rect -1570 12600 -1450 12620
rect -1490 12510 -1450 12600
rect -1530 12490 -1450 12510
rect -1290 12490 -1230 12510
rect -1530 12450 -1510 12490
rect -1470 12450 -1280 12490
rect -1240 12450 -1230 12490
rect -1530 12430 -1450 12450
rect -1290 12430 -1230 12450
rect -1180 12490 -1040 12510
rect -1180 12450 -1170 12490
rect -1130 12450 -1090 12490
rect -1050 12450 -1040 12490
rect -1000 12490 -960 12670
rect -910 12590 -870 12750
rect -420 12710 -380 12750
rect -200 12710 -160 12750
rect 20 12710 60 12750
rect 250 12710 290 12750
rect 470 12710 510 12750
rect -820 12690 -740 12710
rect -480 12690 -380 12710
rect -820 12650 -800 12690
rect -760 12650 -460 12690
rect -420 12650 -380 12690
rect -820 12630 -740 12650
rect -480 12630 -380 12650
rect -240 12670 60 12710
rect -240 12630 -200 12670
rect -910 12550 -600 12590
rect -640 12510 -600 12550
rect -870 12490 -810 12510
rect -1000 12450 -860 12490
rect -820 12450 -810 12490
rect -1180 12430 -1040 12450
rect -870 12430 -810 12450
rect -760 12490 -700 12510
rect -760 12450 -750 12490
rect -710 12450 -700 12490
rect -760 12430 -700 12450
rect -650 12490 -590 12510
rect -650 12450 -640 12490
rect -600 12450 -590 12490
rect -420 12490 -380 12630
rect -280 12610 -200 12630
rect -280 12570 -260 12610
rect -220 12570 -200 12610
rect -280 12550 -200 12570
rect 20 12510 60 12670
rect 100 12690 180 12710
rect 100 12650 120 12690
rect 160 12650 180 12690
rect 250 12670 510 12710
rect 620 12690 700 12710
rect 100 12640 180 12650
rect 620 12650 640 12690
rect 680 12650 700 12690
rect 620 12640 700 12650
rect 740 12590 780 12750
rect 120 12570 780 12590
rect 120 12530 140 12570
rect 180 12550 780 12570
rect 880 12770 930 12810
rect 970 12770 980 12810
rect 880 12750 980 12770
rect 1030 12810 1090 12830
rect 1030 12770 1040 12810
rect 1080 12770 1090 12810
rect 1030 12750 1090 12770
rect 1140 12810 1200 12830
rect 1140 12770 1150 12810
rect 1190 12770 1200 12810
rect 1140 12750 1200 12770
rect 1250 12810 1310 12830
rect 1250 12770 1260 12810
rect 1300 12770 1310 12810
rect 1250 12750 1310 12770
rect 1360 12810 1420 12830
rect 1500 12810 1560 12830
rect 1360 12770 1370 12810
rect 1410 12770 1420 12810
rect 1360 12750 1420 12770
rect 1460 12770 1510 12810
rect 1550 12770 1560 12810
rect 1460 12750 1560 12770
rect 1610 12810 1670 12830
rect 1610 12770 1620 12810
rect 1660 12770 1670 12810
rect 1610 12750 1670 12770
rect 1720 12810 1860 12830
rect 2060 12810 2120 12830
rect 1720 12770 1730 12810
rect 1770 12770 1810 12810
rect 1850 12770 1860 12810
rect 1720 12750 1860 12770
rect 1900 12770 2070 12810
rect 2110 12770 2120 12810
rect 180 12530 200 12550
rect 120 12510 200 12530
rect 250 12510 290 12550
rect 580 12510 620 12550
rect 880 12510 920 12750
rect 1150 12710 1190 12750
rect 1370 12710 1410 12750
rect 970 12690 1410 12710
rect 970 12650 990 12690
rect 1030 12670 1410 12690
rect 1030 12650 1050 12670
rect 970 12640 1050 12650
rect -200 12490 -140 12510
rect -420 12450 -190 12490
rect -150 12450 -140 12490
rect -650 12430 -590 12450
rect -200 12430 -140 12450
rect -90 12490 -30 12510
rect -90 12450 -80 12490
rect -40 12450 -30 12490
rect -90 12430 -30 12450
rect 20 12490 80 12510
rect 20 12450 30 12490
rect 70 12450 80 12490
rect 20 12430 80 12450
rect 240 12490 300 12510
rect 240 12450 250 12490
rect 290 12450 300 12490
rect 240 12430 300 12450
rect 350 12490 410 12510
rect 350 12450 360 12490
rect 400 12450 410 12490
rect 350 12430 410 12450
rect 460 12490 530 12510
rect 460 12450 470 12490
rect 510 12450 530 12490
rect 460 12430 530 12450
rect 570 12490 630 12510
rect 570 12450 580 12490
rect 620 12450 630 12490
rect 570 12430 630 12450
rect 840 12490 920 12510
rect 1080 12490 1140 12510
rect 840 12450 860 12490
rect 900 12450 1090 12490
rect 1130 12450 1140 12490
rect 840 12430 920 12450
rect 1080 12430 1140 12450
rect 1190 12490 1330 12510
rect 1190 12450 1200 12490
rect 1240 12450 1280 12490
rect 1320 12450 1330 12490
rect 1370 12490 1410 12670
rect 1460 12590 1500 12750
rect 1550 12690 1630 12710
rect 1760 12690 1840 12710
rect 1550 12650 1570 12690
rect 1610 12650 1780 12690
rect 1820 12650 1840 12690
rect 1550 12630 1630 12650
rect 1760 12640 1840 12650
rect 1900 12590 1940 12770
rect 2060 12750 2120 12770
rect 2170 12810 2230 12830
rect 2170 12770 2180 12810
rect 2220 12770 2230 12810
rect 2170 12750 2230 12770
rect 2420 12810 2480 12830
rect 2420 12770 2430 12810
rect 2470 12770 2480 12810
rect 2420 12750 2480 12770
rect 2530 12810 2590 12830
rect 2530 12770 2540 12810
rect 2580 12770 2590 12810
rect 2530 12750 2590 12770
rect 2670 12810 2730 12830
rect 2670 12770 2680 12810
rect 2720 12770 2730 12810
rect 2670 12750 2730 12770
rect 2780 12810 2840 12830
rect 2780 12770 2790 12810
rect 2830 12770 2840 12810
rect 2780 12750 2840 12770
rect 2890 12810 2950 12830
rect 2890 12770 2900 12810
rect 2940 12770 2950 12810
rect 2890 12750 2950 12770
rect 3000 12810 3060 12830
rect 3000 12770 3010 12810
rect 3050 12770 3060 12810
rect 3000 12750 3060 12770
rect 3110 12810 3170 12830
rect 3110 12770 3120 12810
rect 3160 12770 3170 12810
rect 3110 12750 3170 12770
rect 3250 12810 3390 12830
rect 3250 12770 3260 12810
rect 3300 12770 3340 12810
rect 3380 12770 3390 12810
rect 3250 12750 3390 12770
rect 3440 12810 3500 12830
rect 3440 12770 3450 12810
rect 3490 12770 3500 12810
rect 3440 12750 3500 12770
rect 3550 12810 3610 12830
rect 3550 12770 3560 12810
rect 3600 12770 3610 12810
rect 3550 12750 3610 12770
rect 3660 12810 3720 12830
rect 3880 12810 3940 12830
rect 3660 12770 3670 12810
rect 3710 12770 3760 12810
rect 3660 12750 3760 12770
rect 2000 12690 2080 12710
rect 2430 12700 2470 12750
rect 2000 12650 2020 12690
rect 2060 12670 2080 12690
rect 2340 12680 2470 12700
rect 2340 12670 2360 12680
rect 2060 12650 2360 12670
rect 2000 12640 2360 12650
rect 2400 12640 2470 12680
rect 2670 12660 2710 12750
rect 2890 12710 2930 12750
rect 3110 12710 3150 12750
rect 2000 12630 2470 12640
rect 2340 12620 2470 12630
rect 1460 12550 1770 12590
rect 1730 12510 1770 12550
rect 1820 12570 2220 12590
rect 1820 12530 1840 12570
rect 1880 12550 2220 12570
rect 1880 12530 1900 12550
rect 1820 12510 1900 12530
rect 1960 12510 2000 12550
rect 2180 12510 2220 12550
rect 2430 12510 2470 12620
rect 2610 12640 2710 12660
rect 2610 12600 2630 12640
rect 2670 12600 2710 12640
rect 2850 12670 3150 12710
rect 2850 12630 2890 12670
rect 2610 12580 2710 12600
rect 1500 12490 1560 12510
rect 1370 12450 1510 12490
rect 1550 12450 1560 12490
rect 1190 12430 1330 12450
rect 1500 12430 1560 12450
rect 1610 12490 1670 12510
rect 1610 12450 1620 12490
rect 1660 12450 1670 12490
rect 1610 12430 1670 12450
rect 1720 12490 1780 12510
rect 1720 12450 1730 12490
rect 1770 12450 1780 12490
rect 1720 12430 1780 12450
rect 1950 12490 2010 12510
rect 1950 12450 1960 12490
rect 2000 12450 2010 12490
rect 1950 12430 2010 12450
rect 2060 12490 2120 12510
rect 2060 12450 2070 12490
rect 2110 12450 2120 12490
rect 2060 12430 2120 12450
rect 2170 12490 2230 12510
rect 2170 12450 2180 12490
rect 2220 12450 2230 12490
rect 2170 12430 2230 12450
rect 2310 12490 2370 12510
rect 2310 12450 2320 12490
rect 2360 12450 2370 12490
rect 2310 12430 2370 12450
rect 2420 12490 2480 12510
rect 2420 12450 2430 12490
rect 2470 12450 2480 12490
rect 2420 12430 2480 12450
rect 2530 12490 2590 12510
rect 2530 12450 2540 12490
rect 2580 12450 2590 12490
rect 2670 12490 2710 12580
rect 2810 12610 2890 12630
rect 2810 12570 2830 12610
rect 2870 12570 2890 12610
rect 2810 12550 2890 12570
rect 3110 12510 3150 12670
rect 3240 12690 3320 12710
rect 3600 12690 3680 12710
rect 3240 12650 3260 12690
rect 3300 12650 3620 12690
rect 3660 12650 3680 12690
rect 3240 12640 3320 12650
rect 3600 12640 3680 12650
rect 3210 12570 3600 12590
rect 3210 12530 3230 12570
rect 3270 12550 3600 12570
rect 3270 12530 3290 12550
rect 3210 12510 3290 12530
rect 3340 12510 3380 12550
rect 3560 12510 3600 12550
rect 2890 12490 2950 12510
rect 2670 12450 2900 12490
rect 2940 12450 2950 12490
rect 2530 12430 2590 12450
rect 2890 12430 2950 12450
rect 3000 12490 3060 12510
rect 3000 12450 3010 12490
rect 3050 12450 3060 12490
rect 3000 12430 3060 12450
rect 3110 12490 3170 12510
rect 3110 12450 3120 12490
rect 3160 12450 3170 12490
rect 3110 12430 3170 12450
rect 3330 12490 3390 12510
rect 3330 12450 3340 12490
rect 3380 12450 3390 12490
rect 3330 12430 3390 12450
rect 3440 12490 3500 12510
rect 3440 12450 3450 12490
rect 3490 12450 3500 12490
rect 3440 12430 3500 12450
rect 3550 12490 3610 12510
rect 3720 12490 3760 12750
rect 3840 12770 3890 12810
rect 3930 12770 3940 12810
rect 3840 12750 3940 12770
rect 3990 12810 4050 12830
rect 3990 12770 4000 12810
rect 4040 12770 4050 12810
rect 3990 12750 4050 12770
rect 4100 12810 4160 12830
rect 4100 12770 4110 12810
rect 4150 12770 4160 12810
rect 4100 12750 4160 12770
rect 4210 12810 4270 12830
rect 4210 12770 4220 12810
rect 4260 12770 4270 12810
rect 4210 12750 4270 12770
rect 4320 12810 4380 12830
rect 4320 12770 4330 12810
rect 4370 12770 4380 12810
rect 4540 12810 4600 12830
rect 4540 12790 4550 12810
rect 4320 12750 4380 12770
rect 4420 12770 4550 12790
rect 4590 12770 4600 12810
rect 4420 12750 4600 12770
rect 4650 12810 4710 12830
rect 4650 12770 4660 12810
rect 4700 12770 4710 12810
rect 4650 12750 4710 12770
rect 4760 12810 4830 12830
rect 4760 12770 4770 12810
rect 4810 12770 4830 12810
rect 4760 12750 4830 12770
rect 4870 12810 4930 12830
rect 4870 12770 4880 12810
rect 4920 12770 4930 12810
rect 4870 12750 4930 12770
rect 3840 12510 3880 12750
rect 4110 12710 4150 12750
rect 4330 12710 4370 12750
rect 3930 12690 4370 12710
rect 3930 12650 3950 12690
rect 3990 12670 4370 12690
rect 3990 12650 4010 12670
rect 3930 12640 4010 12650
rect 4260 12510 4300 12670
rect 4420 12630 4460 12750
rect 4880 12710 4920 12750
rect 4510 12690 4920 12710
rect 4510 12650 4530 12690
rect 4570 12670 4920 12690
rect 4570 12650 4590 12670
rect 4510 12630 4590 12650
rect 4340 12610 4460 12630
rect 4340 12570 4360 12610
rect 4400 12590 4460 12610
rect 4400 12570 4560 12590
rect 4340 12550 4560 12570
rect 4520 12510 4560 12550
rect 4660 12510 4700 12670
rect 4880 12510 4920 12670
rect 4980 12670 5060 12690
rect 4980 12630 5000 12670
rect 5040 12650 5060 12670
rect 5140 12650 5180 12840
rect 5410 12800 5450 12840
rect 5630 12800 5670 12840
rect 5230 12780 5670 12800
rect 5230 12740 5250 12780
rect 5290 12760 5670 12780
rect 5290 12740 5310 12760
rect 5230 12720 5310 12740
rect 5040 12630 5180 12650
rect 4980 12610 5180 12630
rect 3550 12450 3560 12490
rect 3600 12450 3760 12490
rect 3800 12490 3880 12510
rect 3950 12490 4010 12510
rect 3800 12450 3820 12490
rect 3860 12450 3960 12490
rect 4000 12450 4010 12490
rect 3550 12430 3610 12450
rect 3800 12430 3880 12450
rect 3950 12430 4010 12450
rect 4060 12490 4200 12510
rect 4060 12450 4070 12490
rect 4110 12450 4150 12490
rect 4190 12450 4200 12490
rect 4060 12430 4200 12450
rect 4260 12490 4350 12510
rect 4260 12450 4300 12490
rect 4340 12450 4350 12490
rect 4260 12430 4350 12450
rect 4400 12490 4460 12510
rect 4400 12450 4410 12490
rect 4450 12450 4460 12490
rect 4400 12430 4460 12450
rect 4510 12490 4570 12510
rect 4510 12450 4520 12490
rect 4560 12450 4570 12490
rect 4510 12430 4570 12450
rect 4650 12490 4710 12510
rect 4650 12450 4660 12490
rect 4700 12450 4710 12490
rect 4650 12430 4710 12450
rect 4760 12490 4820 12510
rect 4760 12450 4770 12490
rect 4810 12450 4820 12490
rect 4760 12430 4820 12450
rect 4870 12490 4930 12510
rect 4870 12450 4880 12490
rect 4920 12450 4930 12490
rect 5140 12490 5180 12610
rect 5560 12510 5600 12760
rect 5720 12630 5760 12840
rect 6180 12800 6220 12840
rect 5810 12780 6220 12800
rect 5810 12740 5830 12780
rect 5870 12760 6220 12780
rect 5870 12740 5890 12760
rect 5810 12720 5890 12740
rect 5640 12610 5760 12630
rect 5640 12570 5660 12610
rect 5700 12590 5760 12610
rect 5700 12570 5860 12590
rect 5640 12550 5860 12570
rect 5820 12510 5860 12550
rect 5960 12510 6000 12760
rect 6180 12510 6220 12760
rect 6280 12670 6360 12690
rect 6280 12630 6300 12670
rect 6340 12650 6360 12670
rect 6440 12650 6480 12840
rect 6710 12800 6750 12840
rect 6930 12800 6970 12840
rect 6530 12780 6970 12800
rect 6530 12740 6550 12780
rect 6590 12760 6970 12780
rect 6590 12740 6610 12760
rect 6530 12720 6610 12740
rect 6340 12630 6480 12650
rect 6280 12610 6480 12630
rect 5250 12490 5310 12510
rect 5140 12450 5260 12490
rect 5300 12450 5310 12490
rect 4870 12430 4930 12450
rect 5250 12430 5310 12450
rect 5360 12490 5500 12510
rect 5360 12450 5370 12490
rect 5410 12450 5450 12490
rect 5490 12450 5500 12490
rect 5360 12430 5500 12450
rect 5560 12490 5650 12510
rect 5560 12450 5600 12490
rect 5640 12450 5650 12490
rect 5560 12430 5650 12450
rect 5700 12490 5760 12510
rect 5700 12450 5710 12490
rect 5750 12450 5760 12490
rect 5700 12430 5760 12450
rect 5810 12490 5870 12510
rect 5810 12450 5820 12490
rect 5860 12450 5870 12490
rect 5810 12430 5870 12450
rect 5950 12490 6010 12510
rect 5950 12450 5960 12490
rect 6000 12450 6010 12490
rect 5950 12430 6010 12450
rect 6060 12490 6120 12510
rect 6060 12450 6070 12490
rect 6110 12450 6120 12490
rect 6060 12430 6120 12450
rect 6170 12490 6230 12510
rect 6170 12450 6180 12490
rect 6220 12450 6230 12490
rect 6440 12490 6480 12610
rect 6860 12510 6900 12760
rect 7020 12630 7060 12840
rect 7480 12800 7520 12840
rect 7110 12780 7520 12800
rect 7110 12740 7130 12780
rect 7170 12760 7520 12780
rect 7170 12740 7190 12760
rect 7110 12720 7190 12740
rect 6940 12610 7060 12630
rect 6940 12570 6960 12610
rect 7000 12590 7060 12610
rect 7000 12570 7160 12590
rect 6940 12550 7160 12570
rect 7120 12510 7160 12550
rect 7260 12510 7300 12760
rect 7480 12510 7520 12760
rect 7580 12670 7660 12690
rect 7580 12630 7600 12670
rect 7640 12650 7660 12670
rect 7740 12650 7780 12840
rect 8010 12800 8050 12840
rect 8230 12800 8270 12840
rect 7830 12780 8270 12800
rect 7830 12740 7850 12780
rect 7890 12760 8270 12780
rect 7890 12740 7910 12760
rect 7830 12720 7910 12740
rect 7640 12630 7780 12650
rect 7580 12610 7780 12630
rect 6550 12490 6610 12510
rect 6440 12450 6560 12490
rect 6600 12450 6610 12490
rect 6170 12430 6230 12450
rect 6550 12430 6610 12450
rect 6660 12490 6800 12510
rect 6660 12450 6670 12490
rect 6710 12450 6750 12490
rect 6790 12450 6800 12490
rect 6660 12430 6800 12450
rect 6860 12490 6950 12510
rect 6860 12450 6900 12490
rect 6940 12450 6950 12490
rect 6860 12430 6950 12450
rect 7000 12490 7060 12510
rect 7000 12450 7010 12490
rect 7050 12450 7060 12490
rect 7000 12430 7060 12450
rect 7110 12490 7170 12510
rect 7110 12450 7120 12490
rect 7160 12450 7170 12490
rect 7110 12430 7170 12450
rect 7250 12490 7310 12510
rect 7250 12450 7260 12490
rect 7300 12450 7310 12490
rect 7250 12430 7310 12450
rect 7360 12490 7420 12510
rect 7360 12450 7370 12490
rect 7410 12450 7420 12490
rect 7360 12430 7420 12450
rect 7470 12490 7530 12510
rect 7470 12450 7480 12490
rect 7520 12450 7530 12490
rect 7740 12490 7780 12610
rect 8160 12510 8200 12760
rect 8320 12630 8360 12840
rect 8780 12800 8820 12840
rect 8410 12780 8820 12800
rect 8410 12740 8430 12780
rect 8470 12760 8820 12780
rect 8470 12740 8490 12760
rect 8410 12720 8490 12740
rect 8240 12610 8360 12630
rect 8240 12570 8260 12610
rect 8300 12590 8360 12610
rect 8300 12570 8460 12590
rect 8240 12550 8460 12570
rect 8420 12510 8460 12550
rect 8560 12510 8600 12760
rect 8780 12510 8820 12760
rect 9200 12770 9240 13210
rect 9380 13162 9438 13180
rect 9380 13128 9392 13162
rect 9426 13128 9438 13162
rect 9380 13110 9438 13128
rect 9900 13162 9958 13180
rect 9900 13128 9912 13162
rect 9946 13128 9958 13162
rect 9900 13110 9958 13128
rect 10420 13162 10478 13180
rect 10420 13128 10432 13162
rect 10466 13128 10478 13162
rect 10420 13110 10478 13128
rect 9310 13000 9370 13020
rect 9310 12960 9320 13000
rect 9360 12960 9370 13000
rect 9310 12940 9370 12960
rect 9420 13000 9480 13020
rect 9420 12960 9430 13000
rect 9470 12960 9480 13000
rect 9420 12940 9480 12960
rect 9830 13000 9890 13020
rect 9830 12960 9840 13000
rect 9880 12960 9890 13000
rect 9830 12940 9890 12960
rect 9940 13000 10000 13020
rect 9940 12960 9950 13000
rect 9990 12960 10000 13000
rect 9940 12940 10000 12960
rect 10350 13000 10410 13020
rect 10350 12960 10360 13000
rect 10400 12960 10410 13000
rect 10350 12940 10410 12960
rect 10460 13000 10520 13020
rect 10460 12960 10470 13000
rect 10510 12960 10520 13000
rect 10460 12940 10520 12960
rect 9352 12882 9410 12900
rect 9352 12848 9364 12882
rect 9398 12848 9410 12882
rect 9352 12830 9410 12848
rect 9872 12882 9930 12900
rect 9872 12848 9884 12882
rect 9918 12848 9930 12882
rect 9872 12830 9930 12848
rect 10392 12882 10450 12900
rect 10392 12848 10404 12882
rect 10438 12848 10450 12882
rect 10392 12830 10450 12848
rect 11190 12770 11230 13210
rect 9200 12730 10330 12770
rect 10470 12730 11230 12770
rect 8862 12662 8920 12690
rect 8862 12628 8874 12662
rect 8908 12628 8920 12662
rect 8862 12610 8920 12628
rect 9200 12530 10210 12570
rect 10370 12530 11420 12570
rect 7850 12490 7910 12510
rect 7740 12450 7860 12490
rect 7900 12450 7910 12490
rect 7470 12430 7530 12450
rect 7850 12430 7910 12450
rect 7960 12490 8100 12510
rect 7960 12450 7970 12490
rect 8010 12450 8050 12490
rect 8090 12450 8100 12490
rect 7960 12430 8100 12450
rect 8160 12490 8250 12510
rect 8160 12450 8200 12490
rect 8240 12450 8250 12490
rect 8160 12430 8250 12450
rect 8300 12490 8360 12510
rect 8300 12450 8310 12490
rect 8350 12450 8360 12490
rect 8300 12430 8360 12450
rect 8410 12490 8470 12510
rect 8410 12450 8420 12490
rect 8460 12450 8470 12490
rect 8410 12430 8470 12450
rect 8550 12490 8610 12510
rect 8550 12450 8560 12490
rect 8600 12450 8610 12490
rect 8550 12430 8610 12450
rect 8660 12490 8720 12510
rect 8660 12450 8670 12490
rect 8710 12450 8720 12490
rect 8660 12430 8720 12450
rect 8770 12490 8830 12510
rect 8770 12450 8780 12490
rect 8820 12450 8830 12490
rect 8770 12430 8830 12450
rect -1170 12280 -1130 12430
rect -870 12370 -790 12390
rect -870 12330 -850 12370
rect -810 12330 -790 12370
rect -870 12310 -790 12330
rect -750 12280 -710 12430
rect -640 12390 -600 12430
rect -670 12370 -600 12390
rect -670 12330 -660 12370
rect -620 12330 -600 12370
rect -560 12390 -480 12410
rect -560 12350 -540 12390
rect -500 12350 -480 12390
rect -560 12330 -480 12350
rect -670 12310 -600 12330
rect -80 12280 -40 12430
rect 250 12370 330 12390
rect 250 12330 270 12370
rect 310 12330 330 12370
rect 250 12310 330 12330
rect 390 12370 450 12390
rect 390 12330 400 12370
rect 440 12330 450 12370
rect 390 12310 450 12330
rect 490 12280 530 12430
rect 1200 12280 1240 12430
rect 1510 12370 1590 12390
rect 1510 12330 1530 12370
rect 1570 12330 1590 12370
rect 1510 12310 1590 12330
rect 1630 12280 1670 12430
rect 1730 12390 1770 12430
rect 1730 12370 1810 12390
rect 1730 12330 1750 12370
rect 1790 12330 1810 12370
rect 1730 12310 1810 12330
rect 2070 12280 2110 12430
rect 2320 12280 2360 12430
rect 2540 12280 2580 12430
rect 2900 12380 2940 12430
rect 2860 12360 2940 12380
rect 2860 12320 2880 12360
rect 2920 12320 2940 12360
rect 2860 12310 2940 12320
rect 3010 12280 3050 12430
rect 3270 12360 3350 12380
rect 3270 12320 3290 12360
rect 3330 12320 3350 12360
rect 3270 12310 3350 12320
rect 3450 12280 3490 12430
rect 4070 12280 4110 12430
rect 4410 12280 4450 12430
rect 4770 12280 4810 12430
rect 5260 12390 5300 12430
rect 5220 12370 5300 12390
rect 5220 12330 5240 12370
rect 5280 12330 5300 12370
rect 5220 12310 5300 12330
rect 5370 12280 5410 12430
rect 5710 12280 5750 12430
rect 5800 12370 5880 12390
rect 5800 12330 5820 12370
rect 5860 12330 5880 12370
rect 5800 12310 5880 12330
rect 6070 12280 6110 12430
rect 6560 12390 6600 12430
rect 6520 12370 6600 12390
rect 6520 12330 6540 12370
rect 6580 12330 6600 12370
rect 6520 12310 6600 12330
rect 6670 12280 6710 12430
rect 7010 12280 7050 12430
rect 7100 12370 7180 12390
rect 7100 12330 7120 12370
rect 7160 12330 7180 12370
rect 7100 12310 7180 12330
rect 7370 12280 7410 12430
rect 7860 12390 7900 12430
rect 7820 12370 7900 12390
rect 7820 12330 7840 12370
rect 7880 12330 7900 12370
rect 7820 12310 7900 12330
rect 7970 12280 8010 12430
rect 8310 12280 8350 12430
rect 8400 12370 8480 12390
rect 8400 12330 8420 12370
rect 8460 12330 8480 12370
rect 8400 12310 8480 12330
rect 8670 12280 8710 12430
rect -1190 12260 -1110 12280
rect -1190 12220 -1170 12260
rect -1130 12220 -1110 12260
rect -1190 12200 -1110 12220
rect -770 12260 -690 12280
rect -770 12220 -750 12260
rect -710 12220 -690 12260
rect -770 12200 -690 12220
rect -100 12260 -20 12280
rect -100 12220 -80 12260
rect -40 12220 -20 12260
rect -100 12200 -20 12220
rect 470 12260 550 12280
rect 470 12220 490 12260
rect 530 12220 550 12260
rect 470 12200 550 12220
rect 1180 12260 1260 12280
rect 1180 12220 1200 12260
rect 1240 12220 1260 12260
rect 1180 12200 1260 12220
rect 1610 12260 1690 12280
rect 1610 12220 1630 12260
rect 1670 12220 1690 12260
rect 1610 12200 1690 12220
rect 2050 12260 2130 12280
rect 2050 12220 2070 12260
rect 2110 12220 2130 12260
rect 2050 12200 2130 12220
rect 2300 12260 2380 12280
rect 2300 12220 2320 12260
rect 2360 12220 2380 12260
rect 2300 12200 2380 12220
rect 2520 12260 2600 12280
rect 2520 12220 2540 12260
rect 2580 12220 2600 12260
rect 2520 12200 2600 12220
rect 2990 12260 3070 12280
rect 2990 12220 3010 12260
rect 3050 12220 3070 12260
rect 2990 12200 3070 12220
rect 3430 12260 3510 12280
rect 3430 12220 3450 12260
rect 3490 12220 3510 12260
rect 3430 12200 3510 12220
rect 4050 12260 4130 12280
rect 4050 12220 4070 12260
rect 4110 12220 4130 12260
rect 4050 12200 4130 12220
rect 4390 12260 4470 12280
rect 4390 12220 4410 12260
rect 4450 12220 4470 12260
rect 4390 12200 4470 12220
rect 4750 12260 4830 12280
rect 4750 12220 4770 12260
rect 4810 12220 4830 12260
rect 4750 12200 4830 12220
rect 5350 12260 5430 12280
rect 5350 12220 5370 12260
rect 5410 12220 5430 12260
rect 5350 12200 5430 12220
rect 5690 12260 5770 12280
rect 5690 12220 5710 12260
rect 5750 12220 5770 12260
rect 5690 12200 5770 12220
rect 6050 12260 6130 12280
rect 6050 12220 6070 12260
rect 6110 12220 6130 12260
rect 6050 12200 6130 12220
rect 6650 12260 6730 12280
rect 6650 12220 6670 12260
rect 6710 12220 6730 12260
rect 6650 12200 6730 12220
rect 6990 12260 7070 12280
rect 6990 12220 7010 12260
rect 7050 12220 7070 12260
rect 6990 12200 7070 12220
rect 7350 12260 7430 12280
rect 7350 12220 7370 12260
rect 7410 12220 7430 12260
rect 7350 12200 7430 12220
rect 7950 12260 8030 12280
rect 7950 12220 7970 12260
rect 8010 12220 8030 12260
rect 7950 12200 8030 12220
rect 8290 12260 8370 12280
rect 8290 12220 8310 12260
rect 8350 12220 8370 12260
rect 8290 12200 8370 12220
rect 8650 12260 8730 12280
rect 8650 12220 8670 12260
rect 8710 12220 8730 12260
rect 8650 12200 8730 12220
rect 9200 11600 9240 12530
rect 9352 12452 9410 12470
rect 9352 12418 9364 12452
rect 9398 12418 9410 12452
rect 9352 12400 9410 12418
rect 9872 12452 9930 12470
rect 9872 12418 9884 12452
rect 9918 12418 9930 12452
rect 9872 12400 9930 12418
rect 10392 12452 10450 12470
rect 10392 12418 10404 12452
rect 10438 12418 10450 12452
rect 10392 12400 10450 12418
rect 9310 12340 9370 12360
rect 9310 12300 9320 12340
rect 9360 12300 9370 12340
rect 9310 12240 9370 12300
rect 9310 12200 9320 12240
rect 9360 12200 9370 12240
rect 9310 12180 9370 12200
rect 9420 12340 9480 12360
rect 9420 12300 9430 12340
rect 9470 12300 9480 12340
rect 9420 12240 9480 12300
rect 9420 12200 9430 12240
rect 9470 12200 9480 12240
rect 9420 12180 9480 12200
rect 9830 12340 9890 12360
rect 9830 12300 9840 12340
rect 9880 12300 9890 12340
rect 9830 12240 9890 12300
rect 9830 12200 9840 12240
rect 9880 12200 9890 12240
rect 9830 12180 9890 12200
rect 9940 12340 10000 12360
rect 9940 12300 9950 12340
rect 9990 12300 10000 12340
rect 9940 12240 10000 12300
rect 9940 12200 9950 12240
rect 9990 12200 10000 12240
rect 9940 12180 10000 12200
rect 10350 12340 10410 12360
rect 10350 12300 10360 12340
rect 10400 12300 10410 12340
rect 10350 12240 10410 12300
rect 10350 12200 10360 12240
rect 10400 12200 10410 12240
rect 10350 12180 10410 12200
rect 10460 12340 10520 12360
rect 10460 12300 10470 12340
rect 10510 12300 10520 12340
rect 10460 12240 10520 12300
rect 10460 12200 10470 12240
rect 10510 12200 10520 12240
rect 10460 12180 10520 12200
rect 9380 12072 9438 12090
rect 9380 12038 9392 12072
rect 9426 12038 9438 12072
rect 9380 12020 9438 12038
rect 9900 12072 9958 12090
rect 9900 12038 9912 12072
rect 9946 12038 9958 12072
rect 9900 12020 9958 12038
rect 10420 12072 10478 12090
rect 10420 12038 10432 12072
rect 10466 12038 10478 12072
rect 10420 12020 10478 12038
rect 9310 11960 9370 11980
rect 9310 11920 9320 11960
rect 9360 11920 9370 11960
rect 9310 11860 9370 11920
rect 9310 11820 9320 11860
rect 9360 11820 9370 11860
rect 9310 11760 9370 11820
rect 9310 11720 9320 11760
rect 9360 11720 9370 11760
rect 9310 11660 9370 11720
rect 9310 11620 9320 11660
rect 9360 11620 9370 11660
rect 9310 11600 9370 11620
rect 9420 11960 9480 11980
rect 9420 11920 9430 11960
rect 9470 11920 9480 11960
rect 9420 11860 9480 11920
rect 9420 11820 9430 11860
rect 9470 11820 9480 11860
rect 9420 11760 9480 11820
rect 9420 11720 9430 11760
rect 9470 11720 9480 11760
rect 9420 11660 9480 11720
rect 9420 11620 9430 11660
rect 9470 11620 9480 11660
rect 9420 11600 9480 11620
rect 9830 11960 9890 11980
rect 9830 11920 9840 11960
rect 9880 11920 9890 11960
rect 9830 11860 9890 11920
rect 9830 11820 9840 11860
rect 9880 11820 9890 11860
rect 9830 11760 9890 11820
rect 9830 11720 9840 11760
rect 9880 11720 9890 11760
rect 9830 11660 9890 11720
rect 9830 11620 9840 11660
rect 9880 11620 9890 11660
rect 9830 11600 9890 11620
rect 9940 11960 10000 11980
rect 9940 11920 9950 11960
rect 9990 11920 10000 11960
rect 9940 11860 10000 11920
rect 9940 11820 9950 11860
rect 9990 11820 10000 11860
rect 9940 11760 10000 11820
rect 9940 11720 9950 11760
rect 9990 11720 10000 11760
rect 9940 11660 10000 11720
rect 9940 11620 9950 11660
rect 9990 11620 10000 11660
rect 9940 11600 10000 11620
rect 10350 11960 10410 11980
rect 10350 11920 10360 11960
rect 10400 11920 10410 11960
rect 10350 11860 10410 11920
rect 10350 11820 10360 11860
rect 10400 11820 10410 11860
rect 10350 11760 10410 11820
rect 10350 11720 10360 11760
rect 10400 11720 10410 11760
rect 10350 11660 10410 11720
rect 10350 11620 10360 11660
rect 10400 11620 10410 11660
rect 10350 11600 10410 11620
rect 10460 11960 10520 11980
rect 10460 11920 10470 11960
rect 10510 11920 10520 11960
rect 10460 11860 10520 11920
rect 10460 11820 10470 11860
rect 10510 11820 10520 11860
rect 10460 11760 10520 11820
rect 10460 11720 10470 11760
rect 10510 11720 10520 11760
rect 10460 11660 10520 11720
rect 10460 11620 10470 11660
rect 10510 11620 10520 11660
rect 10460 11600 10520 11620
rect 11380 11600 11420 12530
rect 9490 11390 9570 11410
rect 9490 11350 9510 11390
rect 9550 11350 9570 11390
rect 9490 11330 9570 11350
rect 10010 11390 10090 11410
rect 10010 11350 10030 11390
rect 10070 11350 10090 11390
rect 10010 11330 10090 11350
rect 10530 11390 10610 11410
rect 10530 11350 10550 11390
rect 10590 11350 10610 11390
rect 10530 11330 10610 11350
rect 11060 11390 11120 11410
rect 11060 11350 11070 11390
rect 11110 11350 11120 11390
rect 11060 11330 11120 11350
rect 9200 10840 9240 11270
rect 9310 11270 9370 11290
rect 9310 11230 9320 11270
rect 9360 11230 9370 11270
rect 9310 11170 9370 11230
rect 9310 11130 9320 11170
rect 9360 11130 9370 11170
rect 9310 11070 9370 11130
rect 9310 11030 9320 11070
rect 9360 11030 9370 11070
rect 9310 10970 9370 11030
rect 9310 10930 9320 10970
rect 9360 10930 9370 10970
rect 9310 10910 9370 10930
rect 9690 11270 9750 11290
rect 9690 11230 9700 11270
rect 9740 11230 9750 11270
rect 9690 11170 9750 11230
rect 9690 11130 9700 11170
rect 9740 11130 9750 11170
rect 9690 11070 9750 11130
rect 9690 11030 9700 11070
rect 9740 11030 9750 11070
rect 9690 10970 9750 11030
rect 9690 10930 9700 10970
rect 9740 10930 9750 10970
rect 9690 10910 9750 10930
rect 9830 11270 9890 11290
rect 9830 11230 9840 11270
rect 9880 11230 9890 11270
rect 9830 11170 9890 11230
rect 9830 11130 9840 11170
rect 9880 11130 9890 11170
rect 9830 11070 9890 11130
rect 9830 11030 9840 11070
rect 9880 11030 9890 11070
rect 9830 10970 9890 11030
rect 9830 10930 9840 10970
rect 9880 10930 9890 10970
rect 9830 10910 9890 10930
rect 10210 11270 10270 11290
rect 10210 11230 10220 11270
rect 10260 11230 10270 11270
rect 10210 11170 10270 11230
rect 10210 11130 10220 11170
rect 10260 11130 10270 11170
rect 10210 11070 10270 11130
rect 10210 11030 10220 11070
rect 10260 11030 10270 11070
rect 10210 10970 10270 11030
rect 10210 10930 10220 10970
rect 10260 10930 10270 10970
rect 10210 10910 10270 10930
rect 10350 11270 10410 11290
rect 10350 11230 10360 11270
rect 10400 11230 10410 11270
rect 10350 11170 10410 11230
rect 10350 11130 10360 11170
rect 10400 11130 10410 11170
rect 10350 11070 10410 11130
rect 10350 11030 10360 11070
rect 10400 11030 10410 11070
rect 10350 10970 10410 11030
rect 10350 10930 10360 10970
rect 10400 10930 10410 10970
rect 10350 10910 10410 10930
rect 10730 11270 10790 11290
rect 10730 11230 10740 11270
rect 10780 11230 10790 11270
rect 10730 11170 10790 11230
rect 10730 11130 10740 11170
rect 10780 11130 10790 11170
rect 10730 11070 10790 11130
rect 10730 11030 10740 11070
rect 10780 11030 10790 11070
rect 10730 10970 10790 11030
rect 10730 10930 10740 10970
rect 10780 10930 10790 10970
rect 10730 10910 10790 10930
rect 10870 11270 10930 11290
rect 10870 11230 10880 11270
rect 10920 11230 10930 11270
rect 10870 11170 10930 11230
rect 10870 11130 10880 11170
rect 10920 11130 10930 11170
rect 10870 11070 10930 11130
rect 10870 11030 10880 11070
rect 10920 11030 10930 11070
rect 10870 10970 10930 11030
rect 10870 10930 10880 10970
rect 10920 10930 10930 10970
rect 10870 10910 10930 10930
rect 11250 11270 11310 11290
rect 11250 11230 11260 11270
rect 11300 11230 11310 11270
rect 11250 11170 11310 11230
rect 11250 11130 11260 11170
rect 11300 11130 11310 11170
rect 11250 11070 11310 11130
rect 11250 11030 11260 11070
rect 11300 11030 11310 11070
rect 11250 10970 11310 11030
rect 11250 10930 11260 10970
rect 11300 10930 11310 10970
rect 11250 10910 11310 10930
rect 9680 10840 9760 10860
rect 10200 10840 10280 10860
rect 10720 10840 10800 10860
rect 11240 10840 11320 10860
rect 11380 10840 11420 11270
rect 9200 10800 9700 10840
rect 9740 10800 10210 10840
rect 10370 10800 10740 10840
rect 10780 10800 11250 10840
rect 11320 10800 11420 10840
rect 9680 10780 9760 10800
rect 10200 10780 10280 10800
rect 10720 10780 10800 10800
rect 11240 10780 11320 10800
rect 9090 10520 9200 10540
rect -640 10440 -560 10460
rect -640 10400 -620 10440
rect -580 10400 -560 10440
rect -640 10380 -560 10400
rect -420 10440 -340 10460
rect -420 10400 -400 10440
rect -360 10400 -340 10440
rect -420 10380 -340 10400
rect -120 10440 -40 10460
rect -120 10400 -100 10440
rect -60 10400 -40 10440
rect -120 10380 -40 10400
rect 100 10440 180 10460
rect 100 10400 120 10440
rect 160 10400 180 10440
rect 100 10380 180 10400
rect 260 10440 340 10460
rect 260 10400 280 10440
rect 320 10400 340 10440
rect 260 10380 340 10400
rect 480 10440 560 10460
rect 480 10400 500 10440
rect 540 10400 560 10440
rect 480 10380 560 10400
rect 780 10440 860 10460
rect 780 10400 800 10440
rect 840 10400 860 10440
rect 780 10380 860 10400
rect 1000 10440 1080 10460
rect 1000 10400 1020 10440
rect 1060 10400 1080 10440
rect 1000 10380 1080 10400
rect 1300 10440 1380 10460
rect 1300 10400 1320 10440
rect 1360 10400 1380 10440
rect 1300 10380 1380 10400
rect 1740 10440 1820 10460
rect 1740 10400 1760 10440
rect 1800 10400 1820 10440
rect 1740 10380 1820 10400
rect 2070 10440 2150 10460
rect 2070 10400 2090 10440
rect 2130 10400 2150 10440
rect 2070 10380 2150 10400
rect 2500 10440 2580 10460
rect 2500 10400 2520 10440
rect 2560 10400 2580 10440
rect 2500 10380 2580 10400
rect 2890 10440 2970 10460
rect 2890 10400 2910 10440
rect 2950 10400 2970 10440
rect 2890 10380 2970 10400
rect 3280 10440 3360 10460
rect 3280 10400 3300 10440
rect 3340 10400 3360 10440
rect 9090 10450 9110 10520
rect 9180 10450 9200 10520
rect 9090 10430 9200 10450
rect 3280 10380 3360 10400
rect -620 10230 -580 10380
rect -400 10230 -360 10380
rect -230 10330 -150 10350
rect -230 10290 -210 10330
rect -170 10290 -150 10330
rect -230 10270 -150 10290
rect -710 10210 -570 10230
rect -710 10170 -700 10210
rect -660 10170 -620 10210
rect -580 10170 -570 10210
rect -710 10110 -570 10170
rect -710 10070 -700 10110
rect -660 10070 -620 10110
rect -580 10070 -570 10110
rect -710 10050 -570 10070
rect -520 10210 -460 10230
rect -520 10170 -510 10210
rect -470 10170 -460 10210
rect -520 10110 -460 10170
rect -520 10070 -510 10110
rect -470 10070 -460 10110
rect -520 10050 -460 10070
rect -410 10210 -350 10230
rect -410 10170 -400 10210
rect -360 10170 -350 10210
rect -410 10110 -350 10170
rect -410 10070 -400 10110
rect -360 10070 -350 10110
rect -410 10050 -350 10070
rect -760 9950 -680 9970
rect -760 9910 -740 9950
rect -700 9910 -680 9950
rect -760 9890 -680 9910
rect -520 9890 -480 10050
rect -430 9990 -350 10010
rect -430 9950 -410 9990
rect -370 9970 -350 9990
rect -190 9970 -150 10270
rect -100 10230 -60 10380
rect 120 10230 160 10380
rect 280 10230 320 10380
rect 500 10230 540 10380
rect 800 10230 840 10380
rect 1020 10230 1060 10380
rect 1320 10230 1360 10380
rect 1490 10330 1570 10350
rect 1490 10290 1510 10330
rect 1550 10290 1570 10330
rect 1490 10270 1570 10290
rect 1760 10230 1800 10380
rect 2090 10230 2130 10380
rect 2520 10230 2560 10380
rect 2910 10230 2950 10380
rect 3300 10230 3340 10380
rect 3570 10330 3650 10350
rect 3570 10290 3590 10330
rect 3630 10290 3650 10330
rect 3570 10270 3650 10290
rect 3590 10230 3630 10270
rect -110 10210 -50 10230
rect -110 10170 -100 10210
rect -60 10170 -50 10210
rect -110 10110 -50 10170
rect -110 10070 -100 10110
rect -60 10070 -50 10110
rect -110 10050 -50 10070
rect 0 10210 60 10230
rect 0 10170 10 10210
rect 50 10170 60 10210
rect 0 10110 60 10170
rect 0 10070 10 10110
rect 50 10070 60 10110
rect 0 10050 60 10070
rect 110 10210 330 10230
rect 110 10170 120 10210
rect 160 10170 200 10210
rect 240 10170 280 10210
rect 320 10170 330 10210
rect 110 10110 330 10170
rect 110 10070 120 10110
rect 160 10070 200 10110
rect 240 10070 280 10110
rect 320 10070 330 10110
rect 110 10050 330 10070
rect 380 10210 440 10230
rect 380 10170 390 10210
rect 430 10170 440 10210
rect 380 10110 440 10170
rect 380 10070 390 10110
rect 430 10070 440 10110
rect 380 10050 440 10070
rect 490 10210 550 10230
rect 490 10170 500 10210
rect 540 10170 550 10210
rect 490 10110 550 10170
rect 490 10070 500 10110
rect 540 10070 550 10110
rect 490 10050 550 10070
rect 790 10210 850 10230
rect 790 10170 800 10210
rect 840 10170 850 10210
rect 790 10110 850 10170
rect 790 10070 800 10110
rect 840 10070 850 10110
rect 790 10050 850 10070
rect 900 10210 960 10230
rect 900 10170 910 10210
rect 950 10170 960 10210
rect 900 10110 960 10170
rect 900 10070 910 10110
rect 950 10070 960 10110
rect 900 10050 960 10070
rect 1010 10210 1150 10230
rect 1010 10170 1020 10210
rect 1060 10170 1100 10210
rect 1140 10170 1150 10210
rect 1010 10110 1150 10170
rect 1010 10070 1020 10110
rect 1060 10070 1100 10110
rect 1140 10070 1150 10110
rect 1010 10050 1150 10070
rect 1230 10210 1370 10230
rect 1230 10170 1240 10210
rect 1280 10170 1320 10210
rect 1360 10170 1370 10210
rect 1230 10110 1370 10170
rect 1230 10070 1240 10110
rect 1280 10070 1320 10110
rect 1360 10070 1370 10110
rect 1230 10050 1370 10070
rect 1420 10210 1480 10230
rect 1420 10170 1430 10210
rect 1470 10170 1480 10210
rect 1420 10110 1480 10170
rect 1420 10070 1430 10110
rect 1470 10070 1480 10110
rect 1420 10050 1480 10070
rect 1530 10210 1590 10230
rect 1530 10170 1540 10210
rect 1580 10170 1590 10210
rect 1530 10110 1590 10170
rect 1530 10070 1540 10110
rect 1580 10070 1590 10110
rect 1530 10050 1590 10070
rect 1670 10210 1810 10230
rect 1670 10170 1680 10210
rect 1720 10170 1760 10210
rect 1800 10170 1810 10210
rect 1670 10110 1810 10170
rect 1670 10070 1680 10110
rect 1720 10070 1760 10110
rect 1800 10070 1810 10110
rect 1670 10050 1810 10070
rect 1860 10210 1920 10230
rect 1860 10170 1870 10210
rect 1910 10170 1920 10210
rect 1860 10110 1920 10170
rect 1860 10070 1870 10110
rect 1910 10070 1920 10110
rect 1860 10050 1920 10070
rect 2000 10210 2140 10230
rect 2000 10170 2010 10210
rect 2050 10170 2090 10210
rect 2130 10170 2140 10210
rect 2000 10110 2140 10170
rect 2000 10070 2010 10110
rect 2050 10070 2090 10110
rect 2130 10070 2140 10110
rect 2000 10050 2140 10070
rect 2190 10210 2250 10230
rect 2190 10170 2200 10210
rect 2240 10170 2250 10210
rect 2190 10110 2250 10170
rect 2190 10070 2200 10110
rect 2240 10070 2250 10110
rect 2190 10050 2250 10070
rect 2420 10210 2580 10230
rect 2420 10170 2430 10210
rect 2470 10170 2520 10210
rect 2560 10170 2580 10210
rect 2420 10110 2580 10170
rect 2420 10070 2430 10110
rect 2470 10070 2520 10110
rect 2560 10070 2580 10110
rect 2420 10050 2580 10070
rect 2630 10210 2710 10230
rect 2630 10170 2650 10210
rect 2690 10170 2710 10210
rect 2630 10110 2710 10170
rect 2630 10070 2650 10110
rect 2690 10070 2710 10110
rect 2630 10050 2710 10070
rect 2810 10210 2970 10230
rect 2810 10170 2820 10210
rect 2860 10170 2910 10210
rect 2950 10170 2970 10210
rect 2810 10110 2970 10170
rect 2810 10070 2820 10110
rect 2860 10070 2910 10110
rect 2950 10070 2970 10110
rect 2810 10050 2970 10070
rect 3020 10210 3100 10230
rect 3020 10170 3040 10210
rect 3080 10170 3100 10210
rect 3020 10110 3100 10170
rect 3020 10070 3040 10110
rect 3080 10070 3100 10110
rect 3020 10050 3100 10070
rect 3200 10210 3360 10230
rect 3200 10170 3210 10210
rect 3250 10170 3300 10210
rect 3340 10170 3360 10210
rect 3200 10110 3360 10170
rect 3200 10070 3210 10110
rect 3250 10070 3300 10110
rect 3340 10070 3360 10110
rect 3200 10050 3360 10070
rect 3410 10210 3490 10230
rect 3410 10170 3430 10210
rect 3470 10170 3490 10210
rect 3410 10110 3490 10170
rect 3410 10070 3430 10110
rect 3470 10070 3490 10110
rect 3410 10050 3490 10070
rect 3570 10210 3650 10230
rect 3570 10170 3590 10210
rect 3630 10170 3650 10210
rect 3570 10110 3650 10170
rect 3570 10070 3590 10110
rect 3630 10070 3650 10110
rect 3570 10050 3650 10070
rect 3700 10210 3780 10230
rect 3700 10170 3720 10210
rect 3760 10170 3780 10210
rect 3700 10110 3780 10170
rect 3700 10070 3720 10110
rect 3760 10070 3780 10110
rect 3700 10050 3780 10070
rect -370 9950 -150 9970
rect -430 9930 -150 9950
rect -520 9850 -360 9890
rect -400 9810 -360 9850
rect -710 9790 -570 9810
rect -710 9750 -700 9790
rect -660 9750 -620 9790
rect -580 9750 -570 9790
rect -710 9690 -570 9750
rect -710 9650 -700 9690
rect -660 9650 -620 9690
rect -580 9650 -570 9690
rect -710 9590 -570 9650
rect -710 9550 -700 9590
rect -660 9550 -620 9590
rect -580 9550 -570 9590
rect -710 9490 -570 9550
rect -710 9450 -700 9490
rect -660 9450 -620 9490
rect -580 9450 -570 9490
rect -710 9430 -570 9450
rect -520 9790 -460 9810
rect -520 9750 -510 9790
rect -470 9750 -460 9790
rect -520 9690 -460 9750
rect -520 9650 -510 9690
rect -470 9650 -460 9690
rect -520 9590 -460 9650
rect -520 9550 -510 9590
rect -470 9550 -460 9590
rect -520 9490 -460 9550
rect -520 9450 -510 9490
rect -470 9450 -460 9490
rect -520 9430 -460 9450
rect -410 9790 -350 9810
rect -410 9750 -400 9790
rect -360 9750 -350 9790
rect -410 9690 -350 9750
rect -410 9650 -400 9690
rect -360 9650 -350 9690
rect -410 9590 -350 9650
rect -410 9550 -400 9590
rect -360 9550 -350 9590
rect -410 9490 -350 9550
rect -410 9450 -400 9490
rect -360 9480 -350 9490
rect -310 9490 -230 9510
rect -310 9480 -290 9490
rect -360 9450 -290 9480
rect -250 9450 -230 9490
rect -410 9430 -230 9450
rect -190 9470 -150 9930
rect 10 9890 50 10050
rect -100 9850 50 9890
rect 90 9910 170 9930
rect 90 9870 110 9910
rect 150 9890 170 9910
rect 380 9890 420 10050
rect 470 9990 550 10010
rect 470 9950 490 9990
rect 530 9970 550 9990
rect 530 9950 750 9970
rect 470 9930 750 9950
rect 150 9870 540 9890
rect 90 9850 540 9870
rect -100 9810 -60 9850
rect 500 9810 540 9850
rect -110 9790 -50 9810
rect -110 9750 -100 9790
rect -60 9750 -50 9790
rect -110 9690 -50 9750
rect -110 9650 -100 9690
rect -60 9650 -50 9690
rect -110 9590 -50 9650
rect -110 9550 -100 9590
rect -60 9550 -50 9590
rect -110 9490 -50 9550
rect -110 9470 -100 9490
rect -190 9450 -100 9470
rect -60 9450 -50 9490
rect -190 9430 -50 9450
rect 0 9790 60 9810
rect 0 9750 10 9790
rect 50 9750 60 9790
rect 0 9690 60 9750
rect 0 9650 10 9690
rect 50 9650 60 9690
rect 0 9590 60 9650
rect 0 9550 10 9590
rect 50 9550 60 9590
rect 0 9490 60 9550
rect 0 9450 10 9490
rect 50 9450 60 9490
rect 0 9430 60 9450
rect 110 9790 330 9810
rect 110 9750 120 9790
rect 160 9750 200 9790
rect 240 9750 280 9790
rect 320 9750 330 9790
rect 110 9690 330 9750
rect 110 9650 120 9690
rect 160 9650 200 9690
rect 240 9650 280 9690
rect 320 9650 330 9690
rect 110 9590 330 9650
rect 110 9550 120 9590
rect 160 9550 200 9590
rect 240 9550 280 9590
rect 320 9550 330 9590
rect 110 9490 330 9550
rect 110 9450 120 9490
rect 160 9450 200 9490
rect 240 9450 280 9490
rect 320 9450 330 9490
rect 110 9430 330 9450
rect 380 9790 440 9810
rect 380 9750 390 9790
rect 430 9750 440 9790
rect 380 9690 440 9750
rect 380 9650 390 9690
rect 430 9650 440 9690
rect 380 9590 440 9650
rect 380 9550 390 9590
rect 430 9550 440 9590
rect 380 9490 440 9550
rect 380 9450 390 9490
rect 430 9450 440 9490
rect 380 9430 440 9450
rect 490 9790 550 9810
rect 490 9750 500 9790
rect 540 9750 550 9790
rect 490 9690 550 9750
rect 490 9650 500 9690
rect 540 9650 550 9690
rect 490 9590 550 9650
rect 490 9550 500 9590
rect 540 9550 550 9590
rect 490 9490 550 9550
rect 490 9450 500 9490
rect 540 9480 550 9490
rect 590 9490 670 9510
rect 590 9480 610 9490
rect 540 9450 610 9480
rect 650 9450 670 9490
rect 490 9430 670 9450
rect 710 9470 750 9930
rect 910 9890 950 10050
rect 1140 9980 1220 10000
rect 1140 9940 1160 9980
rect 1200 9940 1220 9980
rect 1140 9920 1220 9940
rect 1540 9960 1580 10050
rect 1880 9960 1920 10050
rect 2210 9960 2250 10050
rect 2360 9970 2440 9990
rect 1540 9940 1650 9960
rect 1540 9920 1590 9940
rect 800 9850 950 9890
rect 1430 9900 1590 9920
rect 1630 9900 1650 9940
rect 1430 9880 1650 9900
rect 1880 9940 1980 9960
rect 1880 9900 1920 9940
rect 1960 9900 1980 9940
rect 1880 9880 1980 9900
rect 2210 9940 2310 9960
rect 2210 9900 2250 9940
rect 2290 9900 2310 9940
rect 2360 9930 2380 9970
rect 2420 9930 2440 9970
rect 2360 9910 2440 9930
rect 2670 9940 2710 10050
rect 3060 9970 3100 10050
rect 3320 9990 3400 10010
rect 3320 9970 3340 9990
rect 2930 9940 3010 9960
rect 2210 9880 2310 9900
rect 2670 9900 2950 9940
rect 2990 9900 3010 9940
rect 800 9810 840 9850
rect 1430 9810 1470 9880
rect 1880 9810 1920 9880
rect 2210 9810 2250 9880
rect 2670 9810 2710 9900
rect 2930 9880 3010 9900
rect 3060 9950 3340 9970
rect 3380 9950 3400 9990
rect 3060 9930 3400 9950
rect 3450 9930 3490 10050
rect 3060 9810 3100 9930
rect 3450 9910 3530 9930
rect 3450 9870 3470 9910
rect 3510 9870 3530 9910
rect 3450 9850 3530 9870
rect 3450 9810 3490 9850
rect 3590 9810 3630 10050
rect 3720 10010 3760 10050
rect 3720 9990 4190 10010
rect 3720 9970 4130 9990
rect 3720 9810 3760 9970
rect 4110 9950 4130 9970
rect 4170 9950 4190 9990
rect 4110 9930 4190 9950
rect 3800 9910 3880 9930
rect 3800 9870 3820 9910
rect 3860 9870 3880 9910
rect 3800 9850 3880 9870
rect 4110 9810 4150 9930
rect 5650 9880 5730 9900
rect 5650 9840 5670 9880
rect 5710 9840 5730 9880
rect 5650 9820 5730 9840
rect 8490 9880 8570 9900
rect 8490 9840 8510 9880
rect 8550 9840 8570 9880
rect 8490 9820 8570 9840
rect 790 9790 850 9810
rect 790 9750 800 9790
rect 840 9750 850 9790
rect 790 9690 850 9750
rect 790 9650 800 9690
rect 840 9650 850 9690
rect 790 9590 850 9650
rect 790 9550 800 9590
rect 840 9550 850 9590
rect 790 9490 850 9550
rect 790 9470 800 9490
rect 710 9450 800 9470
rect 840 9450 850 9490
rect 710 9430 850 9450
rect 900 9790 960 9810
rect 900 9750 910 9790
rect 950 9750 960 9790
rect 900 9690 960 9750
rect 900 9650 910 9690
rect 950 9650 960 9690
rect 900 9590 960 9650
rect 900 9550 910 9590
rect 950 9550 960 9590
rect 900 9490 960 9550
rect 900 9450 910 9490
rect 950 9450 960 9490
rect 900 9430 960 9450
rect 1010 9790 1150 9810
rect 1010 9750 1020 9790
rect 1060 9750 1100 9790
rect 1140 9750 1150 9790
rect 1010 9690 1150 9750
rect 1010 9650 1020 9690
rect 1060 9650 1100 9690
rect 1140 9650 1150 9690
rect 1010 9590 1150 9650
rect 1010 9550 1020 9590
rect 1060 9550 1100 9590
rect 1140 9550 1150 9590
rect 1010 9490 1150 9550
rect 1010 9450 1020 9490
rect 1060 9450 1100 9490
rect 1140 9450 1150 9490
rect 1010 9430 1150 9450
rect 1230 9790 1370 9810
rect 1230 9750 1240 9790
rect 1280 9750 1320 9790
rect 1360 9750 1370 9790
rect 1230 9690 1370 9750
rect 1230 9650 1240 9690
rect 1280 9650 1320 9690
rect 1360 9650 1370 9690
rect 1230 9590 1370 9650
rect 1230 9550 1240 9590
rect 1280 9550 1320 9590
rect 1360 9550 1370 9590
rect 1230 9490 1370 9550
rect 1230 9450 1240 9490
rect 1280 9450 1320 9490
rect 1360 9450 1370 9490
rect 1230 9430 1370 9450
rect 1420 9790 1480 9810
rect 1420 9750 1430 9790
rect 1470 9750 1480 9790
rect 1420 9690 1480 9750
rect 1420 9650 1430 9690
rect 1470 9650 1480 9690
rect 1420 9590 1480 9650
rect 1420 9550 1430 9590
rect 1470 9550 1480 9590
rect 1420 9490 1480 9550
rect 1420 9450 1430 9490
rect 1470 9450 1480 9490
rect 1420 9430 1480 9450
rect 1530 9790 1590 9810
rect 1530 9750 1540 9790
rect 1580 9750 1590 9790
rect 1530 9690 1590 9750
rect 1530 9650 1540 9690
rect 1580 9650 1590 9690
rect 1530 9590 1590 9650
rect 1530 9550 1540 9590
rect 1580 9550 1590 9590
rect 1530 9490 1590 9550
rect 1530 9450 1540 9490
rect 1580 9450 1590 9490
rect 1530 9430 1590 9450
rect 1670 9790 1810 9810
rect 1670 9750 1680 9790
rect 1720 9750 1760 9790
rect 1800 9750 1810 9790
rect 1670 9690 1810 9750
rect 1670 9650 1680 9690
rect 1720 9650 1760 9690
rect 1800 9650 1810 9690
rect 1670 9590 1810 9650
rect 1670 9550 1680 9590
rect 1720 9550 1760 9590
rect 1800 9550 1810 9590
rect 1670 9490 1810 9550
rect 1670 9450 1680 9490
rect 1720 9450 1760 9490
rect 1800 9450 1810 9490
rect 1670 9430 1810 9450
rect 1860 9790 1920 9810
rect 1860 9750 1870 9790
rect 1910 9750 1920 9790
rect 1860 9690 1920 9750
rect 1860 9650 1870 9690
rect 1910 9650 1920 9690
rect 1860 9590 1920 9650
rect 1860 9550 1870 9590
rect 1910 9550 1920 9590
rect 1860 9490 1920 9550
rect 1860 9450 1870 9490
rect 1910 9450 1920 9490
rect 1860 9430 1920 9450
rect 2000 9790 2140 9810
rect 2000 9750 2010 9790
rect 2050 9750 2090 9790
rect 2130 9750 2140 9790
rect 2000 9690 2140 9750
rect 2000 9650 2010 9690
rect 2050 9650 2090 9690
rect 2130 9650 2140 9690
rect 2000 9590 2140 9650
rect 2000 9550 2010 9590
rect 2050 9550 2090 9590
rect 2130 9550 2140 9590
rect 2000 9490 2140 9550
rect 2000 9450 2010 9490
rect 2050 9450 2090 9490
rect 2130 9450 2140 9490
rect 2000 9430 2140 9450
rect 2190 9790 2250 9810
rect 2190 9750 2200 9790
rect 2240 9750 2250 9790
rect 2190 9690 2250 9750
rect 2190 9650 2200 9690
rect 2240 9650 2250 9690
rect 2190 9590 2250 9650
rect 2190 9550 2200 9590
rect 2240 9550 2250 9590
rect 2190 9490 2250 9550
rect 2190 9450 2200 9490
rect 2240 9450 2250 9490
rect 2190 9430 2250 9450
rect 2400 9790 2580 9810
rect 2400 9750 2420 9790
rect 2460 9750 2520 9790
rect 2560 9750 2580 9790
rect 2400 9690 2580 9750
rect 2400 9650 2420 9690
rect 2460 9650 2520 9690
rect 2560 9650 2580 9690
rect 2400 9590 2580 9650
rect 2400 9550 2420 9590
rect 2460 9550 2520 9590
rect 2560 9550 2580 9590
rect 2400 9490 2580 9550
rect 2400 9450 2420 9490
rect 2460 9450 2520 9490
rect 2560 9450 2580 9490
rect 2400 9430 2580 9450
rect 2630 9790 2710 9810
rect 2630 9750 2650 9790
rect 2690 9750 2710 9790
rect 2630 9690 2710 9750
rect 2630 9650 2650 9690
rect 2690 9650 2710 9690
rect 2630 9590 2710 9650
rect 2630 9550 2650 9590
rect 2690 9550 2710 9590
rect 2630 9490 2710 9550
rect 2630 9450 2650 9490
rect 2690 9450 2710 9490
rect 2630 9430 2710 9450
rect 2790 9790 2970 9810
rect 2790 9750 2810 9790
rect 2850 9750 2910 9790
rect 2950 9750 2970 9790
rect 2790 9690 2970 9750
rect 2790 9650 2810 9690
rect 2850 9650 2910 9690
rect 2950 9650 2970 9690
rect 2790 9590 2970 9650
rect 2790 9550 2810 9590
rect 2850 9550 2910 9590
rect 2950 9550 2970 9590
rect 2790 9490 2970 9550
rect 2790 9450 2810 9490
rect 2850 9450 2910 9490
rect 2950 9450 2970 9490
rect 2790 9430 2970 9450
rect 3020 9790 3100 9810
rect 3020 9750 3040 9790
rect 3080 9750 3100 9790
rect 3020 9690 3100 9750
rect 3020 9650 3040 9690
rect 3080 9650 3100 9690
rect 3020 9590 3100 9650
rect 3020 9550 3040 9590
rect 3080 9550 3100 9590
rect 3020 9490 3100 9550
rect 3020 9450 3040 9490
rect 3080 9450 3100 9490
rect 3020 9430 3100 9450
rect 3180 9790 3360 9810
rect 3180 9750 3200 9790
rect 3240 9750 3300 9790
rect 3340 9750 3360 9790
rect 3180 9690 3360 9750
rect 3180 9650 3200 9690
rect 3240 9650 3300 9690
rect 3340 9650 3360 9690
rect 3180 9590 3360 9650
rect 3180 9550 3200 9590
rect 3240 9550 3300 9590
rect 3340 9550 3360 9590
rect 3180 9490 3360 9550
rect 3180 9450 3200 9490
rect 3240 9450 3300 9490
rect 3340 9450 3360 9490
rect 3180 9430 3360 9450
rect 3410 9790 3490 9810
rect 3410 9750 3430 9790
rect 3470 9750 3490 9790
rect 3410 9690 3490 9750
rect 3410 9650 3430 9690
rect 3470 9650 3490 9690
rect 3410 9590 3490 9650
rect 3410 9550 3430 9590
rect 3470 9550 3490 9590
rect 3410 9490 3490 9550
rect 3410 9450 3430 9490
rect 3470 9450 3490 9490
rect 3410 9430 3490 9450
rect 3570 9790 3650 9810
rect 3570 9750 3590 9790
rect 3630 9750 3650 9790
rect 3570 9690 3650 9750
rect 3570 9650 3590 9690
rect 3630 9650 3650 9690
rect 3570 9590 3650 9650
rect 3570 9550 3590 9590
rect 3630 9550 3650 9590
rect 3570 9490 3650 9550
rect 3570 9450 3590 9490
rect 3630 9450 3650 9490
rect 3570 9430 3650 9450
rect 3700 9790 3780 9810
rect 3700 9750 3720 9790
rect 3760 9750 3780 9790
rect 3700 9690 3780 9750
rect 3700 9650 3720 9690
rect 3760 9650 3780 9690
rect 3700 9590 3780 9650
rect 3700 9550 3720 9590
rect 3760 9550 3780 9590
rect 3700 9490 3780 9550
rect 3700 9450 3720 9490
rect 3760 9450 3780 9490
rect 3700 9430 3780 9450
rect 3860 9790 4040 9810
rect 3860 9750 3880 9790
rect 3920 9750 3980 9790
rect 4020 9750 4040 9790
rect 3860 9690 4040 9750
rect 3860 9650 3880 9690
rect 3920 9650 3980 9690
rect 4020 9650 4040 9690
rect 3860 9590 4040 9650
rect 3860 9550 3880 9590
rect 3920 9550 3980 9590
rect 4020 9550 4040 9590
rect 3860 9490 4040 9550
rect 3860 9450 3880 9490
rect 3920 9450 3980 9490
rect 4020 9450 4040 9490
rect 3860 9430 4040 9450
rect 4090 9790 4170 9810
rect 4090 9750 4110 9790
rect 4150 9750 4170 9790
rect 4090 9690 4170 9750
rect 4090 9650 4110 9690
rect 4150 9650 4170 9690
rect 4090 9590 4170 9650
rect 4090 9550 4110 9590
rect 4150 9550 4170 9590
rect 4090 9490 4170 9550
rect 4090 9450 4110 9490
rect 4150 9450 4170 9490
rect 4090 9430 4170 9450
rect 5550 9760 5730 9780
rect 5550 9720 5570 9760
rect 5610 9720 5670 9760
rect 5710 9720 5730 9760
rect 5550 9660 5730 9720
rect 5550 9620 5570 9660
rect 5610 9620 5670 9660
rect 5710 9620 5730 9660
rect 5550 9560 5730 9620
rect 5550 9520 5570 9560
rect 5610 9520 5670 9560
rect 5710 9520 5730 9560
rect 5550 9460 5730 9520
rect -620 9280 -580 9430
rect 120 9280 160 9430
rect 280 9280 320 9430
rect 1020 9280 1060 9430
rect 1280 9280 1320 9430
rect 1360 9370 1440 9390
rect 1360 9330 1380 9370
rect 1420 9330 1440 9370
rect 1360 9320 1440 9330
rect 1540 9280 1580 9430
rect 1760 9280 1800 9430
rect 2090 9280 2130 9430
rect 2520 9280 2560 9430
rect 2910 9280 2950 9430
rect 3300 9280 3340 9430
rect 3980 9280 4020 9430
rect 5550 9420 5570 9460
rect 5610 9420 5670 9460
rect 5710 9420 5730 9460
rect 5550 9400 5730 9420
rect 5870 9760 5950 9780
rect 5870 9720 5890 9760
rect 5930 9720 5950 9760
rect 5870 9660 5950 9720
rect 5870 9620 5890 9660
rect 5930 9620 5950 9660
rect 5870 9560 5950 9620
rect 5870 9520 5890 9560
rect 5930 9520 5950 9560
rect 5870 9460 5950 9520
rect 5870 9420 5890 9460
rect 5930 9420 5950 9460
rect 5870 9400 5950 9420
rect 6090 9760 6170 9780
rect 6090 9720 6110 9760
rect 6150 9720 6170 9760
rect 6090 9660 6170 9720
rect 6090 9620 6110 9660
rect 6150 9620 6170 9660
rect 6090 9560 6170 9620
rect 6090 9520 6110 9560
rect 6150 9520 6170 9560
rect 6090 9460 6170 9520
rect 6090 9420 6110 9460
rect 6150 9420 6170 9460
rect 6090 9400 6170 9420
rect 6310 9760 6390 9780
rect 6310 9720 6330 9760
rect 6370 9720 6390 9760
rect 6310 9660 6390 9720
rect 6310 9620 6330 9660
rect 6370 9620 6390 9660
rect 6310 9560 6390 9620
rect 6310 9520 6330 9560
rect 6370 9520 6390 9560
rect 6310 9460 6390 9520
rect 6310 9420 6330 9460
rect 6370 9420 6390 9460
rect 6310 9400 6390 9420
rect 6530 9760 6610 9780
rect 6530 9720 6550 9760
rect 6590 9720 6610 9760
rect 6530 9660 6610 9720
rect 6530 9620 6550 9660
rect 6590 9620 6610 9660
rect 6530 9560 6610 9620
rect 6530 9520 6550 9560
rect 6590 9520 6610 9560
rect 6530 9460 6610 9520
rect 6530 9420 6550 9460
rect 6590 9420 6610 9460
rect 6530 9400 6610 9420
rect 6750 9760 6830 9780
rect 6750 9720 6770 9760
rect 6810 9720 6830 9760
rect 6750 9660 6830 9720
rect 6750 9620 6770 9660
rect 6810 9620 6830 9660
rect 6750 9560 6830 9620
rect 6750 9520 6770 9560
rect 6810 9520 6830 9560
rect 6750 9460 6830 9520
rect 6750 9420 6770 9460
rect 6810 9420 6830 9460
rect 6750 9400 6830 9420
rect 6970 9760 7250 9780
rect 6970 9720 6990 9760
rect 7030 9720 7090 9760
rect 7130 9720 7190 9760
rect 7230 9720 7250 9760
rect 6970 9660 7250 9720
rect 6970 9620 6990 9660
rect 7030 9620 7090 9660
rect 7130 9620 7190 9660
rect 7230 9620 7250 9660
rect 6970 9560 7250 9620
rect 6970 9520 6990 9560
rect 7030 9520 7090 9560
rect 7130 9520 7190 9560
rect 7230 9520 7250 9560
rect 6970 9460 7250 9520
rect 6970 9420 6990 9460
rect 7030 9420 7090 9460
rect 7130 9420 7190 9460
rect 7230 9420 7250 9460
rect 6970 9400 7250 9420
rect 7390 9760 7470 9780
rect 7390 9720 7410 9760
rect 7450 9720 7470 9760
rect 7390 9660 7470 9720
rect 7390 9620 7410 9660
rect 7450 9620 7470 9660
rect 7390 9560 7470 9620
rect 7390 9520 7410 9560
rect 7450 9520 7470 9560
rect 7390 9460 7470 9520
rect 7390 9420 7410 9460
rect 7450 9420 7470 9460
rect 7390 9400 7470 9420
rect 7610 9760 7690 9780
rect 7610 9720 7630 9760
rect 7670 9720 7690 9760
rect 7610 9660 7690 9720
rect 7610 9620 7630 9660
rect 7670 9620 7690 9660
rect 7610 9560 7690 9620
rect 7610 9520 7630 9560
rect 7670 9520 7690 9560
rect 7610 9460 7690 9520
rect 7610 9420 7630 9460
rect 7670 9420 7690 9460
rect 7610 9400 7690 9420
rect 7830 9760 7910 9780
rect 7830 9720 7850 9760
rect 7890 9720 7910 9760
rect 7830 9660 7910 9720
rect 7830 9620 7850 9660
rect 7890 9620 7910 9660
rect 7830 9560 7910 9620
rect 7830 9520 7850 9560
rect 7890 9520 7910 9560
rect 7830 9460 7910 9520
rect 7830 9420 7850 9460
rect 7890 9420 7910 9460
rect 7830 9400 7910 9420
rect 8050 9760 8130 9780
rect 8050 9720 8070 9760
rect 8110 9720 8130 9760
rect 8050 9660 8130 9720
rect 8050 9620 8070 9660
rect 8110 9620 8130 9660
rect 8050 9560 8130 9620
rect 8050 9520 8070 9560
rect 8110 9520 8130 9560
rect 8050 9460 8130 9520
rect 8050 9420 8070 9460
rect 8110 9420 8130 9460
rect 8050 9400 8130 9420
rect 8270 9760 8350 9780
rect 8270 9720 8290 9760
rect 8330 9720 8350 9760
rect 8270 9660 8350 9720
rect 8270 9620 8290 9660
rect 8330 9620 8350 9660
rect 8270 9560 8350 9620
rect 8270 9520 8290 9560
rect 8330 9520 8350 9560
rect 8270 9460 8350 9520
rect 8270 9420 8290 9460
rect 8330 9420 8350 9460
rect 8270 9400 8350 9420
rect 8490 9760 8670 9780
rect 8490 9720 8510 9760
rect 8550 9720 8610 9760
rect 8650 9720 8670 9760
rect 8490 9660 8670 9720
rect 8490 9620 8510 9660
rect 8550 9620 8610 9660
rect 8650 9620 8670 9660
rect 8490 9560 8670 9620
rect 8490 9520 8510 9560
rect 8550 9520 8610 9560
rect 8650 9520 8670 9560
rect 8490 9460 8670 9520
rect 8490 9420 8510 9460
rect 8550 9420 8610 9460
rect 8650 9420 8670 9460
rect 8490 9400 8670 9420
rect 6310 9340 6390 9360
rect 6310 9300 6330 9340
rect 6370 9300 6390 9340
rect 6310 9280 6390 9300
rect 7070 9340 7150 9400
rect 7070 9300 7090 9340
rect 7130 9300 7150 9340
rect 8850 9340 8960 9360
rect 7070 9280 7150 9300
rect 7480 9310 7560 9330
rect -640 9260 -560 9280
rect -640 9220 -620 9260
rect -580 9220 -560 9260
rect -640 9200 -560 9220
rect 100 9260 180 9280
rect 100 9220 120 9260
rect 160 9220 180 9260
rect 100 9200 180 9220
rect 260 9260 340 9280
rect 260 9220 280 9260
rect 320 9220 340 9260
rect 260 9200 340 9220
rect 1000 9260 1080 9280
rect 1000 9220 1020 9260
rect 1060 9220 1080 9260
rect 1000 9200 1080 9220
rect 1250 9260 1330 9280
rect 1250 9220 1270 9260
rect 1310 9220 1330 9260
rect 1250 9200 1330 9220
rect 1440 9260 1600 9280
rect 1440 9220 1460 9260
rect 1500 9220 1540 9260
rect 1580 9220 1600 9260
rect 1440 9200 1600 9220
rect 1730 9260 1810 9280
rect 1730 9220 1750 9260
rect 1790 9220 1810 9260
rect 1730 9200 1810 9220
rect 2060 9260 2140 9280
rect 2060 9220 2080 9260
rect 2120 9220 2140 9260
rect 2060 9200 2140 9220
rect 2500 9260 2580 9280
rect 2500 9220 2520 9260
rect 2560 9220 2580 9260
rect 2500 9200 2580 9220
rect 2890 9260 2970 9280
rect 2890 9220 2910 9260
rect 2950 9220 2970 9260
rect 2890 9200 2970 9220
rect 3280 9260 3360 9280
rect 3280 9220 3300 9260
rect 3340 9220 3360 9260
rect 3280 9200 3360 9220
rect 3960 9260 4040 9280
rect 3960 9220 3980 9260
rect 4020 9220 4040 9260
rect 7480 9270 7500 9310
rect 7540 9270 7560 9310
rect 7480 9250 7560 9270
rect 8180 9310 8260 9330
rect 8180 9270 8200 9310
rect 8240 9270 8260 9310
rect 8180 9250 8260 9270
rect 8850 9270 8870 9340
rect 8940 9270 8960 9340
rect 8850 9250 8960 9270
rect 3960 9200 4040 9220
rect -620 9050 -580 9200
rect -190 9150 -110 9170
rect -190 9110 -170 9150
rect -130 9110 -110 9150
rect -190 9090 -110 9110
rect -190 9050 -150 9090
rect 120 9050 160 9200
rect 280 9050 320 9200
rect 1020 9050 1060 9200
rect 1440 9050 1480 9200
rect 1750 9050 1790 9200
rect 2080 9050 2120 9200
rect 2520 9050 2560 9200
rect 2930 9150 3010 9160
rect 2930 9110 2950 9150
rect 2990 9110 3010 9150
rect 2930 9090 3010 9110
rect 3300 9050 3340 9200
rect 3570 9150 3650 9170
rect 3570 9110 3590 9150
rect 3630 9110 3650 9150
rect 3570 9090 3650 9110
rect 3590 9050 3630 9090
rect -710 9030 -570 9050
rect -710 8990 -700 9030
rect -660 8990 -620 9030
rect -580 8990 -570 9030
rect -710 8930 -570 8990
rect -710 8890 -700 8930
rect -660 8890 -620 8930
rect -580 8890 -570 8930
rect -710 8830 -570 8890
rect -710 8790 -700 8830
rect -660 8790 -620 8830
rect -580 8790 -570 8830
rect -710 8730 -570 8790
rect -710 8690 -700 8730
rect -660 8690 -620 8730
rect -580 8690 -570 8730
rect -710 8670 -570 8690
rect -520 9030 -460 9050
rect -520 8990 -510 9030
rect -470 8990 -460 9030
rect -520 8930 -460 8990
rect -520 8890 -510 8930
rect -470 8890 -460 8930
rect -520 8830 -460 8890
rect -520 8790 -510 8830
rect -470 8790 -460 8830
rect -520 8730 -460 8790
rect -520 8690 -510 8730
rect -470 8690 -460 8730
rect -520 8670 -460 8690
rect -410 9030 -230 9050
rect -410 8990 -400 9030
rect -360 9000 -290 9030
rect -360 8990 -350 9000
rect -410 8930 -350 8990
rect -310 8990 -290 9000
rect -250 8990 -230 9030
rect -310 8970 -230 8990
rect -190 9030 -50 9050
rect -190 9010 -100 9030
rect -410 8890 -400 8930
rect -360 8890 -350 8930
rect -410 8830 -350 8890
rect -410 8790 -400 8830
rect -360 8790 -350 8830
rect -410 8730 -350 8790
rect -410 8690 -400 8730
rect -360 8690 -350 8730
rect -410 8670 -350 8690
rect -400 8630 -360 8670
rect -520 8590 -360 8630
rect -760 8570 -680 8590
rect -760 8530 -740 8570
rect -700 8530 -680 8570
rect -760 8510 -680 8530
rect -520 8430 -480 8590
rect -190 8550 -150 9010
rect -110 8990 -100 9010
rect -60 8990 -50 9030
rect -110 8930 -50 8990
rect -110 8890 -100 8930
rect -60 8890 -50 8930
rect -110 8830 -50 8890
rect -110 8790 -100 8830
rect -60 8790 -50 8830
rect -110 8730 -50 8790
rect -110 8690 -100 8730
rect -60 8690 -50 8730
rect -110 8670 -50 8690
rect 0 9030 60 9050
rect 0 8990 10 9030
rect 50 8990 60 9030
rect 0 8930 60 8990
rect 0 8890 10 8930
rect 50 8890 60 8930
rect 0 8830 60 8890
rect 0 8790 10 8830
rect 50 8790 60 8830
rect 0 8730 60 8790
rect 0 8690 10 8730
rect 50 8690 60 8730
rect 0 8670 60 8690
rect 110 9030 330 9050
rect 110 8990 120 9030
rect 160 8990 200 9030
rect 240 8990 280 9030
rect 320 8990 330 9030
rect 110 8930 330 8990
rect 110 8890 120 8930
rect 160 8890 200 8930
rect 240 8890 280 8930
rect 320 8890 330 8930
rect 110 8830 330 8890
rect 110 8790 120 8830
rect 160 8790 200 8830
rect 240 8790 280 8830
rect 320 8790 330 8830
rect 110 8730 330 8790
rect 110 8690 120 8730
rect 160 8690 200 8730
rect 240 8690 280 8730
rect 320 8690 330 8730
rect 110 8670 330 8690
rect 380 9030 440 9050
rect 380 8990 390 9030
rect 430 8990 440 9030
rect 380 8930 440 8990
rect 380 8890 390 8930
rect 430 8890 440 8930
rect 380 8830 440 8890
rect 380 8790 390 8830
rect 430 8790 440 8830
rect 380 8730 440 8790
rect 380 8690 390 8730
rect 430 8690 440 8730
rect 380 8670 440 8690
rect 490 9030 670 9050
rect 490 8990 500 9030
rect 540 9000 610 9030
rect 540 8990 550 9000
rect 490 8930 550 8990
rect 590 8990 610 9000
rect 650 8990 670 9030
rect 590 8970 670 8990
rect 710 9030 850 9050
rect 710 9010 800 9030
rect 490 8890 500 8930
rect 540 8890 550 8930
rect 490 8830 550 8890
rect 490 8790 500 8830
rect 540 8790 550 8830
rect 490 8730 550 8790
rect 490 8690 500 8730
rect 540 8690 550 8730
rect 490 8670 550 8690
rect -100 8630 -60 8670
rect 500 8630 540 8670
rect -100 8590 50 8630
rect -430 8530 -150 8550
rect -430 8490 -410 8530
rect -370 8510 -150 8530
rect -370 8490 -350 8510
rect -430 8470 -350 8490
rect 10 8430 50 8590
rect 90 8610 540 8630
rect 90 8570 110 8610
rect 150 8590 540 8610
rect 150 8570 170 8590
rect 90 8550 170 8570
rect 380 8430 420 8590
rect 710 8550 750 9010
rect 790 8990 800 9010
rect 840 8990 850 9030
rect 790 8930 850 8990
rect 790 8890 800 8930
rect 840 8890 850 8930
rect 790 8830 850 8890
rect 790 8790 800 8830
rect 840 8790 850 8830
rect 790 8730 850 8790
rect 790 8690 800 8730
rect 840 8690 850 8730
rect 790 8670 850 8690
rect 900 9030 960 9050
rect 900 8990 910 9030
rect 950 8990 960 9030
rect 900 8930 960 8990
rect 900 8890 910 8930
rect 950 8890 960 8930
rect 900 8830 960 8890
rect 900 8790 910 8830
rect 950 8790 960 8830
rect 900 8730 960 8790
rect 900 8690 910 8730
rect 950 8690 960 8730
rect 900 8670 960 8690
rect 1010 9030 1150 9050
rect 1010 8990 1020 9030
rect 1060 8990 1100 9030
rect 1140 8990 1150 9030
rect 1010 8930 1150 8990
rect 1010 8890 1020 8930
rect 1060 8890 1100 8930
rect 1140 8890 1150 8930
rect 1010 8830 1150 8890
rect 1010 8790 1020 8830
rect 1060 8790 1100 8830
rect 1140 8790 1150 8830
rect 1010 8730 1150 8790
rect 1010 8690 1020 8730
rect 1060 8690 1100 8730
rect 1140 8690 1150 8730
rect 1010 8670 1150 8690
rect 1300 9030 1360 9050
rect 1300 8990 1310 9030
rect 1350 8990 1360 9030
rect 1300 8930 1360 8990
rect 1300 8890 1310 8930
rect 1350 8890 1360 8930
rect 1300 8830 1360 8890
rect 1300 8790 1310 8830
rect 1350 8790 1360 8830
rect 1300 8730 1360 8790
rect 1300 8690 1310 8730
rect 1350 8690 1360 8730
rect 1300 8670 1360 8690
rect 1410 9030 1550 9050
rect 1410 8990 1420 9030
rect 1460 8990 1500 9030
rect 1540 8990 1550 9030
rect 1410 8930 1550 8990
rect 1410 8890 1420 8930
rect 1460 8890 1500 8930
rect 1540 8890 1550 8930
rect 1410 8830 1550 8890
rect 1410 8790 1420 8830
rect 1460 8790 1500 8830
rect 1540 8790 1550 8830
rect 1410 8730 1550 8790
rect 1410 8690 1420 8730
rect 1460 8690 1500 8730
rect 1540 8690 1550 8730
rect 1410 8670 1550 8690
rect 1630 9030 1690 9050
rect 1630 8990 1640 9030
rect 1680 8990 1690 9030
rect 1630 8930 1690 8990
rect 1630 8890 1640 8930
rect 1680 8890 1690 8930
rect 1630 8830 1690 8890
rect 1630 8790 1640 8830
rect 1680 8790 1690 8830
rect 1630 8730 1690 8790
rect 1630 8690 1640 8730
rect 1680 8690 1690 8730
rect 1630 8670 1690 8690
rect 1740 9030 1880 9050
rect 1740 8990 1750 9030
rect 1790 8990 1830 9030
rect 1870 8990 1880 9030
rect 1740 8930 1880 8990
rect 1740 8890 1750 8930
rect 1790 8890 1830 8930
rect 1870 8890 1880 8930
rect 1740 8830 1880 8890
rect 1740 8790 1750 8830
rect 1790 8790 1830 8830
rect 1870 8790 1880 8830
rect 1740 8730 1880 8790
rect 1740 8690 1750 8730
rect 1790 8690 1830 8730
rect 1870 8690 1880 8730
rect 1740 8670 1880 8690
rect 1960 9030 2020 9050
rect 1960 8990 1970 9030
rect 2010 8990 2020 9030
rect 1960 8930 2020 8990
rect 1960 8890 1970 8930
rect 2010 8890 2020 8930
rect 1960 8830 2020 8890
rect 1960 8790 1970 8830
rect 2010 8790 2020 8830
rect 1960 8730 2020 8790
rect 1960 8690 1970 8730
rect 2010 8690 2020 8730
rect 1960 8670 2020 8690
rect 2070 9030 2210 9050
rect 2070 8990 2080 9030
rect 2120 8990 2160 9030
rect 2200 8990 2210 9030
rect 2070 8930 2210 8990
rect 2070 8890 2080 8930
rect 2120 8890 2160 8930
rect 2200 8890 2210 8930
rect 2070 8830 2210 8890
rect 2070 8790 2080 8830
rect 2120 8790 2160 8830
rect 2200 8790 2210 8830
rect 2070 8730 2210 8790
rect 2070 8690 2080 8730
rect 2120 8690 2160 8730
rect 2200 8690 2210 8730
rect 2070 8670 2210 8690
rect 2400 9030 2580 9050
rect 2400 8990 2420 9030
rect 2460 8990 2520 9030
rect 2560 8990 2580 9030
rect 2400 8930 2580 8990
rect 2400 8890 2420 8930
rect 2460 8890 2520 8930
rect 2560 8890 2580 8930
rect 2400 8830 2580 8890
rect 2400 8790 2420 8830
rect 2460 8790 2520 8830
rect 2560 8790 2580 8830
rect 2400 8730 2580 8790
rect 2400 8690 2420 8730
rect 2460 8690 2520 8730
rect 2560 8690 2580 8730
rect 2400 8670 2580 8690
rect 2630 9030 2710 9050
rect 2630 8990 2650 9030
rect 2690 8990 2710 9030
rect 2630 8930 2710 8990
rect 2630 8890 2650 8930
rect 2690 8890 2710 8930
rect 2630 8830 2710 8890
rect 2630 8790 2650 8830
rect 2690 8790 2710 8830
rect 2630 8730 2710 8790
rect 2630 8690 2650 8730
rect 2690 8690 2710 8730
rect 2630 8670 2710 8690
rect 2890 9030 2970 9050
rect 2890 8990 2910 9030
rect 2950 8990 2970 9030
rect 2890 8930 2970 8990
rect 2890 8890 2910 8930
rect 2950 8890 2970 8930
rect 2890 8830 2970 8890
rect 2890 8790 2910 8830
rect 2950 8790 2970 8830
rect 2890 8730 2970 8790
rect 2890 8690 2910 8730
rect 2950 8690 2970 8730
rect 2890 8670 2970 8690
rect 3020 9030 3100 9050
rect 3020 8990 3040 9030
rect 3080 8990 3100 9030
rect 3020 8930 3100 8990
rect 3020 8890 3040 8930
rect 3080 8890 3100 8930
rect 3020 8830 3100 8890
rect 3020 8790 3040 8830
rect 3080 8790 3100 8830
rect 3020 8730 3100 8790
rect 3020 8690 3040 8730
rect 3080 8690 3100 8730
rect 3020 8670 3100 8690
rect 3180 9030 3360 9050
rect 3180 8990 3200 9030
rect 3240 8990 3300 9030
rect 3340 8990 3360 9030
rect 3180 8930 3360 8990
rect 3180 8890 3200 8930
rect 3240 8890 3300 8930
rect 3340 8890 3360 8930
rect 3180 8830 3360 8890
rect 3180 8790 3200 8830
rect 3240 8790 3300 8830
rect 3340 8790 3360 8830
rect 3180 8730 3360 8790
rect 3180 8690 3200 8730
rect 3240 8690 3300 8730
rect 3340 8690 3360 8730
rect 3180 8670 3360 8690
rect 3410 9030 3490 9050
rect 3410 8990 3430 9030
rect 3470 8990 3490 9030
rect 3410 8930 3490 8990
rect 3410 8890 3430 8930
rect 3470 8890 3490 8930
rect 3410 8830 3490 8890
rect 3410 8790 3430 8830
rect 3470 8790 3490 8830
rect 3410 8730 3490 8790
rect 3410 8690 3430 8730
rect 3470 8690 3490 8730
rect 3410 8670 3490 8690
rect 3570 9030 3650 9050
rect 3570 8990 3590 9030
rect 3630 8990 3650 9030
rect 3570 8930 3650 8990
rect 3570 8890 3590 8930
rect 3630 8890 3650 8930
rect 3570 8830 3650 8890
rect 3570 8790 3590 8830
rect 3630 8790 3650 8830
rect 3570 8730 3650 8790
rect 3570 8690 3590 8730
rect 3630 8690 3650 8730
rect 3570 8670 3650 8690
rect 3700 9030 3780 9050
rect 3700 8990 3720 9030
rect 3760 8990 3780 9030
rect 3700 8930 3780 8990
rect 3700 8890 3720 8930
rect 3760 8890 3780 8930
rect 3700 8830 3780 8890
rect 3700 8790 3720 8830
rect 3760 8790 3780 8830
rect 7920 8810 8000 8830
rect 3700 8730 3780 8790
rect 3700 8690 3720 8730
rect 3760 8690 3780 8730
rect 3700 8670 3780 8690
rect 5890 8770 5970 8790
rect 5890 8730 5910 8770
rect 5950 8730 5970 8770
rect 800 8630 840 8670
rect 800 8590 950 8630
rect 1300 8600 1340 8670
rect 1630 8600 1670 8670
rect 1960 8600 2000 8670
rect 2650 8630 2690 8670
rect 2910 8630 2950 8670
rect 470 8530 750 8550
rect 470 8490 490 8530
rect 530 8510 750 8530
rect 530 8490 550 8510
rect 470 8470 550 8490
rect 910 8430 950 8590
rect 1160 8580 1340 8600
rect 1160 8540 1180 8580
rect 1220 8540 1260 8580
rect 1300 8540 1340 8580
rect 1160 8520 1340 8540
rect 1570 8580 1670 8600
rect 1570 8540 1590 8580
rect 1630 8540 1670 8580
rect 1570 8520 1670 8540
rect 1900 8580 2000 8600
rect 1900 8540 1920 8580
rect 1960 8540 2000 8580
rect 1900 8520 2000 8540
rect 2190 8580 2270 8600
rect 2650 8590 2950 8630
rect 2190 8540 2210 8580
rect 2250 8540 2270 8580
rect 2190 8520 2270 8540
rect 2340 8570 2420 8590
rect 2340 8530 2360 8570
rect 2400 8530 2420 8570
rect 1300 8430 1340 8520
rect 1630 8430 1670 8520
rect 1960 8430 2000 8520
rect 2340 8510 2420 8530
rect 2650 8430 2690 8590
rect 2910 8430 2950 8590
rect 3040 8620 3080 8670
rect 3040 8600 3140 8620
rect 3040 8560 3080 8600
rect 3120 8560 3140 8600
rect 3040 8540 3140 8560
rect 3040 8430 3080 8540
rect 3450 8530 3490 8670
rect 3450 8520 3530 8530
rect 3450 8480 3470 8520
rect 3510 8480 3530 8520
rect 3450 8460 3530 8480
rect 3450 8430 3490 8460
rect 3590 8430 3630 8670
rect 3720 8550 3760 8670
rect 5350 8660 5530 8680
rect 5350 8620 5370 8660
rect 5410 8620 5470 8660
rect 5510 8620 5530 8660
rect 5350 8560 5530 8620
rect 3720 8530 4190 8550
rect 3720 8510 4130 8530
rect 3720 8430 3760 8510
rect 4110 8490 4130 8510
rect 4170 8490 4190 8530
rect 4110 8470 4190 8490
rect 5350 8520 5370 8560
rect 5410 8520 5470 8560
rect 5510 8520 5530 8560
rect 4110 8430 4150 8470
rect 5350 8460 5530 8520
rect -710 8410 -570 8430
rect -710 8370 -700 8410
rect -660 8370 -620 8410
rect -580 8370 -570 8410
rect -710 8310 -570 8370
rect -710 8270 -700 8310
rect -660 8270 -620 8310
rect -580 8270 -570 8310
rect -710 8250 -570 8270
rect -520 8410 -460 8430
rect -520 8370 -510 8410
rect -470 8370 -460 8410
rect -520 8310 -460 8370
rect -520 8270 -510 8310
rect -470 8270 -460 8310
rect -520 8250 -460 8270
rect -410 8410 -350 8430
rect -410 8370 -400 8410
rect -360 8370 -350 8410
rect -410 8310 -350 8370
rect -410 8270 -400 8310
rect -360 8270 -350 8310
rect -410 8250 -350 8270
rect -110 8410 -50 8430
rect -110 8370 -100 8410
rect -60 8370 -50 8410
rect -110 8310 -50 8370
rect -110 8270 -100 8310
rect -60 8270 -50 8310
rect -110 8250 -50 8270
rect 0 8410 60 8430
rect 0 8370 10 8410
rect 50 8370 60 8410
rect 0 8310 60 8370
rect 0 8270 10 8310
rect 50 8270 60 8310
rect 0 8250 60 8270
rect 110 8410 330 8430
rect 110 8370 120 8410
rect 160 8370 200 8410
rect 240 8370 280 8410
rect 320 8370 330 8410
rect 110 8310 330 8370
rect 110 8270 120 8310
rect 160 8270 200 8310
rect 240 8270 280 8310
rect 320 8270 330 8310
rect 110 8250 330 8270
rect 380 8410 440 8430
rect 380 8370 390 8410
rect 430 8370 440 8410
rect 380 8310 440 8370
rect 380 8270 390 8310
rect 430 8270 440 8310
rect 380 8250 440 8270
rect 490 8410 550 8430
rect 490 8370 500 8410
rect 540 8370 550 8410
rect 490 8310 550 8370
rect 490 8270 500 8310
rect 540 8270 550 8310
rect 490 8250 550 8270
rect 790 8410 850 8430
rect 790 8370 800 8410
rect 840 8370 850 8410
rect 790 8310 850 8370
rect 790 8270 800 8310
rect 840 8270 850 8310
rect 790 8250 850 8270
rect 900 8410 960 8430
rect 900 8370 910 8410
rect 950 8370 960 8410
rect 900 8310 960 8370
rect 900 8270 910 8310
rect 950 8270 960 8310
rect 900 8250 960 8270
rect 1010 8410 1150 8430
rect 1010 8370 1020 8410
rect 1060 8370 1100 8410
rect 1140 8370 1150 8410
rect 1010 8310 1150 8370
rect 1010 8270 1020 8310
rect 1060 8270 1100 8310
rect 1140 8270 1150 8310
rect 1010 8250 1150 8270
rect 1300 8410 1360 8430
rect 1300 8370 1310 8410
rect 1350 8370 1360 8410
rect 1300 8310 1360 8370
rect 1300 8270 1310 8310
rect 1350 8270 1360 8310
rect 1300 8250 1360 8270
rect 1410 8410 1550 8430
rect 1410 8370 1420 8410
rect 1460 8370 1500 8410
rect 1540 8370 1550 8410
rect 1410 8310 1550 8370
rect 1410 8270 1420 8310
rect 1460 8270 1500 8310
rect 1540 8270 1550 8310
rect 1410 8250 1550 8270
rect 1630 8410 1690 8430
rect 1630 8370 1640 8410
rect 1680 8370 1690 8410
rect 1630 8310 1690 8370
rect 1630 8270 1640 8310
rect 1680 8270 1690 8310
rect 1630 8250 1690 8270
rect 1740 8410 1880 8430
rect 1740 8370 1750 8410
rect 1790 8370 1830 8410
rect 1870 8370 1880 8410
rect 1740 8310 1880 8370
rect 1740 8270 1750 8310
rect 1790 8270 1830 8310
rect 1870 8270 1880 8310
rect 1740 8250 1880 8270
rect 1960 8410 2020 8430
rect 1960 8370 1970 8410
rect 2010 8370 2020 8410
rect 1960 8310 2020 8370
rect 1960 8270 1970 8310
rect 2010 8270 2020 8310
rect 1960 8250 2020 8270
rect 2070 8410 2210 8430
rect 2070 8370 2080 8410
rect 2120 8370 2160 8410
rect 2200 8370 2210 8410
rect 2070 8310 2210 8370
rect 2070 8270 2080 8310
rect 2120 8270 2160 8310
rect 2200 8270 2210 8310
rect 2070 8250 2210 8270
rect 2400 8410 2580 8430
rect 2400 8370 2420 8410
rect 2460 8370 2520 8410
rect 2560 8370 2580 8410
rect 2400 8310 2580 8370
rect 2400 8270 2420 8310
rect 2460 8270 2520 8310
rect 2560 8270 2580 8310
rect 2400 8250 2580 8270
rect 2630 8410 2710 8430
rect 2630 8370 2650 8410
rect 2690 8370 2710 8410
rect 2630 8310 2710 8370
rect 2630 8270 2650 8310
rect 2690 8270 2710 8310
rect 2630 8250 2710 8270
rect 2890 8410 2970 8430
rect 2890 8370 2910 8410
rect 2950 8370 2970 8410
rect 2890 8310 2970 8370
rect 2890 8270 2910 8310
rect 2950 8270 2970 8310
rect 2890 8250 2970 8270
rect 3020 8410 3100 8430
rect 3020 8370 3040 8410
rect 3080 8370 3100 8410
rect 3020 8310 3100 8370
rect 3020 8270 3040 8310
rect 3080 8270 3100 8310
rect 3020 8250 3100 8270
rect 3180 8410 3360 8430
rect 3180 8370 3200 8410
rect 3240 8370 3300 8410
rect 3340 8370 3360 8410
rect 3180 8310 3360 8370
rect 3180 8270 3200 8310
rect 3240 8270 3300 8310
rect 3340 8270 3360 8310
rect 3180 8250 3360 8270
rect 3410 8410 3490 8430
rect 3410 8370 3430 8410
rect 3470 8370 3490 8410
rect 3410 8310 3490 8370
rect 3410 8270 3430 8310
rect 3470 8270 3490 8310
rect 3410 8250 3490 8270
rect 3570 8410 3650 8430
rect 3570 8370 3590 8410
rect 3630 8370 3650 8410
rect 3570 8310 3650 8370
rect 3570 8270 3590 8310
rect 3630 8270 3650 8310
rect 3570 8250 3650 8270
rect 3700 8410 3780 8430
rect 3700 8370 3720 8410
rect 3760 8370 3780 8410
rect 3700 8310 3780 8370
rect 3700 8270 3720 8310
rect 3760 8270 3780 8310
rect 3700 8250 3780 8270
rect 3860 8410 4040 8430
rect 3860 8370 3880 8410
rect 3920 8370 3980 8410
rect 4020 8370 4040 8410
rect 3860 8310 4040 8370
rect 3860 8270 3880 8310
rect 3920 8270 3980 8310
rect 4020 8270 4040 8310
rect 3860 8250 4040 8270
rect 4090 8410 4170 8430
rect 4090 8370 4110 8410
rect 4150 8370 4170 8410
rect 4090 8310 4170 8370
rect 4090 8270 4110 8310
rect 4150 8270 4170 8310
rect 5350 8420 5370 8460
rect 5410 8420 5470 8460
rect 5510 8420 5530 8460
rect 5350 8360 5530 8420
rect 5350 8320 5370 8360
rect 5410 8320 5470 8360
rect 5510 8320 5530 8360
rect 5350 8300 5530 8320
rect 5670 8660 5750 8680
rect 5670 8620 5690 8660
rect 5730 8620 5750 8660
rect 5670 8560 5750 8620
rect 5670 8520 5690 8560
rect 5730 8520 5750 8560
rect 5670 8460 5750 8520
rect 5670 8420 5690 8460
rect 5730 8420 5750 8460
rect 5670 8360 5750 8420
rect 5670 8320 5690 8360
rect 5730 8320 5750 8360
rect 5670 8300 5750 8320
rect 5890 8660 5970 8730
rect 6430 8780 6510 8800
rect 6430 8740 6450 8780
rect 6490 8740 6510 8780
rect 6430 8680 6510 8740
rect 7510 8780 7590 8800
rect 7510 8740 7530 8780
rect 7570 8740 7590 8780
rect 7920 8770 7940 8810
rect 7980 8770 8000 8810
rect 7920 8750 8000 8770
rect 8180 8810 8260 8830
rect 8180 8770 8200 8810
rect 8240 8770 8260 8810
rect 8180 8750 8260 8770
rect 8850 8810 8960 8830
rect 7510 8680 7590 8740
rect 8850 8740 8870 8810
rect 8940 8740 8960 8810
rect 8850 8720 8960 8740
rect 5890 8620 5910 8660
rect 5950 8620 5970 8660
rect 5890 8560 5970 8620
rect 5890 8520 5910 8560
rect 5950 8520 5970 8560
rect 5890 8460 5970 8520
rect 5890 8420 5910 8460
rect 5950 8420 5970 8460
rect 5890 8360 5970 8420
rect 5890 8320 5910 8360
rect 5950 8320 5970 8360
rect 5890 8300 5970 8320
rect 6110 8660 6190 8680
rect 6110 8620 6130 8660
rect 6170 8620 6190 8660
rect 6110 8560 6190 8620
rect 6110 8520 6130 8560
rect 6170 8520 6190 8560
rect 6110 8460 6190 8520
rect 6110 8420 6130 8460
rect 6170 8420 6190 8460
rect 6110 8360 6190 8420
rect 6110 8320 6130 8360
rect 6170 8320 6190 8360
rect 6110 8300 6190 8320
rect 6330 8660 6610 8680
rect 6330 8620 6350 8660
rect 6390 8620 6450 8660
rect 6490 8620 6550 8660
rect 6590 8620 6610 8660
rect 6330 8560 6610 8620
rect 6330 8520 6350 8560
rect 6390 8520 6450 8560
rect 6490 8520 6550 8560
rect 6590 8520 6610 8560
rect 6330 8460 6610 8520
rect 6330 8420 6350 8460
rect 6390 8420 6450 8460
rect 6490 8420 6550 8460
rect 6590 8420 6610 8460
rect 6330 8360 6610 8420
rect 6330 8320 6350 8360
rect 6390 8320 6450 8360
rect 6490 8320 6550 8360
rect 6590 8320 6610 8360
rect 6330 8300 6610 8320
rect 6750 8660 6830 8680
rect 6750 8620 6770 8660
rect 6810 8620 6830 8660
rect 6750 8560 6830 8620
rect 6750 8520 6770 8560
rect 6810 8520 6830 8560
rect 6750 8460 6830 8520
rect 6750 8420 6770 8460
rect 6810 8420 6830 8460
rect 6750 8360 6830 8420
rect 6750 8320 6770 8360
rect 6810 8320 6830 8360
rect 6750 8300 6830 8320
rect 6970 8660 7050 8680
rect 6970 8620 6990 8660
rect 7030 8620 7050 8660
rect 6970 8560 7050 8620
rect 6970 8520 6990 8560
rect 7030 8520 7050 8560
rect 6970 8460 7050 8520
rect 6970 8420 6990 8460
rect 7030 8420 7050 8460
rect 6970 8360 7050 8420
rect 6970 8320 6990 8360
rect 7030 8320 7050 8360
rect 6970 8300 7050 8320
rect 7190 8660 7270 8680
rect 7190 8620 7210 8660
rect 7250 8620 7270 8660
rect 7190 8560 7270 8620
rect 7190 8520 7210 8560
rect 7250 8520 7270 8560
rect 7190 8460 7270 8520
rect 7190 8420 7210 8460
rect 7250 8420 7270 8460
rect 7190 8360 7270 8420
rect 7190 8320 7210 8360
rect 7250 8320 7270 8360
rect 7190 8300 7270 8320
rect 7410 8660 7690 8680
rect 7410 8620 7430 8660
rect 7470 8620 7530 8660
rect 7570 8620 7630 8660
rect 7670 8620 7690 8660
rect 7410 8560 7690 8620
rect 7410 8520 7430 8560
rect 7470 8520 7530 8560
rect 7570 8520 7630 8560
rect 7670 8520 7690 8560
rect 7410 8460 7690 8520
rect 7410 8420 7430 8460
rect 7470 8420 7530 8460
rect 7570 8420 7630 8460
rect 7670 8420 7690 8460
rect 7410 8360 7690 8420
rect 7410 8320 7430 8360
rect 7470 8320 7530 8360
rect 7570 8320 7630 8360
rect 7670 8320 7690 8360
rect 7410 8300 7690 8320
rect 7830 8660 7910 8680
rect 7830 8620 7850 8660
rect 7890 8620 7910 8660
rect 7830 8560 7910 8620
rect 7830 8520 7850 8560
rect 7890 8520 7910 8560
rect 7830 8460 7910 8520
rect 7830 8420 7850 8460
rect 7890 8420 7910 8460
rect 7830 8360 7910 8420
rect 7830 8320 7850 8360
rect 7890 8320 7910 8360
rect 7830 8300 7910 8320
rect 8050 8660 8130 8680
rect 8050 8620 8070 8660
rect 8110 8620 8130 8660
rect 8050 8560 8130 8620
rect 8050 8520 8070 8560
rect 8110 8520 8130 8560
rect 8050 8460 8130 8520
rect 8050 8420 8070 8460
rect 8110 8420 8130 8460
rect 8050 8360 8130 8420
rect 8050 8320 8070 8360
rect 8110 8320 8130 8360
rect 8050 8300 8130 8320
rect 8270 8660 8350 8680
rect 8270 8620 8290 8660
rect 8330 8620 8350 8660
rect 8270 8560 8350 8620
rect 8270 8520 8290 8560
rect 8330 8520 8350 8560
rect 8270 8460 8350 8520
rect 8270 8420 8290 8460
rect 8330 8420 8350 8460
rect 8270 8360 8350 8420
rect 8270 8320 8290 8360
rect 8330 8320 8350 8360
rect 8270 8300 8350 8320
rect 8490 8660 8670 8680
rect 8490 8620 8510 8660
rect 8550 8620 8610 8660
rect 8650 8620 8670 8660
rect 8490 8560 8670 8620
rect 8490 8520 8510 8560
rect 8550 8520 8610 8560
rect 8650 8520 8670 8560
rect 8490 8460 8670 8520
rect 8490 8420 8510 8460
rect 8550 8420 8610 8460
rect 8650 8420 8670 8460
rect 8490 8360 8670 8420
rect 8490 8320 8510 8360
rect 8550 8320 8610 8360
rect 8650 8320 8670 8360
rect 8490 8300 8670 8320
rect 4090 8250 4170 8270
rect -620 8100 -580 8250
rect -400 8100 -360 8250
rect -100 8100 -60 8250
rect 130 8100 170 8250
rect 280 8100 320 8250
rect 500 8100 540 8250
rect 800 8100 840 8250
rect 1020 8100 1060 8250
rect 1420 8100 1460 8250
rect 1750 8100 1790 8250
rect 2080 8100 2120 8250
rect 2520 8100 2560 8250
rect 3010 8190 3090 8210
rect 3010 8150 3030 8190
rect 3070 8150 3090 8190
rect 3010 8130 3090 8150
rect 3300 8100 3340 8250
rect 3640 8190 3720 8210
rect 3640 8150 3660 8190
rect 3700 8150 3720 8190
rect 3640 8130 3720 8150
rect 3980 8100 4020 8250
rect 5450 8240 5530 8260
rect 5450 8200 5470 8240
rect 5510 8200 5530 8240
rect 5450 8180 5530 8200
rect 8490 8240 8570 8260
rect 8490 8200 8510 8240
rect 8550 8200 8570 8240
rect 8490 8180 8570 8200
rect -640 8080 -560 8100
rect -640 8040 -620 8080
rect -580 8040 -560 8080
rect -640 8020 -560 8040
rect -420 8080 -340 8100
rect -420 8040 -400 8080
rect -360 8040 -340 8080
rect -420 8020 -340 8040
rect -120 8080 -40 8100
rect -120 8040 -100 8080
rect -60 8040 -40 8080
rect -120 8020 -40 8040
rect 110 8080 190 8100
rect 110 8040 130 8080
rect 170 8040 190 8080
rect 110 8020 190 8040
rect 260 8080 340 8100
rect 260 8040 280 8080
rect 320 8040 340 8080
rect 260 8020 340 8040
rect 480 8080 560 8100
rect 480 8040 500 8080
rect 540 8040 560 8080
rect 480 8020 560 8040
rect 780 8080 860 8100
rect 780 8040 800 8080
rect 840 8040 860 8080
rect 780 8020 860 8040
rect 1000 8080 1080 8100
rect 1000 8040 1020 8080
rect 1060 8040 1080 8080
rect 1000 8020 1080 8040
rect 1400 8080 1480 8100
rect 1400 8040 1420 8080
rect 1460 8040 1480 8080
rect 1400 8020 1480 8040
rect 1730 8080 1810 8100
rect 1730 8040 1750 8080
rect 1790 8040 1810 8080
rect 1730 8020 1810 8040
rect 2060 8080 2140 8100
rect 2060 8040 2080 8080
rect 2120 8040 2140 8080
rect 2060 8020 2140 8040
rect 2500 8080 2580 8100
rect 2500 8040 2520 8080
rect 2560 8040 2580 8080
rect 2500 8020 2580 8040
rect 3280 8080 3360 8100
rect 3280 8040 3300 8080
rect 3340 8040 3360 8080
rect 3280 8020 3360 8040
rect 3960 8080 4040 8100
rect 3960 8040 3980 8080
rect 4020 8040 4040 8080
rect 3960 8020 4040 8040
rect 9200 8020 9310 8040
rect 9200 7950 9220 8020
rect 9290 7950 9310 8020
rect 9200 7930 9310 7950
rect 9320 7260 9420 7280
rect 9320 7200 9340 7260
rect 9400 7200 9420 7260
rect 9320 7180 9420 7200
rect -1360 6960 -1280 6980
rect -1360 6920 -1340 6960
rect -1300 6920 -1280 6960
rect -1360 6900 -1280 6920
rect -40 6960 40 6980
rect -40 6920 -20 6960
rect 20 6920 40 6960
rect -40 6900 40 6920
rect 540 6960 620 6980
rect 540 6920 560 6960
rect 600 6920 620 6960
rect 540 6900 620 6920
rect 1860 6960 1940 6980
rect 1860 6920 1880 6960
rect 1920 6920 1940 6960
rect 1860 6900 1940 6920
rect -1430 6840 -1290 6860
rect -1430 6800 -1420 6840
rect -1380 6800 -1340 6840
rect -1300 6800 -1290 6840
rect -1430 6740 -1290 6800
rect -1430 6700 -1420 6740
rect -1380 6700 -1340 6740
rect -1300 6700 -1290 6740
rect -1430 6680 -1290 6700
rect -1240 6840 -1180 6860
rect -1240 6800 -1230 6840
rect -1190 6800 -1180 6840
rect -1240 6740 -1180 6800
rect -1240 6700 -1230 6740
rect -1190 6700 -1180 6740
rect -1240 6680 -1180 6700
rect -1130 6840 -1070 6860
rect -1130 6800 -1120 6840
rect -1080 6800 -1070 6840
rect -1130 6740 -1070 6800
rect -1130 6700 -1120 6740
rect -1080 6700 -1070 6740
rect -1130 6680 -1070 6700
rect -1020 6840 -960 6860
rect -1020 6800 -1010 6840
rect -970 6800 -960 6840
rect -1020 6740 -960 6800
rect -1020 6700 -1010 6740
rect -970 6700 -960 6740
rect -1020 6680 -960 6700
rect -910 6840 -850 6860
rect -910 6800 -900 6840
rect -860 6800 -850 6840
rect -910 6740 -850 6800
rect -910 6700 -900 6740
rect -860 6700 -850 6740
rect -910 6680 -850 6700
rect -800 6840 -740 6860
rect -800 6800 -790 6840
rect -750 6800 -740 6840
rect -800 6740 -740 6800
rect -800 6700 -790 6740
rect -750 6700 -740 6740
rect -800 6680 -740 6700
rect -690 6840 -630 6860
rect -690 6800 -680 6840
rect -640 6800 -630 6840
rect -690 6740 -630 6800
rect -690 6700 -680 6740
rect -640 6700 -630 6740
rect -690 6680 -630 6700
rect -580 6840 -520 6860
rect -580 6800 -570 6840
rect -530 6800 -520 6840
rect -580 6740 -520 6800
rect -580 6700 -570 6740
rect -530 6700 -520 6740
rect -580 6680 -520 6700
rect -470 6840 -410 6860
rect -470 6800 -460 6840
rect -420 6800 -410 6840
rect -470 6740 -410 6800
rect -470 6700 -460 6740
rect -420 6700 -410 6740
rect -470 6680 -410 6700
rect -360 6840 -300 6860
rect -360 6800 -350 6840
rect -310 6800 -300 6840
rect -360 6740 -300 6800
rect -360 6700 -350 6740
rect -310 6700 -300 6740
rect -360 6680 -300 6700
rect -250 6840 -190 6860
rect -250 6800 -240 6840
rect -200 6800 -190 6840
rect -250 6740 -190 6800
rect -250 6700 -240 6740
rect -200 6700 -190 6740
rect -250 6680 -190 6700
rect -140 6840 -80 6860
rect -140 6800 -130 6840
rect -90 6800 -80 6840
rect -140 6740 -80 6800
rect -140 6700 -130 6740
rect -90 6700 -80 6740
rect -140 6680 -80 6700
rect -30 6840 110 6860
rect -30 6800 -20 6840
rect 20 6800 60 6840
rect 100 6800 110 6840
rect -30 6740 110 6800
rect -30 6700 -20 6740
rect 20 6700 60 6740
rect 100 6700 110 6740
rect -30 6680 110 6700
rect 470 6840 610 6860
rect 470 6800 480 6840
rect 520 6800 560 6840
rect 600 6800 610 6840
rect 470 6740 610 6800
rect 470 6700 480 6740
rect 520 6700 560 6740
rect 600 6700 610 6740
rect 470 6680 610 6700
rect 660 6840 720 6860
rect 660 6800 670 6840
rect 710 6800 720 6840
rect 660 6740 720 6800
rect 660 6700 670 6740
rect 710 6700 720 6740
rect 660 6680 720 6700
rect 770 6840 830 6860
rect 770 6800 780 6840
rect 820 6800 830 6840
rect 770 6740 830 6800
rect 770 6700 780 6740
rect 820 6700 830 6740
rect 770 6680 830 6700
rect 880 6840 940 6860
rect 880 6800 890 6840
rect 930 6800 940 6840
rect 880 6740 940 6800
rect 880 6700 890 6740
rect 930 6700 940 6740
rect 880 6680 940 6700
rect 990 6840 1050 6860
rect 990 6800 1000 6840
rect 1040 6800 1050 6840
rect 990 6740 1050 6800
rect 990 6700 1000 6740
rect 1040 6700 1050 6740
rect 990 6680 1050 6700
rect 1100 6840 1160 6860
rect 1100 6800 1110 6840
rect 1150 6800 1160 6840
rect 1100 6740 1160 6800
rect 1100 6700 1110 6740
rect 1150 6700 1160 6740
rect 1100 6680 1160 6700
rect 1210 6840 1270 6860
rect 1210 6800 1220 6840
rect 1260 6800 1270 6840
rect 1210 6740 1270 6800
rect 1210 6700 1220 6740
rect 1260 6700 1270 6740
rect 1210 6680 1270 6700
rect 1320 6840 1380 6860
rect 1320 6800 1330 6840
rect 1370 6800 1380 6840
rect 1320 6740 1380 6800
rect 1320 6700 1330 6740
rect 1370 6700 1380 6740
rect 1320 6680 1380 6700
rect 1430 6840 1490 6860
rect 1430 6800 1440 6840
rect 1480 6800 1490 6840
rect 1430 6740 1490 6800
rect 1430 6700 1440 6740
rect 1480 6700 1490 6740
rect 1430 6680 1490 6700
rect 1540 6840 1600 6860
rect 1540 6800 1550 6840
rect 1590 6800 1600 6840
rect 1540 6740 1600 6800
rect 1540 6700 1550 6740
rect 1590 6700 1600 6740
rect 1540 6680 1600 6700
rect 1650 6840 1710 6860
rect 1650 6800 1660 6840
rect 1700 6800 1710 6840
rect 1650 6740 1710 6800
rect 1650 6700 1660 6740
rect 1700 6700 1710 6740
rect 1650 6680 1710 6700
rect 1760 6840 1820 6860
rect 1760 6800 1770 6840
rect 1810 6800 1820 6840
rect 1760 6740 1820 6800
rect 1760 6700 1770 6740
rect 1810 6700 1820 6740
rect 1760 6680 1820 6700
rect 1870 6840 2010 6860
rect 1870 6800 1880 6840
rect 1920 6800 1960 6840
rect 2000 6800 2010 6840
rect 1870 6740 2010 6800
rect 1870 6700 1880 6740
rect 1920 6700 1960 6740
rect 2000 6700 2010 6740
rect 1870 6680 2010 6700
rect 9120 6730 9200 6750
rect 9120 6690 9140 6730
rect 9180 6690 9200 6730
rect 9120 6670 9200 6690
rect -1184 6622 -1126 6640
rect -1184 6588 -1172 6622
rect -1138 6588 -1126 6622
rect -1184 6570 -1126 6588
rect -1074 6622 -1016 6640
rect -1074 6588 -1062 6622
rect -1028 6588 -1016 6622
rect -1074 6570 -1016 6588
rect -964 6622 -906 6640
rect -964 6588 -952 6622
rect -918 6588 -906 6622
rect -964 6570 -906 6588
rect -854 6622 -796 6640
rect -854 6588 -842 6622
rect -808 6588 -796 6622
rect -854 6570 -796 6588
rect -744 6622 -686 6640
rect -744 6588 -732 6622
rect -698 6588 -686 6622
rect -744 6570 -686 6588
rect -634 6622 -576 6640
rect -634 6588 -622 6622
rect -588 6588 -576 6622
rect -634 6570 -576 6588
rect -524 6622 -466 6640
rect -524 6588 -512 6622
rect -478 6588 -466 6622
rect -524 6570 -466 6588
rect -414 6622 -356 6640
rect -414 6588 -402 6622
rect -368 6588 -356 6622
rect -414 6570 -356 6588
rect -304 6622 -246 6640
rect -304 6588 -292 6622
rect -258 6588 -246 6622
rect -304 6570 -246 6588
rect -194 6622 -136 6640
rect -194 6588 -182 6622
rect -148 6588 -136 6622
rect -194 6570 -136 6588
rect 716 6622 774 6640
rect 716 6588 728 6622
rect 762 6588 774 6622
rect 716 6570 774 6588
rect 826 6622 884 6640
rect 826 6588 838 6622
rect 872 6588 884 6622
rect 826 6570 884 6588
rect 936 6622 994 6640
rect 936 6588 948 6622
rect 982 6588 994 6622
rect 936 6570 994 6588
rect 1046 6622 1104 6640
rect 1046 6588 1058 6622
rect 1092 6588 1104 6622
rect 1046 6570 1104 6588
rect 1156 6622 1214 6640
rect 1156 6588 1168 6622
rect 1202 6588 1214 6622
rect 1156 6570 1214 6588
rect 1266 6622 1324 6640
rect 1266 6588 1278 6622
rect 1312 6588 1324 6622
rect 1266 6570 1324 6588
rect 1376 6622 1434 6640
rect 1376 6588 1388 6622
rect 1422 6588 1434 6622
rect 1376 6570 1434 6588
rect 1486 6622 1544 6640
rect 1486 6588 1498 6622
rect 1532 6588 1544 6622
rect 1486 6570 1544 6588
rect 1596 6622 1654 6640
rect 1596 6588 1608 6622
rect 1642 6588 1654 6622
rect 1596 6570 1654 6588
rect 1706 6622 1764 6640
rect 1706 6588 1718 6622
rect 1752 6588 1764 6622
rect 1706 6570 1764 6588
rect -1370 6360 -1290 6380
rect -1370 6320 -1350 6360
rect -1310 6320 -1290 6360
rect -1370 6300 -1290 6320
rect -1010 6360 -930 6380
rect -1010 6320 -990 6360
rect -950 6320 -930 6360
rect -1010 6300 -930 6320
rect -650 6360 -570 6380
rect -650 6320 -630 6360
rect -590 6320 -570 6360
rect -650 6300 -570 6320
rect -290 6360 -210 6380
rect -290 6320 -270 6360
rect -230 6320 -210 6360
rect -290 6300 -210 6320
rect 70 6360 150 6380
rect 70 6320 90 6360
rect 130 6320 150 6360
rect 70 6300 150 6320
rect 430 6360 510 6380
rect 430 6320 450 6360
rect 490 6320 510 6360
rect 430 6300 510 6320
rect 790 6360 870 6380
rect 790 6320 810 6360
rect 850 6320 870 6360
rect 790 6300 870 6320
rect 1150 6360 1230 6380
rect 1150 6320 1170 6360
rect 1210 6320 1230 6360
rect 1150 6300 1230 6320
rect 1510 6360 1590 6380
rect 1510 6320 1530 6360
rect 1570 6320 1590 6360
rect 1510 6300 1590 6320
rect 1870 6360 1950 6380
rect 1870 6320 1890 6360
rect 1930 6320 1950 6360
rect 1870 6300 1950 6320
rect 5250 6356 5370 6360
rect 6670 6356 6790 6360
rect 5250 6340 5404 6356
rect 5250 6300 5270 6340
rect 5310 6306 5370 6340
rect 5310 6300 5404 6306
rect -1350 6260 -1310 6300
rect -990 6260 -950 6300
rect -630 6260 -590 6300
rect -270 6260 -230 6300
rect 90 6260 130 6300
rect 450 6260 490 6300
rect 810 6260 850 6300
rect 1170 6260 1210 6300
rect 1530 6260 1570 6300
rect 1890 6260 1930 6300
rect 5250 6290 5404 6300
rect 6644 6340 6790 6356
rect 6678 6306 6790 6340
rect 6644 6290 6790 6306
rect 5250 6280 5370 6290
rect -1440 6240 -1300 6260
rect -1440 6200 -1430 6240
rect -1390 6200 -1350 6240
rect -1310 6200 -1300 6240
rect -1440 6140 -1300 6200
rect -1440 6100 -1430 6140
rect -1390 6100 -1350 6140
rect -1310 6100 -1300 6140
rect -1440 6040 -1300 6100
rect -1440 6000 -1430 6040
rect -1390 6000 -1350 6040
rect -1310 6000 -1300 6040
rect -1440 5940 -1300 6000
rect -1440 5900 -1430 5940
rect -1390 5900 -1350 5940
rect -1310 5900 -1300 5940
rect -1440 5840 -1300 5900
rect -1440 5800 -1430 5840
rect -1390 5800 -1350 5840
rect -1310 5800 -1300 5840
rect -1440 5740 -1300 5800
rect -1440 5700 -1430 5740
rect -1390 5700 -1350 5740
rect -1310 5700 -1300 5740
rect -1440 5680 -1300 5700
rect -1180 6240 -1120 6260
rect -1180 6200 -1170 6240
rect -1130 6200 -1120 6240
rect -1180 6140 -1120 6200
rect -1180 6100 -1170 6140
rect -1130 6100 -1120 6140
rect -1180 6040 -1120 6100
rect -1180 6000 -1170 6040
rect -1130 6000 -1120 6040
rect -1180 5940 -1120 6000
rect -1180 5900 -1170 5940
rect -1130 5900 -1120 5940
rect -1180 5840 -1120 5900
rect -1180 5800 -1170 5840
rect -1130 5800 -1120 5840
rect -1180 5740 -1120 5800
rect -1180 5700 -1170 5740
rect -1130 5700 -1120 5740
rect -1180 5680 -1120 5700
rect -1000 6240 -940 6260
rect -1000 6200 -990 6240
rect -950 6200 -940 6240
rect -1000 6140 -940 6200
rect -1000 6100 -990 6140
rect -950 6100 -940 6140
rect -1000 6040 -940 6100
rect -1000 6000 -990 6040
rect -950 6000 -940 6040
rect -1000 5940 -940 6000
rect -1000 5900 -990 5940
rect -950 5900 -940 5940
rect -1000 5840 -940 5900
rect -1000 5800 -990 5840
rect -950 5800 -940 5840
rect -1000 5740 -940 5800
rect -1000 5700 -990 5740
rect -950 5700 -940 5740
rect -1000 5680 -940 5700
rect -820 6240 -760 6260
rect -820 6200 -810 6240
rect -770 6200 -760 6240
rect -820 6140 -760 6200
rect -820 6100 -810 6140
rect -770 6100 -760 6140
rect -820 6040 -760 6100
rect -820 6000 -810 6040
rect -770 6000 -760 6040
rect -820 5940 -760 6000
rect -820 5900 -810 5940
rect -770 5900 -760 5940
rect -820 5840 -760 5900
rect -820 5800 -810 5840
rect -770 5800 -760 5840
rect -820 5740 -760 5800
rect -820 5700 -810 5740
rect -770 5700 -760 5740
rect -820 5680 -760 5700
rect -640 6240 -580 6260
rect -640 6200 -630 6240
rect -590 6200 -580 6240
rect -640 6140 -580 6200
rect -640 6100 -630 6140
rect -590 6100 -580 6140
rect -640 6040 -580 6100
rect -640 6000 -630 6040
rect -590 6000 -580 6040
rect -640 5940 -580 6000
rect -640 5900 -630 5940
rect -590 5900 -580 5940
rect -640 5840 -580 5900
rect -640 5800 -630 5840
rect -590 5800 -580 5840
rect -640 5740 -580 5800
rect -640 5700 -630 5740
rect -590 5700 -580 5740
rect -640 5680 -580 5700
rect -460 6240 -400 6260
rect -460 6200 -450 6240
rect -410 6200 -400 6240
rect -460 6140 -400 6200
rect -460 6100 -450 6140
rect -410 6100 -400 6140
rect -460 6040 -400 6100
rect -460 6000 -450 6040
rect -410 6000 -400 6040
rect -460 5940 -400 6000
rect -460 5900 -450 5940
rect -410 5900 -400 5940
rect -460 5840 -400 5900
rect -460 5800 -450 5840
rect -410 5800 -400 5840
rect -460 5740 -400 5800
rect -460 5700 -450 5740
rect -410 5700 -400 5740
rect -460 5680 -400 5700
rect -280 6240 -220 6260
rect -280 6200 -270 6240
rect -230 6200 -220 6240
rect -280 6140 -220 6200
rect -280 6100 -270 6140
rect -230 6100 -220 6140
rect -280 6040 -220 6100
rect -280 6000 -270 6040
rect -230 6000 -220 6040
rect -280 5940 -220 6000
rect -280 5900 -270 5940
rect -230 5900 -220 5940
rect -280 5840 -220 5900
rect -280 5800 -270 5840
rect -230 5800 -220 5840
rect -280 5740 -220 5800
rect -280 5700 -270 5740
rect -230 5700 -220 5740
rect -280 5680 -220 5700
rect -100 6240 -40 6260
rect -100 6200 -90 6240
rect -50 6200 -40 6240
rect -100 6140 -40 6200
rect -100 6100 -90 6140
rect -50 6100 -40 6140
rect -100 6040 -40 6100
rect -100 6000 -90 6040
rect -50 6000 -40 6040
rect -100 5940 -40 6000
rect -100 5900 -90 5940
rect -50 5900 -40 5940
rect -100 5840 -40 5900
rect -100 5800 -90 5840
rect -50 5800 -40 5840
rect -100 5740 -40 5800
rect -100 5700 -90 5740
rect -50 5700 -40 5740
rect -100 5680 -40 5700
rect 80 6240 140 6260
rect 80 6200 90 6240
rect 130 6200 140 6240
rect 80 6140 140 6200
rect 80 6100 90 6140
rect 130 6100 140 6140
rect 80 6040 140 6100
rect 80 6000 90 6040
rect 130 6000 140 6040
rect 80 5940 140 6000
rect 80 5900 90 5940
rect 130 5900 140 5940
rect 80 5840 140 5900
rect 80 5800 90 5840
rect 130 5800 140 5840
rect 80 5740 140 5800
rect 80 5700 90 5740
rect 130 5700 140 5740
rect 80 5680 140 5700
rect 260 6240 320 6260
rect 260 6200 270 6240
rect 310 6200 320 6240
rect 260 6140 320 6200
rect 260 6100 270 6140
rect 310 6100 320 6140
rect 260 6040 320 6100
rect 260 6000 270 6040
rect 310 6000 320 6040
rect 260 5940 320 6000
rect 260 5900 270 5940
rect 310 5900 320 5940
rect 260 5840 320 5900
rect 260 5800 270 5840
rect 310 5800 320 5840
rect 260 5740 320 5800
rect 260 5700 270 5740
rect 310 5700 320 5740
rect 260 5680 320 5700
rect 440 6240 500 6260
rect 440 6200 450 6240
rect 490 6200 500 6240
rect 440 6140 500 6200
rect 440 6100 450 6140
rect 490 6100 500 6140
rect 440 6040 500 6100
rect 440 6000 450 6040
rect 490 6000 500 6040
rect 440 5940 500 6000
rect 440 5900 450 5940
rect 490 5900 500 5940
rect 440 5840 500 5900
rect 440 5800 450 5840
rect 490 5800 500 5840
rect 440 5740 500 5800
rect 440 5700 450 5740
rect 490 5700 500 5740
rect 440 5680 500 5700
rect 620 6240 680 6260
rect 620 6200 630 6240
rect 670 6200 680 6240
rect 620 6140 680 6200
rect 620 6100 630 6140
rect 670 6100 680 6140
rect 620 6040 680 6100
rect 620 6000 630 6040
rect 670 6000 680 6040
rect 620 5940 680 6000
rect 620 5900 630 5940
rect 670 5900 680 5940
rect 620 5840 680 5900
rect 620 5800 630 5840
rect 670 5800 680 5840
rect 620 5740 680 5800
rect 620 5700 630 5740
rect 670 5700 680 5740
rect 620 5680 680 5700
rect 800 6240 860 6260
rect 800 6200 810 6240
rect 850 6200 860 6240
rect 800 6140 860 6200
rect 800 6100 810 6140
rect 850 6100 860 6140
rect 800 6040 860 6100
rect 800 6000 810 6040
rect 850 6000 860 6040
rect 800 5940 860 6000
rect 800 5900 810 5940
rect 850 5900 860 5940
rect 800 5840 860 5900
rect 800 5800 810 5840
rect 850 5800 860 5840
rect 800 5740 860 5800
rect 800 5700 810 5740
rect 850 5700 860 5740
rect 800 5680 860 5700
rect 980 6240 1040 6260
rect 980 6200 990 6240
rect 1030 6200 1040 6240
rect 980 6140 1040 6200
rect 980 6100 990 6140
rect 1030 6100 1040 6140
rect 980 6040 1040 6100
rect 980 6000 990 6040
rect 1030 6000 1040 6040
rect 980 5940 1040 6000
rect 980 5900 990 5940
rect 1030 5900 1040 5940
rect 980 5840 1040 5900
rect 980 5800 990 5840
rect 1030 5800 1040 5840
rect 980 5740 1040 5800
rect 980 5700 990 5740
rect 1030 5700 1040 5740
rect 980 5680 1040 5700
rect 1160 6240 1220 6260
rect 1160 6200 1170 6240
rect 1210 6200 1220 6240
rect 1160 6140 1220 6200
rect 1160 6100 1170 6140
rect 1210 6100 1220 6140
rect 1160 6040 1220 6100
rect 1160 6000 1170 6040
rect 1210 6000 1220 6040
rect 1160 5940 1220 6000
rect 1160 5900 1170 5940
rect 1210 5900 1220 5940
rect 1160 5840 1220 5900
rect 1160 5800 1170 5840
rect 1210 5800 1220 5840
rect 1160 5740 1220 5800
rect 1160 5700 1170 5740
rect 1210 5700 1220 5740
rect 1160 5680 1220 5700
rect 1340 6240 1400 6260
rect 1340 6200 1350 6240
rect 1390 6200 1400 6240
rect 1340 6140 1400 6200
rect 1340 6100 1350 6140
rect 1390 6100 1400 6140
rect 1340 6040 1400 6100
rect 1340 6000 1350 6040
rect 1390 6000 1400 6040
rect 1340 5940 1400 6000
rect 1340 5900 1350 5940
rect 1390 5900 1400 5940
rect 1340 5840 1400 5900
rect 1340 5800 1350 5840
rect 1390 5800 1400 5840
rect 1340 5740 1400 5800
rect 1340 5700 1350 5740
rect 1390 5700 1400 5740
rect 1340 5680 1400 5700
rect 1520 6240 1580 6260
rect 1520 6200 1530 6240
rect 1570 6200 1580 6240
rect 1520 6140 1580 6200
rect 1520 6100 1530 6140
rect 1570 6100 1580 6140
rect 1520 6040 1580 6100
rect 1520 6000 1530 6040
rect 1570 6000 1580 6040
rect 1520 5940 1580 6000
rect 1520 5900 1530 5940
rect 1570 5900 1580 5940
rect 1520 5840 1580 5900
rect 1520 5800 1530 5840
rect 1570 5800 1580 5840
rect 1520 5740 1580 5800
rect 1520 5700 1530 5740
rect 1570 5700 1580 5740
rect 1520 5680 1580 5700
rect 1700 6240 1760 6260
rect 1700 6200 1710 6240
rect 1750 6200 1760 6240
rect 1700 6140 1760 6200
rect 1700 6100 1710 6140
rect 1750 6100 1760 6140
rect 1700 6040 1760 6100
rect 1700 6000 1710 6040
rect 1750 6000 1760 6040
rect 1700 5940 1760 6000
rect 1700 5900 1710 5940
rect 1750 5900 1760 5940
rect 1700 5840 1760 5900
rect 1700 5800 1710 5840
rect 1750 5800 1760 5840
rect 1700 5740 1760 5800
rect 1700 5700 1710 5740
rect 1750 5700 1760 5740
rect 1700 5680 1760 5700
rect 1880 6240 2020 6260
rect 1880 6200 1890 6240
rect 1930 6200 1970 6240
rect 2010 6200 2020 6240
rect 1880 6140 2020 6200
rect 1880 6100 1890 6140
rect 1930 6100 1970 6140
rect 2010 6100 2020 6140
rect 2500 6160 2580 6180
rect 2500 6120 2520 6160
rect 2560 6120 2580 6160
rect 2500 6100 2580 6120
rect 2720 6160 2800 6180
rect 2720 6120 2740 6160
rect 2780 6120 2800 6160
rect 2720 6100 2800 6120
rect 2950 6160 3010 6180
rect 6700 6170 6790 6290
rect 2950 6120 2960 6160
rect 3000 6120 3010 6160
rect 2950 6100 3010 6120
rect 6310 6150 6790 6170
rect 6310 6110 6330 6150
rect 6370 6110 6730 6150
rect 6770 6110 6790 6150
rect 1880 6040 2020 6100
rect 6310 6090 6790 6110
rect 1880 6000 1890 6040
rect 1930 6000 1970 6040
rect 2010 6000 2020 6040
rect 1880 5940 2020 6000
rect 1880 5900 1890 5940
rect 1930 5900 1970 5940
rect 2010 5900 2020 5940
rect 1880 5840 2020 5900
rect 2420 6040 2570 6060
rect 2420 6000 2430 6040
rect 2470 6000 2520 6040
rect 2560 6000 2570 6040
rect 2420 5940 2570 6000
rect 2420 5900 2430 5940
rect 2470 5900 2520 5940
rect 2560 5900 2570 5940
rect 2420 5880 2570 5900
rect 2620 6040 2680 6060
rect 2620 6000 2630 6040
rect 2670 6000 2680 6040
rect 2620 5940 2680 6000
rect 2620 5900 2630 5940
rect 2670 5900 2680 5940
rect 2620 5880 2680 5900
rect 2730 6040 2790 6060
rect 2730 6000 2740 6040
rect 2780 6000 2790 6040
rect 2730 5940 2790 6000
rect 2730 5900 2740 5940
rect 2780 5900 2790 5940
rect 2730 5880 2790 5900
rect 2840 6040 2900 6060
rect 2840 6000 2850 6040
rect 2890 6000 2900 6040
rect 2840 5940 2900 6000
rect 2840 5900 2850 5940
rect 2890 5900 2900 5940
rect 2840 5880 2900 5900
rect 2950 6040 3090 6060
rect 6330 6050 6370 6090
rect 6730 6050 6770 6090
rect 2950 6000 2960 6040
rect 3000 6000 3040 6040
rect 3080 6000 3090 6040
rect 2950 5940 3090 6000
rect 2950 5900 2960 5940
rect 3000 5900 3040 5940
rect 3080 5900 3090 5940
rect 2950 5880 3090 5900
rect 5410 6030 5590 6050
rect 5410 5980 5430 6030
rect 5470 5980 5530 6030
rect 5570 5980 5590 6030
rect 5410 5890 5590 5980
rect 5410 5840 5430 5890
rect 5470 5840 5530 5890
rect 5570 5840 5590 5890
rect 1880 5800 1890 5840
rect 1930 5800 1970 5840
rect 2010 5800 2020 5840
rect 1880 5740 2020 5800
rect 2600 5820 2680 5840
rect 2600 5780 2620 5820
rect 2660 5780 2680 5820
rect 2600 5760 2680 5780
rect 2720 5820 2800 5840
rect 2720 5780 2740 5820
rect 2780 5780 2800 5820
rect 2720 5760 2800 5780
rect 2840 5820 2920 5840
rect 5410 5820 5590 5840
rect 5710 6030 5790 6050
rect 5710 5980 5730 6030
rect 5770 5980 5790 6030
rect 5710 5890 5790 5980
rect 5710 5840 5730 5890
rect 5770 5840 5790 5890
rect 5710 5820 5790 5840
rect 5910 6030 5990 6050
rect 5910 5980 5930 6030
rect 5970 5980 5990 6030
rect 5910 5890 5990 5980
rect 5910 5840 5930 5890
rect 5970 5840 5990 5890
rect 5910 5820 5990 5840
rect 6110 6030 6190 6050
rect 6110 5980 6130 6030
rect 6170 5980 6190 6030
rect 6110 5890 6190 5980
rect 6110 5840 6130 5890
rect 6170 5840 6190 5890
rect 6110 5820 6190 5840
rect 6310 6030 6390 6050
rect 6310 5980 6330 6030
rect 6370 5980 6390 6030
rect 6310 5890 6390 5980
rect 6310 5840 6330 5890
rect 6370 5840 6390 5890
rect 6310 5820 6390 5840
rect 6510 6030 6590 6050
rect 6510 5980 6530 6030
rect 6570 5980 6590 6030
rect 6510 5890 6590 5980
rect 6510 5840 6530 5890
rect 6570 5840 6590 5890
rect 6510 5820 6590 5840
rect 6710 6030 6790 6050
rect 6710 5980 6730 6030
rect 6770 5980 6790 6030
rect 6710 5890 6790 5980
rect 6710 5840 6730 5890
rect 6770 5840 6790 5890
rect 6710 5820 6790 5840
rect 6910 6030 6990 6050
rect 6910 5980 6930 6030
rect 6970 5980 6990 6030
rect 6910 5890 6990 5980
rect 6910 5840 6930 5890
rect 6970 5840 6990 5890
rect 6910 5820 6990 5840
rect 7110 6030 7190 6050
rect 7110 5980 7130 6030
rect 7170 5980 7190 6030
rect 7110 5890 7190 5980
rect 7110 5840 7130 5890
rect 7170 5840 7190 5890
rect 7110 5820 7190 5840
rect 7310 6030 7390 6050
rect 7310 5980 7330 6030
rect 7370 5980 7390 6030
rect 7310 5890 7390 5980
rect 7310 5840 7330 5890
rect 7370 5840 7390 5890
rect 7310 5820 7390 5840
rect 7510 6030 7690 6050
rect 7510 5980 7530 6030
rect 7570 5980 7630 6030
rect 7670 5980 7690 6030
rect 7510 5890 7690 5980
rect 7510 5840 7530 5890
rect 7570 5840 7630 5890
rect 7670 5840 7690 5890
rect 7510 5820 7690 5840
rect 2840 5780 2860 5820
rect 2900 5780 2920 5820
rect 5530 5780 5570 5820
rect 5930 5780 5970 5820
rect 7130 5780 7170 5820
rect 7530 5780 7570 5820
rect 2840 5760 2920 5780
rect 5510 5760 5590 5780
rect 1880 5700 1890 5740
rect 1930 5700 1970 5740
rect 2010 5700 2020 5740
rect 5510 5720 5530 5760
rect 5570 5720 5590 5760
rect 5930 5740 7170 5780
rect 5510 5700 5590 5720
rect 7090 5720 7170 5740
rect 1880 5680 2020 5700
rect 7090 5680 7110 5720
rect 7150 5680 7170 5720
rect 7510 5760 7590 5780
rect 7510 5720 7530 5760
rect 7570 5720 7590 5760
rect 7510 5700 7590 5720
rect 7090 5660 7170 5680
rect -1090 5620 -1020 5640
rect -1090 5580 -1080 5620
rect -1040 5580 -1020 5620
rect -1090 5560 -1020 5580
rect -920 5620 -840 5640
rect -920 5580 -900 5620
rect -860 5580 -840 5620
rect -920 5560 -840 5580
rect -740 5620 -660 5640
rect -740 5580 -720 5620
rect -680 5580 -660 5620
rect -740 5560 -660 5580
rect -560 5620 -480 5640
rect -560 5580 -540 5620
rect -500 5580 -480 5620
rect -560 5560 -480 5580
rect -380 5620 -300 5640
rect -380 5580 -360 5620
rect -320 5580 -300 5620
rect -380 5560 -300 5580
rect -200 5620 -120 5640
rect -200 5580 -180 5620
rect -140 5580 -120 5620
rect -200 5560 -120 5580
rect -20 5620 60 5640
rect -20 5580 0 5620
rect 40 5580 60 5620
rect -20 5560 60 5580
rect 160 5620 230 5640
rect 160 5580 180 5620
rect 220 5580 230 5620
rect 160 5560 230 5580
rect 350 5620 420 5640
rect 350 5580 360 5620
rect 400 5580 420 5620
rect 350 5560 420 5580
rect 520 5620 600 5640
rect 520 5580 540 5620
rect 580 5580 600 5620
rect 520 5560 600 5580
rect 700 5620 780 5640
rect 700 5580 720 5620
rect 760 5580 780 5620
rect 700 5560 780 5580
rect 880 5620 960 5640
rect 880 5580 900 5620
rect 940 5580 960 5620
rect 880 5560 960 5580
rect 1060 5620 1140 5640
rect 1060 5580 1080 5620
rect 1120 5580 1140 5620
rect 1060 5560 1140 5580
rect 1240 5620 1320 5640
rect 1240 5580 1260 5620
rect 1300 5580 1320 5620
rect 1240 5560 1320 5580
rect 1420 5620 1500 5640
rect 1420 5580 1440 5620
rect 1480 5580 1500 5620
rect 1420 5560 1500 5580
rect 1600 5620 1670 5640
rect 1600 5580 1620 5620
rect 1660 5580 1670 5620
rect 1600 5560 1670 5580
rect 5950 5610 6030 5630
rect 5950 5570 5970 5610
rect 6010 5570 6030 5610
rect 5950 5550 6030 5570
rect 8230 5610 8310 5630
rect 8230 5570 8250 5610
rect 8290 5570 8310 5610
rect 8230 5550 8310 5570
rect 5620 5470 5710 5490
rect 5620 5440 5640 5470
rect 5580 5420 5640 5440
rect 5690 5440 5710 5470
rect 5970 5440 6010 5550
rect 7090 5500 7170 5520
rect 6270 5470 6360 5490
rect 6270 5440 6290 5470
rect 5690 5420 6290 5440
rect 6340 5440 6360 5470
rect 6760 5460 6840 5480
rect 6760 5440 6780 5460
rect 6340 5420 6400 5440
rect 5580 5400 6400 5420
rect 5580 5360 5620 5400
rect 5710 5360 5750 5400
rect 5970 5360 6010 5400
rect 6230 5360 6270 5400
rect 6360 5360 6400 5400
rect 6720 5420 6780 5440
rect 6820 5440 6840 5460
rect 7090 5460 7110 5500
rect 7150 5460 7170 5500
rect 7090 5440 7170 5460
rect 7420 5460 7500 5480
rect 7420 5440 7440 5460
rect 6820 5420 7440 5440
rect 7480 5440 7500 5460
rect 7900 5460 7980 5480
rect 7900 5450 7920 5460
rect 7480 5420 7540 5440
rect 6720 5400 7540 5420
rect 6720 5360 6760 5400
rect 6850 5360 6890 5400
rect 7110 5360 7150 5400
rect 7370 5360 7410 5400
rect 7500 5360 7540 5400
rect 7860 5420 7920 5450
rect 7960 5450 7980 5460
rect 8250 5450 8290 5550
rect 8560 5460 8640 5480
rect 8560 5450 8580 5460
rect 7960 5420 8580 5450
rect 8620 5450 8640 5460
rect 8620 5420 8680 5450
rect 7860 5400 8680 5420
rect 7860 5360 7900 5400
rect 7990 5360 8030 5400
rect 8250 5360 8290 5400
rect 8510 5360 8550 5400
rect 8640 5360 8680 5400
rect 5460 5340 5640 5360
rect 5460 5300 5480 5340
rect 5520 5300 5580 5340
rect 5620 5300 5640 5340
rect 5460 5280 5640 5300
rect 5690 5340 5770 5360
rect 5690 5300 5710 5340
rect 5750 5300 5770 5340
rect 5690 5280 5770 5300
rect 5820 5340 5900 5360
rect 5820 5300 5840 5340
rect 5880 5300 5900 5340
rect 5820 5280 5900 5300
rect 5950 5340 6030 5360
rect 5950 5300 5970 5340
rect 6010 5300 6030 5340
rect 5950 5280 6030 5300
rect 6080 5340 6160 5360
rect 6080 5300 6100 5340
rect 6140 5300 6160 5340
rect 6080 5280 6160 5300
rect 6210 5340 6290 5360
rect 6210 5300 6230 5340
rect 6270 5300 6290 5340
rect 6210 5280 6290 5300
rect 6340 5340 6520 5360
rect 6340 5300 6360 5340
rect 6400 5300 6460 5340
rect 6500 5300 6520 5340
rect 6340 5280 6520 5300
rect 6700 5340 6780 5360
rect 6700 5300 6720 5340
rect 6760 5300 6780 5340
rect 6700 5280 6780 5300
rect 6830 5340 6910 5360
rect 6830 5300 6850 5340
rect 6890 5300 6910 5340
rect 6830 5280 6910 5300
rect 6960 5340 7040 5360
rect 6960 5300 6980 5340
rect 7020 5300 7040 5340
rect 6960 5280 7040 5300
rect 7090 5340 7170 5360
rect 7090 5300 7110 5340
rect 7150 5300 7170 5340
rect 7090 5280 7170 5300
rect 7220 5340 7300 5360
rect 7220 5300 7240 5340
rect 7280 5300 7300 5340
rect 7220 5280 7300 5300
rect 7350 5340 7430 5360
rect 7350 5300 7370 5340
rect 7410 5300 7430 5340
rect 7350 5280 7430 5300
rect 7480 5340 7560 5360
rect 7480 5300 7500 5340
rect 7540 5300 7560 5340
rect 7480 5280 7560 5300
rect 7740 5340 7920 5360
rect 7740 5300 7760 5340
rect 7800 5300 7860 5340
rect 7900 5300 7920 5340
rect 7740 5280 7920 5300
rect 7970 5340 8050 5360
rect 7970 5300 7990 5340
rect 8030 5300 8050 5340
rect 7970 5280 8050 5300
rect 8100 5340 8180 5360
rect 8100 5300 8120 5340
rect 8160 5300 8180 5340
rect 8100 5280 8180 5300
rect 8230 5340 8310 5360
rect 8230 5300 8250 5340
rect 8290 5300 8310 5340
rect 8230 5280 8310 5300
rect 8360 5340 8440 5360
rect 8360 5300 8380 5340
rect 8420 5300 8440 5340
rect 8360 5280 8440 5300
rect 8490 5340 8570 5360
rect 8490 5300 8510 5340
rect 8550 5300 8570 5340
rect 8490 5280 8570 5300
rect 8620 5340 8800 5360
rect 8620 5300 8640 5340
rect 8680 5300 8740 5340
rect 8780 5300 8800 5340
rect 8620 5280 8800 5300
rect 9550 5330 9660 5350
rect 5820 5220 5900 5240
rect 5820 5180 5840 5220
rect 5880 5180 5900 5220
rect 5820 5160 5900 5180
rect 6870 5220 6950 5240
rect 6870 5180 6890 5220
rect 6930 5180 6950 5220
rect 6870 5160 6950 5180
rect 7310 5220 7390 5240
rect 7310 5180 7330 5220
rect 7370 5180 7390 5220
rect 7310 5160 7390 5180
rect 8140 5120 8180 5280
rect 8360 5120 8400 5280
rect 9550 5260 9570 5330
rect 9640 5260 9660 5330
rect 9550 5240 9660 5260
rect 8850 5220 8930 5240
rect 8850 5180 8870 5220
rect 8910 5180 8930 5220
rect 8850 5160 8930 5180
rect 9550 5120 9590 5240
rect 8010 5100 8090 5120
rect 8010 5060 8030 5100
rect 8070 5060 8090 5100
rect 8140 5080 9760 5120
rect 8010 5040 8090 5060
rect 9720 5070 9760 5080
rect 9720 5050 9800 5070
rect 9720 5010 9740 5050
rect 9780 5010 9800 5050
rect 9720 4990 9800 5010
rect 9720 4980 9760 4990
rect 8140 4940 9760 4980
rect 5730 4880 5810 4900
rect 5730 4840 5750 4880
rect 5790 4840 5810 4880
rect 5730 4820 5810 4840
rect 6170 4880 6250 4900
rect 6170 4840 6190 4880
rect 6230 4840 6250 4880
rect 6170 4820 6250 4840
rect 6960 4890 7040 4910
rect 6960 4850 6980 4890
rect 7020 4850 7040 4890
rect 6960 4830 7040 4850
rect 8010 4880 8090 4900
rect 8010 4840 8030 4880
rect 8070 4840 8090 4880
rect 8010 4820 8090 4840
rect -2460 4800 -2400 4820
rect -2460 4760 -2450 4800
rect -2410 4760 -2400 4800
rect -2460 4740 -2400 4760
rect -60 4800 0 4820
rect -60 4760 -50 4800
rect -10 4760 0 4800
rect -60 4740 0 4760
rect 580 4800 640 4820
rect 580 4760 590 4800
rect 630 4760 640 4800
rect 580 4740 640 4760
rect 2980 4800 3040 4820
rect 2980 4760 2990 4800
rect 3030 4760 3040 4800
rect 8140 4780 8180 4940
rect 8360 4780 8400 4940
rect 8850 4880 8930 4900
rect 8850 4840 8870 4880
rect 8910 4840 8930 4880
rect 8850 4820 8930 4840
rect 9550 4840 9590 4940
rect 9550 4820 9660 4840
rect 2980 4740 3040 4760
rect 5560 4760 5640 4780
rect 5560 4720 5580 4760
rect 5620 4720 5640 4760
rect -2540 4680 -2400 4700
rect -2540 4640 -2530 4680
rect -2490 4640 -2450 4680
rect -2410 4640 -2400 4680
rect -2540 4580 -2400 4640
rect -2540 4540 -2530 4580
rect -2490 4540 -2450 4580
rect -2410 4540 -2400 4580
rect -2540 4520 -2400 4540
rect -2340 4680 -2280 4700
rect -2340 4640 -2330 4680
rect -2290 4640 -2280 4680
rect -2340 4580 -2280 4640
rect -2340 4540 -2330 4580
rect -2290 4540 -2280 4580
rect -2340 4520 -2280 4540
rect -2220 4680 -2160 4700
rect -2220 4640 -2210 4680
rect -2170 4640 -2160 4680
rect -2220 4580 -2160 4640
rect -2220 4540 -2210 4580
rect -2170 4540 -2160 4580
rect -2220 4520 -2160 4540
rect -2100 4680 -2040 4700
rect -2100 4640 -2090 4680
rect -2050 4640 -2040 4680
rect -2100 4580 -2040 4640
rect -2100 4540 -2090 4580
rect -2050 4540 -2040 4580
rect -2100 4520 -2040 4540
rect -1980 4680 -1920 4700
rect -1980 4640 -1970 4680
rect -1930 4640 -1920 4680
rect -1980 4580 -1920 4640
rect -1980 4540 -1970 4580
rect -1930 4540 -1920 4580
rect -1980 4520 -1920 4540
rect -1860 4680 -1800 4700
rect -1860 4640 -1850 4680
rect -1810 4640 -1800 4680
rect -1860 4580 -1800 4640
rect -1860 4540 -1850 4580
rect -1810 4540 -1800 4580
rect -1860 4520 -1800 4540
rect -1740 4680 -1680 4700
rect -1740 4640 -1730 4680
rect -1690 4640 -1680 4680
rect -1740 4580 -1680 4640
rect -1740 4540 -1730 4580
rect -1690 4540 -1680 4580
rect -1740 4520 -1680 4540
rect -1620 4680 -1560 4700
rect -1620 4640 -1610 4680
rect -1570 4640 -1560 4680
rect -1620 4580 -1560 4640
rect -1620 4540 -1610 4580
rect -1570 4540 -1560 4580
rect -1620 4520 -1560 4540
rect -1500 4680 -1440 4700
rect -1500 4640 -1490 4680
rect -1450 4640 -1440 4680
rect -1500 4580 -1440 4640
rect -1500 4540 -1490 4580
rect -1450 4540 -1440 4580
rect -1500 4520 -1440 4540
rect -1380 4680 -1320 4700
rect -1380 4640 -1370 4680
rect -1330 4640 -1320 4680
rect -1380 4580 -1320 4640
rect -1380 4540 -1370 4580
rect -1330 4540 -1320 4580
rect -1380 4520 -1320 4540
rect -1260 4680 -1200 4700
rect -1260 4640 -1250 4680
rect -1210 4640 -1200 4680
rect -1260 4580 -1200 4640
rect -1260 4540 -1250 4580
rect -1210 4540 -1200 4580
rect -1260 4520 -1200 4540
rect -1140 4680 -1080 4700
rect -1140 4640 -1130 4680
rect -1090 4640 -1080 4680
rect -1140 4580 -1080 4640
rect -1140 4540 -1130 4580
rect -1090 4540 -1080 4580
rect -1140 4520 -1080 4540
rect -1020 4680 -960 4700
rect -1020 4640 -1010 4680
rect -970 4640 -960 4680
rect -1020 4580 -960 4640
rect -1020 4540 -1010 4580
rect -970 4540 -960 4580
rect -1020 4520 -960 4540
rect -900 4680 -840 4700
rect -900 4640 -890 4680
rect -850 4640 -840 4680
rect -900 4580 -840 4640
rect -900 4540 -890 4580
rect -850 4540 -840 4580
rect -900 4520 -840 4540
rect -780 4680 -720 4700
rect -780 4640 -770 4680
rect -730 4640 -720 4680
rect -780 4580 -720 4640
rect -780 4540 -770 4580
rect -730 4540 -720 4580
rect -780 4520 -720 4540
rect -660 4680 -600 4700
rect -660 4640 -650 4680
rect -610 4640 -600 4680
rect -660 4580 -600 4640
rect -660 4540 -650 4580
rect -610 4540 -600 4580
rect -660 4520 -600 4540
rect -540 4680 -480 4700
rect -540 4640 -530 4680
rect -490 4640 -480 4680
rect -540 4580 -480 4640
rect -540 4540 -530 4580
rect -490 4540 -480 4580
rect -540 4520 -480 4540
rect -420 4680 -360 4700
rect -420 4640 -410 4680
rect -370 4640 -360 4680
rect -420 4580 -360 4640
rect -420 4540 -410 4580
rect -370 4540 -360 4580
rect -420 4520 -360 4540
rect -300 4680 -240 4700
rect -300 4640 -290 4680
rect -250 4640 -240 4680
rect -300 4580 -240 4640
rect -300 4540 -290 4580
rect -250 4540 -240 4580
rect -300 4520 -240 4540
rect -180 4680 -120 4700
rect -180 4640 -170 4680
rect -130 4640 -120 4680
rect -180 4580 -120 4640
rect -180 4540 -170 4580
rect -130 4540 -120 4580
rect -180 4520 -120 4540
rect -60 4680 80 4700
rect -60 4640 -50 4680
rect -10 4640 30 4680
rect 70 4640 80 4680
rect -60 4580 80 4640
rect -60 4540 -50 4580
rect -10 4540 30 4580
rect 70 4540 80 4580
rect -60 4520 80 4540
rect 500 4680 640 4700
rect 500 4640 510 4680
rect 550 4640 590 4680
rect 630 4640 640 4680
rect 500 4580 640 4640
rect 500 4540 510 4580
rect 550 4540 590 4580
rect 630 4540 640 4580
rect 500 4520 640 4540
rect 700 4680 760 4700
rect 700 4640 710 4680
rect 750 4640 760 4680
rect 700 4580 760 4640
rect 700 4540 710 4580
rect 750 4540 760 4580
rect 700 4520 760 4540
rect 820 4680 880 4700
rect 820 4640 830 4680
rect 870 4640 880 4680
rect 820 4580 880 4640
rect 820 4540 830 4580
rect 870 4540 880 4580
rect 820 4520 880 4540
rect 940 4680 1000 4700
rect 940 4640 950 4680
rect 990 4640 1000 4680
rect 940 4580 1000 4640
rect 940 4540 950 4580
rect 990 4540 1000 4580
rect 940 4520 1000 4540
rect 1060 4680 1120 4700
rect 1060 4640 1070 4680
rect 1110 4640 1120 4680
rect 1060 4580 1120 4640
rect 1060 4540 1070 4580
rect 1110 4540 1120 4580
rect 1060 4520 1120 4540
rect 1180 4680 1240 4700
rect 1180 4640 1190 4680
rect 1230 4640 1240 4680
rect 1180 4580 1240 4640
rect 1180 4540 1190 4580
rect 1230 4540 1240 4580
rect 1180 4520 1240 4540
rect 1300 4680 1360 4700
rect 1300 4640 1310 4680
rect 1350 4640 1360 4680
rect 1300 4580 1360 4640
rect 1300 4540 1310 4580
rect 1350 4540 1360 4580
rect 1300 4520 1360 4540
rect 1420 4680 1480 4700
rect 1420 4640 1430 4680
rect 1470 4640 1480 4680
rect 1420 4580 1480 4640
rect 1420 4540 1430 4580
rect 1470 4540 1480 4580
rect 1420 4520 1480 4540
rect 1540 4680 1600 4700
rect 1540 4640 1550 4680
rect 1590 4640 1600 4680
rect 1540 4580 1600 4640
rect 1540 4540 1550 4580
rect 1590 4540 1600 4580
rect 1540 4520 1600 4540
rect 1660 4680 1720 4700
rect 1660 4640 1670 4680
rect 1710 4640 1720 4680
rect 1660 4580 1720 4640
rect 1660 4540 1670 4580
rect 1710 4540 1720 4580
rect 1660 4520 1720 4540
rect 1780 4680 1840 4700
rect 1780 4640 1790 4680
rect 1830 4640 1840 4680
rect 1780 4580 1840 4640
rect 1780 4540 1790 4580
rect 1830 4540 1840 4580
rect 1780 4520 1840 4540
rect 1900 4680 1960 4700
rect 1900 4640 1910 4680
rect 1950 4640 1960 4680
rect 1900 4580 1960 4640
rect 1900 4540 1910 4580
rect 1950 4540 1960 4580
rect 1900 4520 1960 4540
rect 2020 4680 2080 4700
rect 2020 4640 2030 4680
rect 2070 4640 2080 4680
rect 2020 4580 2080 4640
rect 2020 4540 2030 4580
rect 2070 4540 2080 4580
rect 2020 4520 2080 4540
rect 2140 4680 2200 4700
rect 2140 4640 2150 4680
rect 2190 4640 2200 4680
rect 2140 4580 2200 4640
rect 2140 4540 2150 4580
rect 2190 4540 2200 4580
rect 2140 4520 2200 4540
rect 2260 4680 2320 4700
rect 2260 4640 2270 4680
rect 2310 4640 2320 4680
rect 2260 4580 2320 4640
rect 2260 4540 2270 4580
rect 2310 4540 2320 4580
rect 2260 4520 2320 4540
rect 2380 4680 2440 4700
rect 2380 4640 2390 4680
rect 2430 4640 2440 4680
rect 2380 4580 2440 4640
rect 2380 4540 2390 4580
rect 2430 4540 2440 4580
rect 2380 4520 2440 4540
rect 2500 4680 2560 4700
rect 2500 4640 2510 4680
rect 2550 4640 2560 4680
rect 2500 4580 2560 4640
rect 2500 4540 2510 4580
rect 2550 4540 2560 4580
rect 2500 4520 2560 4540
rect 2620 4680 2680 4700
rect 2620 4640 2630 4680
rect 2670 4640 2680 4680
rect 2620 4580 2680 4640
rect 2620 4540 2630 4580
rect 2670 4540 2680 4580
rect 2620 4520 2680 4540
rect 2740 4680 2800 4700
rect 2740 4640 2750 4680
rect 2790 4640 2800 4680
rect 2740 4580 2800 4640
rect 2740 4540 2750 4580
rect 2790 4540 2800 4580
rect 2740 4520 2800 4540
rect 2860 4680 2920 4700
rect 2860 4640 2870 4680
rect 2910 4640 2920 4680
rect 2860 4580 2920 4640
rect 2860 4540 2870 4580
rect 2910 4540 2920 4580
rect 2860 4520 2920 4540
rect 2980 4680 3120 4700
rect 2980 4640 2990 4680
rect 3030 4640 3070 4680
rect 3110 4640 3120 4680
rect 2980 4580 3120 4640
rect 5560 4660 5640 4720
rect 5560 4620 5580 4660
rect 5620 4620 5640 4660
rect 5560 4600 5640 4620
rect 5690 4760 5770 4780
rect 5690 4720 5710 4760
rect 5750 4720 5770 4760
rect 5690 4660 5770 4720
rect 5690 4620 5710 4660
rect 5750 4620 5770 4660
rect 5690 4600 5770 4620
rect 5820 4760 5900 4780
rect 5820 4720 5840 4760
rect 5880 4720 5900 4760
rect 5820 4660 5900 4720
rect 5820 4620 5840 4660
rect 5880 4620 5900 4660
rect 5820 4600 5900 4620
rect 5950 4760 6030 4780
rect 5950 4720 5970 4760
rect 6010 4720 6030 4760
rect 5950 4660 6030 4720
rect 5950 4620 5970 4660
rect 6010 4620 6030 4660
rect 5950 4600 6030 4620
rect 6080 4760 6160 4780
rect 6080 4720 6100 4760
rect 6140 4720 6160 4760
rect 6080 4660 6160 4720
rect 6080 4620 6100 4660
rect 6140 4620 6160 4660
rect 6080 4600 6160 4620
rect 6210 4760 6300 4780
rect 6210 4720 6230 4760
rect 6270 4720 6300 4760
rect 6210 4660 6300 4720
rect 6210 4620 6230 4660
rect 6270 4620 6300 4660
rect 6210 4600 6300 4620
rect 6340 4760 6420 4780
rect 6340 4720 6360 4760
rect 6400 4720 6420 4760
rect 6340 4660 6420 4720
rect 6340 4620 6360 4660
rect 6400 4620 6420 4660
rect 6340 4600 6420 4620
rect 6600 4760 6780 4780
rect 6600 4720 6620 4760
rect 6660 4720 6720 4760
rect 6760 4720 6780 4760
rect 6600 4660 6780 4720
rect 6600 4620 6620 4660
rect 6660 4620 6720 4660
rect 6760 4620 6780 4660
rect 6600 4600 6780 4620
rect 6830 4760 6910 4780
rect 6830 4720 6850 4760
rect 6890 4720 6910 4760
rect 6830 4660 6910 4720
rect 6830 4620 6850 4660
rect 6890 4620 6910 4660
rect 6830 4600 6910 4620
rect 6960 4760 7040 4780
rect 6960 4720 6980 4760
rect 7020 4720 7040 4760
rect 6960 4660 7040 4720
rect 6960 4620 6980 4660
rect 7020 4620 7040 4660
rect 6960 4600 7040 4620
rect 7090 4760 7170 4780
rect 7090 4720 7110 4760
rect 7150 4720 7170 4760
rect 7090 4660 7170 4720
rect 7090 4620 7110 4660
rect 7150 4620 7170 4660
rect 7090 4600 7170 4620
rect 7220 4760 7300 4780
rect 7220 4720 7240 4760
rect 7280 4720 7300 4760
rect 7220 4660 7300 4720
rect 7220 4620 7240 4660
rect 7280 4620 7300 4660
rect 7220 4600 7300 4620
rect 7350 4760 7430 4780
rect 7350 4720 7370 4760
rect 7410 4720 7430 4760
rect 7350 4660 7430 4720
rect 7350 4620 7370 4660
rect 7410 4620 7430 4660
rect 7350 4600 7430 4620
rect 7480 4760 7660 4780
rect 7480 4720 7500 4760
rect 7540 4720 7600 4760
rect 7640 4720 7660 4760
rect 7480 4660 7660 4720
rect 7480 4620 7500 4660
rect 7540 4620 7600 4660
rect 7640 4620 7660 4660
rect 7480 4600 7660 4620
rect 7740 4760 7920 4780
rect 7740 4720 7760 4760
rect 7800 4720 7860 4760
rect 7900 4720 7920 4760
rect 7740 4660 7920 4720
rect 7740 4620 7760 4660
rect 7800 4620 7860 4660
rect 7900 4620 7920 4660
rect 7740 4600 7920 4620
rect 7970 4760 8050 4780
rect 7970 4720 7990 4760
rect 8030 4720 8050 4760
rect 7970 4660 8050 4720
rect 7970 4620 7990 4660
rect 8030 4620 8050 4660
rect 7970 4600 8050 4620
rect 8100 4760 8180 4780
rect 8100 4720 8120 4760
rect 8160 4720 8180 4760
rect 8100 4660 8180 4720
rect 8100 4620 8120 4660
rect 8160 4620 8180 4660
rect 8100 4600 8180 4620
rect 8230 4760 8310 4780
rect 8230 4720 8250 4760
rect 8290 4720 8310 4760
rect 8230 4660 8310 4720
rect 8230 4620 8250 4660
rect 8290 4620 8310 4660
rect 8230 4600 8310 4620
rect 8360 4760 8440 4780
rect 8360 4720 8380 4760
rect 8420 4720 8440 4760
rect 8360 4660 8440 4720
rect 8360 4620 8380 4660
rect 8420 4620 8440 4660
rect 8360 4600 8440 4620
rect 8490 4760 8570 4780
rect 8490 4720 8510 4760
rect 8550 4720 8570 4760
rect 8490 4660 8570 4720
rect 8490 4620 8510 4660
rect 8550 4620 8570 4660
rect 8490 4600 8570 4620
rect 8620 4760 8800 4780
rect 8620 4720 8640 4760
rect 8680 4720 8740 4760
rect 8780 4720 8800 4760
rect 9550 4750 9570 4820
rect 9640 4750 9660 4820
rect 9550 4730 9660 4750
rect 8620 4660 8800 4720
rect 8620 4620 8640 4660
rect 8680 4620 8740 4660
rect 8780 4620 8800 4660
rect 8620 4600 8800 4620
rect 2980 4540 2990 4580
rect 3030 4540 3070 4580
rect 3110 4540 3120 4580
rect 2980 4520 3120 4540
rect 5580 4560 5620 4600
rect 5710 4560 5750 4600
rect 5970 4560 6010 4600
rect 6230 4560 6270 4600
rect 6360 4560 6400 4600
rect 5580 4540 6400 4560
rect 5580 4520 5640 4540
rect 5620 4500 5640 4520
rect 5680 4520 6300 4540
rect 5680 4500 5700 4520
rect 5620 4480 5700 4500
rect 6030 4500 6110 4520
rect -2280 4450 -2220 4470
rect -2280 4410 -2270 4450
rect -2230 4410 -2220 4450
rect -2280 4390 -2220 4410
rect -2110 4460 -2030 4480
rect -2110 4420 -2090 4460
rect -2050 4420 -2030 4460
rect -2110 4400 -2030 4420
rect -1620 4460 -1560 4480
rect -1620 4420 -1610 4460
rect -1570 4420 -1560 4460
rect -1620 4400 -1560 4420
rect -1390 4460 -1310 4480
rect -1390 4420 -1370 4460
rect -1330 4420 -1310 4460
rect -1390 4400 -1310 4420
rect -900 4460 -840 4480
rect -900 4420 -890 4460
rect -850 4420 -840 4460
rect -900 4400 -840 4420
rect -670 4460 -590 4480
rect -670 4420 -650 4460
rect -610 4420 -590 4460
rect -670 4400 -590 4420
rect -240 4460 -180 4480
rect -240 4420 -230 4460
rect -190 4420 -180 4460
rect -240 4400 -180 4420
rect 760 4460 820 4480
rect 760 4420 770 4460
rect 810 4420 820 4460
rect 760 4400 820 4420
rect 1170 4460 1250 4480
rect 1170 4420 1190 4460
rect 1230 4420 1250 4460
rect 1170 4400 1250 4420
rect 1420 4460 1480 4480
rect 1420 4420 1430 4460
rect 1470 4420 1480 4460
rect 1420 4400 1480 4420
rect 1890 4460 1970 4480
rect 1890 4420 1910 4460
rect 1950 4420 1970 4460
rect 1890 4400 1970 4420
rect 2140 4460 2200 4480
rect 2140 4420 2150 4460
rect 2190 4420 2200 4460
rect 2140 4400 2200 4420
rect 2610 4460 2690 4480
rect 2610 4420 2630 4460
rect 2670 4420 2690 4460
rect 2610 4400 2690 4420
rect 2800 4450 2860 4470
rect 2800 4410 2810 4450
rect 2850 4410 2860 4450
rect 6030 4460 6050 4500
rect 6090 4460 6110 4500
rect 6280 4500 6300 4520
rect 6340 4520 6400 4540
rect 6720 4560 6760 4600
rect 6850 4560 6890 4600
rect 7110 4560 7150 4600
rect 7370 4560 7410 4600
rect 7500 4560 7540 4600
rect 6720 4540 7540 4560
rect 6720 4520 6780 4540
rect 6340 4500 6360 4520
rect 6280 4480 6360 4500
rect 6760 4500 6780 4520
rect 6820 4520 7440 4540
rect 6820 4500 6840 4520
rect 6760 4480 6840 4500
rect 6030 4440 6110 4460
rect 2800 4390 2860 4410
rect 7110 4410 7150 4520
rect 7420 4500 7440 4520
rect 7480 4520 7540 4540
rect 7860 4560 7900 4600
rect 7990 4560 8030 4600
rect 8250 4560 8290 4600
rect 8510 4560 8550 4600
rect 8640 4560 8680 4600
rect 7860 4540 8680 4560
rect 7860 4520 7920 4540
rect 7480 4500 7500 4520
rect 7420 4480 7500 4500
rect 7900 4500 7920 4520
rect 7960 4520 8580 4540
rect 7960 4500 7980 4520
rect 7900 4480 7980 4500
rect 8250 4410 8290 4520
rect 8560 4500 8580 4520
rect 8620 4520 8680 4540
rect 8620 4500 8640 4520
rect 8560 4480 8640 4500
rect 7110 4390 7190 4410
rect 7110 4350 7130 4390
rect 7170 4350 7190 4390
rect 7110 4330 7190 4350
rect 8230 4390 8310 4410
rect 8230 4350 8250 4390
rect 8290 4350 8310 4390
rect 8230 4330 8310 4350
rect 5630 4230 5710 4250
rect 5630 4190 5650 4230
rect 5690 4190 5710 4230
rect 5630 4130 5710 4190
rect 7630 4230 7710 4250
rect 7630 4190 7650 4230
rect 7690 4190 7710 4230
rect 7630 4170 7710 4190
rect 5530 4110 5710 4130
rect 5530 4070 5550 4110
rect 5590 4070 5650 4110
rect 5690 4070 5710 4110
rect 5530 4010 5710 4070
rect 5530 3970 5550 4010
rect 5590 3970 5650 4010
rect 5690 3970 5710 4010
rect 5530 3910 5710 3970
rect 5530 3870 5550 3910
rect 5590 3870 5650 3910
rect 5690 3870 5710 3910
rect -1458 3852 -1400 3870
rect -1458 3818 -1446 3852
rect -1412 3818 -1400 3852
rect -1458 3800 -1400 3818
rect -1300 3852 -1242 3870
rect -1300 3818 -1288 3852
rect -1254 3818 -1242 3852
rect -1300 3800 -1242 3818
rect -976 3852 -918 3870
rect -976 3818 -964 3852
rect -930 3818 -918 3852
rect -976 3800 -918 3818
rect -822 3852 -764 3870
rect -822 3818 -810 3852
rect -776 3818 -764 3852
rect -822 3800 -764 3818
rect -498 3852 -440 3870
rect -498 3818 -486 3852
rect -452 3818 -440 3852
rect 1020 3852 1078 3870
rect -498 3800 -440 3818
rect -190 3810 -110 3830
rect -190 3770 -170 3810
rect -130 3770 -110 3810
rect -1620 3740 -1560 3760
rect -1620 3700 -1610 3740
rect -1570 3700 -1560 3740
rect -1620 3680 -1560 3700
rect -1500 3740 -1440 3760
rect -1500 3700 -1490 3740
rect -1450 3700 -1440 3740
rect -1500 3680 -1440 3700
rect -1380 3740 -1320 3760
rect -1380 3700 -1370 3740
rect -1330 3700 -1320 3740
rect -1380 3680 -1320 3700
rect -1260 3740 -1200 3760
rect -1260 3700 -1250 3740
rect -1210 3700 -1200 3740
rect -1260 3680 -1200 3700
rect -1140 3740 -1080 3760
rect -1140 3700 -1130 3740
rect -1090 3700 -1080 3740
rect -1140 3680 -1080 3700
rect -1020 3740 -960 3760
rect -1020 3700 -1010 3740
rect -970 3700 -960 3740
rect -1020 3680 -960 3700
rect -900 3740 -840 3760
rect -900 3700 -890 3740
rect -850 3700 -840 3740
rect -900 3680 -840 3700
rect -780 3740 -720 3760
rect -780 3700 -770 3740
rect -730 3700 -720 3740
rect -780 3680 -720 3700
rect -660 3740 -600 3760
rect -660 3700 -650 3740
rect -610 3700 -600 3740
rect -660 3680 -600 3700
rect -540 3740 -480 3760
rect -540 3700 -530 3740
rect -490 3700 -480 3740
rect -540 3680 -480 3700
rect -420 3740 -360 3760
rect -420 3700 -410 3740
rect -370 3700 -360 3740
rect -420 3680 -360 3700
rect -190 3730 -110 3770
rect -190 3690 -170 3730
rect -130 3690 -110 3730
rect -190 3650 -110 3690
rect -1559 3622 -1501 3640
rect -1559 3588 -1547 3622
rect -1513 3588 -1501 3622
rect -1559 3570 -1501 3588
rect -1199 3622 -1141 3640
rect -1199 3588 -1187 3622
rect -1153 3588 -1141 3622
rect -1199 3570 -1141 3588
rect -1079 3622 -1021 3640
rect -1079 3588 -1067 3622
rect -1033 3588 -1021 3622
rect -1079 3570 -1021 3588
rect -719 3622 -661 3640
rect -719 3588 -707 3622
rect -673 3588 -661 3622
rect -719 3570 -661 3588
rect -599 3622 -541 3640
rect -599 3588 -587 3622
rect -553 3588 -541 3622
rect -190 3610 -170 3650
rect -130 3610 -110 3650
rect -190 3590 -110 3610
rect 690 3810 770 3830
rect 690 3770 710 3810
rect 750 3770 770 3810
rect 1020 3818 1032 3852
rect 1066 3818 1078 3852
rect 1020 3800 1078 3818
rect 1344 3852 1402 3870
rect 1344 3818 1356 3852
rect 1390 3818 1402 3852
rect 1344 3800 1402 3818
rect 1498 3852 1556 3870
rect 1498 3818 1510 3852
rect 1544 3818 1556 3852
rect 1498 3800 1556 3818
rect 1822 3852 1880 3870
rect 1822 3818 1834 3852
rect 1868 3818 1880 3852
rect 1822 3800 1880 3818
rect 1980 3852 2038 3870
rect 1980 3818 1992 3852
rect 2026 3818 2038 3852
rect 1980 3800 2038 3818
rect 5530 3810 5710 3870
rect 690 3730 770 3770
rect 5530 3770 5550 3810
rect 5590 3770 5650 3810
rect 5690 3770 5710 3810
rect 690 3690 710 3730
rect 750 3690 770 3730
rect 690 3650 770 3690
rect 940 3740 1000 3760
rect 940 3700 950 3740
rect 990 3700 1000 3740
rect 940 3680 1000 3700
rect 1060 3740 1120 3760
rect 1060 3700 1070 3740
rect 1110 3700 1120 3740
rect 1060 3680 1120 3700
rect 1180 3740 1240 3760
rect 1180 3700 1190 3740
rect 1230 3700 1240 3740
rect 1180 3680 1240 3700
rect 1300 3740 1360 3760
rect 1300 3700 1310 3740
rect 1350 3700 1360 3740
rect 1300 3680 1360 3700
rect 1420 3740 1480 3760
rect 1420 3700 1430 3740
rect 1470 3700 1480 3740
rect 1420 3680 1480 3700
rect 1540 3740 1600 3760
rect 1540 3700 1550 3740
rect 1590 3700 1600 3740
rect 1540 3680 1600 3700
rect 1660 3740 1720 3760
rect 1660 3700 1670 3740
rect 1710 3700 1720 3740
rect 1660 3680 1720 3700
rect 1780 3740 1840 3760
rect 1780 3700 1790 3740
rect 1830 3700 1840 3740
rect 1780 3680 1840 3700
rect 1900 3740 1960 3760
rect 1900 3700 1910 3740
rect 1950 3700 1960 3740
rect 1900 3680 1960 3700
rect 2020 3740 2080 3760
rect 2020 3700 2030 3740
rect 2070 3700 2080 3740
rect 2020 3680 2080 3700
rect 2140 3740 2200 3760
rect 2140 3700 2150 3740
rect 2190 3700 2200 3740
rect 2140 3680 2200 3700
rect 5530 3710 5710 3770
rect 5530 3670 5550 3710
rect 5590 3670 5650 3710
rect 5690 3670 5710 3710
rect 5530 3650 5710 3670
rect 5830 4110 5910 4130
rect 5830 4070 5850 4110
rect 5890 4070 5910 4110
rect 5830 4010 5910 4070
rect 5830 3970 5850 4010
rect 5890 3970 5910 4010
rect 5830 3910 5910 3970
rect 5830 3870 5850 3910
rect 5890 3870 5910 3910
rect 5830 3810 5910 3870
rect 5830 3770 5850 3810
rect 5890 3770 5910 3810
rect 5830 3710 5910 3770
rect 5830 3670 5850 3710
rect 5890 3670 5910 3710
rect 5830 3650 5910 3670
rect 6030 4110 6110 4130
rect 6030 4070 6050 4110
rect 6090 4070 6110 4110
rect 6030 4010 6110 4070
rect 6030 3970 6050 4010
rect 6090 3970 6110 4010
rect 6030 3910 6110 3970
rect 6030 3870 6050 3910
rect 6090 3870 6110 3910
rect 6030 3810 6110 3870
rect 6030 3770 6050 3810
rect 6090 3770 6110 3810
rect 6030 3710 6110 3770
rect 6030 3670 6050 3710
rect 6090 3670 6110 3710
rect 6030 3650 6110 3670
rect 6230 4110 6310 4130
rect 6230 4070 6250 4110
rect 6290 4070 6310 4110
rect 6230 4010 6310 4070
rect 6230 3970 6250 4010
rect 6290 3970 6310 4010
rect 6230 3910 6310 3970
rect 6230 3870 6250 3910
rect 6290 3870 6310 3910
rect 6230 3810 6310 3870
rect 6230 3770 6250 3810
rect 6290 3770 6310 3810
rect 6230 3710 6310 3770
rect 6230 3670 6250 3710
rect 6290 3670 6310 3710
rect 6230 3650 6310 3670
rect 6430 4110 6510 4130
rect 6430 4070 6450 4110
rect 6490 4070 6510 4110
rect 6430 4010 6510 4070
rect 6430 3970 6450 4010
rect 6490 3970 6510 4010
rect 6430 3910 6510 3970
rect 6430 3870 6450 3910
rect 6490 3870 6510 3910
rect 6430 3810 6510 3870
rect 6430 3770 6450 3810
rect 6490 3770 6510 3810
rect 6430 3710 6510 3770
rect 6430 3670 6450 3710
rect 6490 3670 6510 3710
rect 6430 3650 6510 3670
rect 6630 4110 6710 4130
rect 6630 4070 6650 4110
rect 6690 4070 6710 4110
rect 6630 4010 6710 4070
rect 6630 3970 6650 4010
rect 6690 3970 6710 4010
rect 6630 3910 6710 3970
rect 6630 3870 6650 3910
rect 6690 3870 6710 3910
rect 6630 3810 6710 3870
rect 6630 3770 6650 3810
rect 6690 3770 6710 3810
rect 6630 3710 6710 3770
rect 6630 3670 6650 3710
rect 6690 3670 6710 3710
rect 6630 3650 6710 3670
rect 6830 4110 6910 4130
rect 6830 4070 6850 4110
rect 6890 4070 6910 4110
rect 6830 4010 6910 4070
rect 6830 3970 6850 4010
rect 6890 3970 6910 4010
rect 6830 3910 6910 3970
rect 6830 3870 6850 3910
rect 6890 3870 6910 3910
rect 6830 3810 6910 3870
rect 6830 3770 6850 3810
rect 6890 3770 6910 3810
rect 6830 3710 6910 3770
rect 6830 3670 6850 3710
rect 6890 3670 6910 3710
rect 6830 3650 6910 3670
rect 7030 4110 7110 4130
rect 7030 4070 7050 4110
rect 7090 4070 7110 4110
rect 7030 4010 7110 4070
rect 7030 3970 7050 4010
rect 7090 3970 7110 4010
rect 7030 3910 7110 3970
rect 7030 3870 7050 3910
rect 7090 3870 7110 3910
rect 7030 3810 7110 3870
rect 7030 3770 7050 3810
rect 7090 3770 7110 3810
rect 7030 3710 7110 3770
rect 7030 3670 7050 3710
rect 7090 3670 7110 3710
rect 7030 3650 7110 3670
rect 7230 4110 7310 4130
rect 7230 4070 7250 4110
rect 7290 4070 7310 4110
rect 7230 4010 7310 4070
rect 7230 3970 7250 4010
rect 7290 3970 7310 4010
rect 7230 3910 7310 3970
rect 7230 3870 7250 3910
rect 7290 3870 7310 3910
rect 7230 3810 7310 3870
rect 7230 3770 7250 3810
rect 7290 3770 7310 3810
rect 7230 3710 7310 3770
rect 7230 3670 7250 3710
rect 7290 3670 7310 3710
rect 7230 3650 7310 3670
rect 7430 4110 7510 4130
rect 7430 4070 7450 4110
rect 7490 4070 7510 4110
rect 7430 4010 7510 4070
rect 7430 3970 7450 4010
rect 7490 3970 7510 4010
rect 7430 3910 7510 3970
rect 7430 3870 7450 3910
rect 7490 3870 7510 3910
rect 7430 3810 7510 3870
rect 7430 3770 7450 3810
rect 7490 3770 7510 3810
rect 7430 3710 7510 3770
rect 7430 3670 7450 3710
rect 7490 3670 7510 3710
rect 7430 3650 7510 3670
rect 7630 4110 7810 4130
rect 7630 4070 7650 4110
rect 7690 4070 7750 4110
rect 7790 4070 7810 4110
rect 7630 4010 7810 4070
rect 7630 3970 7650 4010
rect 7690 3970 7750 4010
rect 7790 3970 7810 4010
rect 7630 3910 7810 3970
rect 7630 3870 7650 3910
rect 7690 3870 7750 3910
rect 7790 3870 7810 3910
rect 7630 3810 7810 3870
rect 7630 3770 7650 3810
rect 7690 3770 7750 3810
rect 7790 3770 7810 3810
rect 7630 3710 7810 3770
rect 7630 3670 7650 3710
rect 7690 3670 7750 3710
rect 7790 3670 7810 3710
rect 7630 3650 7810 3670
rect 690 3610 710 3650
rect 750 3610 770 3650
rect 690 3590 770 3610
rect 1121 3622 1179 3640
rect -599 3570 -541 3588
rect 1121 3588 1133 3622
rect 1167 3588 1179 3622
rect 1121 3570 1179 3588
rect 1241 3622 1299 3640
rect 1241 3588 1253 3622
rect 1287 3588 1299 3622
rect 1241 3570 1299 3588
rect 1601 3622 1659 3640
rect 1601 3588 1613 3622
rect 1647 3588 1659 3622
rect 1601 3570 1659 3588
rect 1721 3622 1779 3640
rect 1721 3588 1733 3622
rect 1767 3588 1779 3622
rect 1721 3570 1779 3588
rect 2081 3622 2139 3640
rect 2081 3588 2093 3622
rect 2127 3588 2139 3622
rect 2081 3570 2139 3588
rect 6430 3590 6510 3610
rect 6430 3550 6450 3590
rect 6490 3550 6510 3590
rect 6430 3530 6510 3550
rect 6830 3590 6910 3610
rect 6830 3550 6850 3590
rect 6890 3550 6910 3590
rect 6830 3530 6910 3550
rect -2070 3250 -1990 3270
rect -2250 3210 -2170 3230
rect -2250 3170 -2230 3210
rect -2190 3170 -2170 3210
rect -2070 3210 -2050 3250
rect -2010 3210 -1990 3250
rect -2070 3190 -1990 3210
rect -1830 3250 -1750 3270
rect -1830 3210 -1810 3250
rect -1770 3210 -1750 3250
rect -1830 3190 -1750 3210
rect -1590 3250 -1510 3270
rect -1590 3210 -1570 3250
rect -1530 3210 -1510 3250
rect -1590 3190 -1510 3210
rect -1350 3250 -1270 3270
rect -1350 3210 -1330 3250
rect -1290 3210 -1270 3250
rect -1350 3190 -1270 3210
rect -710 3250 -630 3270
rect -710 3210 -690 3250
rect -650 3210 -630 3250
rect -710 3190 -630 3210
rect -470 3250 -390 3270
rect -470 3210 -450 3250
rect -410 3210 -390 3250
rect -470 3190 -390 3210
rect -230 3250 -150 3270
rect -230 3210 -210 3250
rect -170 3210 -150 3250
rect 730 3250 810 3270
rect -230 3190 -150 3210
rect 80 3220 140 3240
rect -2250 3150 -2170 3170
rect 80 3180 90 3220
rect 130 3180 140 3220
rect -2240 3130 -2180 3150
rect -2240 3090 -2230 3130
rect -2190 3090 -2180 3130
rect -2240 3030 -2180 3090
rect -2240 2990 -2230 3030
rect -2190 2990 -2180 3030
rect -2240 2930 -2180 2990
rect -2240 2890 -2230 2930
rect -2190 2890 -2180 2930
rect -2240 2830 -2180 2890
rect -2240 2790 -2230 2830
rect -2190 2790 -2180 2830
rect -2240 2730 -2180 2790
rect -2240 2690 -2230 2730
rect -2190 2690 -2180 2730
rect -2240 2670 -2180 2690
rect -1160 3130 -940 3150
rect -1160 3090 -1150 3130
rect -1110 3090 -1070 3130
rect -1030 3090 -990 3130
rect -950 3090 -940 3130
rect -1160 3030 -940 3090
rect -1160 2990 -1150 3030
rect -1110 2990 -1070 3030
rect -1030 2990 -990 3030
rect -950 2990 -940 3030
rect -1160 2930 -940 2990
rect -1160 2890 -1150 2930
rect -1110 2890 -1070 2930
rect -1030 2890 -990 2930
rect -950 2890 -940 2930
rect -1160 2830 -940 2890
rect -1160 2790 -1150 2830
rect -1110 2790 -1070 2830
rect -1030 2790 -990 2830
rect -950 2790 -940 2830
rect -1160 2730 -940 2790
rect -1160 2690 -1150 2730
rect -1110 2690 -1070 2730
rect -1030 2690 -990 2730
rect -950 2690 -940 2730
rect -1160 2670 -940 2690
rect 80 3130 140 3180
rect 80 3090 90 3130
rect 130 3090 140 3130
rect 80 3030 140 3090
rect 80 2990 90 3030
rect 130 2990 140 3030
rect 80 2930 140 2990
rect 80 2890 90 2930
rect 130 2890 140 2930
rect 80 2830 140 2890
rect 80 2790 90 2830
rect 130 2790 140 2830
rect 80 2730 140 2790
rect 80 2690 90 2730
rect 130 2690 140 2730
rect 80 2670 140 2690
rect 440 3220 500 3240
rect 440 3180 450 3220
rect 490 3180 500 3220
rect 730 3210 750 3250
rect 790 3210 810 3250
rect 730 3190 810 3210
rect 970 3250 1050 3270
rect 970 3210 990 3250
rect 1030 3210 1050 3250
rect 970 3190 1050 3210
rect 1210 3250 1290 3270
rect 1210 3210 1230 3250
rect 1270 3210 1290 3250
rect 1210 3190 1290 3210
rect 1850 3250 1930 3270
rect 1850 3210 1870 3250
rect 1910 3210 1930 3250
rect 1850 3190 1930 3210
rect 2090 3250 2170 3270
rect 2090 3210 2110 3250
rect 2150 3210 2170 3250
rect 2090 3190 2170 3210
rect 2330 3250 2410 3270
rect 2330 3210 2350 3250
rect 2390 3210 2410 3250
rect 2330 3190 2410 3210
rect 2570 3250 2650 3270
rect 2570 3210 2590 3250
rect 2630 3210 2650 3250
rect 2570 3190 2650 3210
rect 9120 3200 9200 3220
rect 440 3130 500 3180
rect 9120 3160 9140 3200
rect 9180 3160 9200 3200
rect 440 3090 450 3130
rect 490 3090 500 3130
rect 440 3030 500 3090
rect 440 2990 450 3030
rect 490 2990 500 3030
rect 440 2930 500 2990
rect 440 2890 450 2930
rect 490 2890 500 2930
rect 440 2830 500 2890
rect 440 2790 450 2830
rect 490 2790 500 2830
rect 440 2730 500 2790
rect 440 2690 450 2730
rect 490 2690 500 2730
rect 440 2670 500 2690
rect 1520 3130 1740 3150
rect 1520 3090 1530 3130
rect 1570 3090 1610 3130
rect 1650 3090 1690 3130
rect 1730 3090 1740 3130
rect 1520 3030 1740 3090
rect 1520 2990 1530 3030
rect 1570 2990 1610 3030
rect 1650 2990 1690 3030
rect 1730 2990 1740 3030
rect 1520 2930 1740 2990
rect 1520 2890 1530 2930
rect 1570 2890 1610 2930
rect 1650 2890 1690 2930
rect 1730 2890 1740 2930
rect 1520 2830 1740 2890
rect 1520 2790 1530 2830
rect 1570 2790 1610 2830
rect 1650 2790 1690 2830
rect 1730 2790 1740 2830
rect 1520 2730 1740 2790
rect 1520 2690 1530 2730
rect 1570 2690 1610 2730
rect 1650 2690 1690 2730
rect 1730 2690 1740 2730
rect 1520 2670 1740 2690
rect 2760 3130 2820 3150
rect 9120 3140 9200 3160
rect 2760 3090 2770 3130
rect 2810 3090 2820 3130
rect 2760 3030 2820 3090
rect 2760 2990 2770 3030
rect 2810 2990 2820 3030
rect 2760 2930 2820 2990
rect 2760 2890 2770 2930
rect 2810 2890 2820 2930
rect 2760 2830 2820 2890
rect 2760 2790 2770 2830
rect 2810 2790 2820 2830
rect 9320 2880 9420 2900
rect 9320 2820 9340 2880
rect 9400 2820 9420 2880
rect 9320 2800 9420 2820
rect 2760 2730 2820 2790
rect 2760 2690 2770 2730
rect 2810 2690 2820 2730
rect 2760 2670 2820 2690
rect -1070 2630 -1030 2670
rect 1610 2630 1650 2670
rect -1090 2610 -1010 2630
rect -1090 2570 -1070 2610
rect -1030 2570 -1010 2610
rect -1090 2550 -1010 2570
rect 1590 2610 1670 2630
rect 1590 2570 1610 2610
rect 1650 2570 1670 2610
rect 1590 2550 1670 2570
rect -1830 2340 -1750 2360
rect -1830 2300 -1810 2340
rect -1770 2300 -1750 2340
rect -1830 2280 -1750 2300
rect -1670 2340 -1590 2360
rect -1670 2300 -1650 2340
rect -1610 2300 -1590 2340
rect -1670 2280 -1590 2300
rect -1510 2340 -1430 2360
rect -1510 2300 -1490 2340
rect -1450 2300 -1430 2340
rect -1510 2280 -1430 2300
rect -1350 2340 -1270 2360
rect -1350 2300 -1330 2340
rect -1290 2300 -1270 2340
rect -1350 2280 -1270 2300
rect -1190 2340 -1110 2360
rect -1190 2300 -1170 2340
rect -1130 2300 -1110 2340
rect -1190 2280 -1110 2300
rect -1030 2340 -950 2360
rect -1030 2300 -1010 2340
rect -970 2300 -950 2340
rect -1030 2280 -950 2300
rect -870 2340 -790 2360
rect -870 2300 -850 2340
rect -810 2300 -790 2340
rect -870 2280 -790 2300
rect -710 2340 -630 2360
rect -710 2300 -690 2340
rect -650 2300 -630 2340
rect -710 2280 -630 2300
rect -550 2340 -470 2360
rect -550 2300 -530 2340
rect -490 2300 -470 2340
rect -550 2280 -470 2300
rect -390 2340 -310 2360
rect -390 2300 -370 2340
rect -330 2300 -310 2340
rect -390 2280 -310 2300
rect -230 2340 -150 2360
rect -230 2300 -210 2340
rect -170 2300 -150 2340
rect -230 2280 -150 2300
rect -70 2340 10 2360
rect -70 2300 -50 2340
rect -10 2300 10 2340
rect -70 2280 10 2300
rect 90 2340 170 2360
rect 90 2300 110 2340
rect 150 2300 170 2340
rect 90 2280 170 2300
rect 250 2340 330 2360
rect 250 2300 270 2340
rect 310 2300 330 2340
rect 250 2280 330 2300
rect 410 2340 490 2360
rect 410 2300 430 2340
rect 470 2300 490 2340
rect 410 2280 490 2300
rect 570 2340 650 2360
rect 570 2300 590 2340
rect 630 2300 650 2340
rect 570 2280 650 2300
rect 730 2340 810 2360
rect 730 2300 750 2340
rect 790 2300 810 2340
rect 730 2280 810 2300
rect 890 2340 970 2360
rect 890 2300 910 2340
rect 950 2300 970 2340
rect 890 2280 970 2300
rect 1050 2340 1130 2360
rect 1050 2300 1070 2340
rect 1110 2300 1130 2340
rect 1050 2280 1130 2300
rect 1210 2340 1290 2360
rect 1210 2300 1230 2340
rect 1270 2300 1290 2340
rect 1210 2280 1290 2300
rect 1370 2340 1450 2360
rect 1370 2300 1390 2340
rect 1430 2300 1450 2340
rect 1370 2280 1450 2300
rect 1530 2340 1610 2360
rect 1530 2300 1550 2340
rect 1590 2300 1610 2340
rect 1530 2280 1610 2300
rect 1690 2340 1770 2360
rect 1690 2300 1710 2340
rect 1750 2300 1770 2340
rect 1690 2280 1770 2300
rect 1850 2340 1930 2360
rect 1850 2300 1870 2340
rect 1910 2300 1930 2340
rect 1850 2280 1930 2300
rect 2010 2340 2090 2360
rect 2010 2300 2030 2340
rect 2070 2300 2090 2340
rect 2010 2280 2090 2300
rect 2170 2340 2250 2360
rect 2170 2300 2190 2340
rect 2230 2300 2250 2340
rect 2170 2280 2250 2300
rect -1810 2240 -1770 2280
rect 270 2240 310 2280
rect -1820 2220 -1760 2240
rect -1820 2190 -1810 2220
rect -1910 2180 -1810 2190
rect -1770 2180 -1760 2220
rect -1910 2170 -1760 2180
rect -1910 2130 -1890 2170
rect -1850 2130 -1760 2170
rect -1910 2120 -1760 2130
rect -1910 2110 -1810 2120
rect -1820 2080 -1810 2110
rect -1770 2080 -1760 2120
rect -1820 2060 -1760 2080
rect 260 2220 320 2240
rect 260 2180 270 2220
rect 310 2180 320 2220
rect 260 2120 320 2180
rect 260 2080 270 2120
rect 310 2080 320 2120
rect 260 2060 320 2080
rect 2340 2230 2480 2240
rect 2340 2220 2560 2230
rect 2340 2180 2350 2220
rect 2390 2180 2430 2220
rect 2470 2210 2560 2220
rect 2470 2180 2500 2210
rect 2340 2170 2500 2180
rect 2540 2170 2560 2210
rect 2340 2130 2560 2170
rect 2340 2120 2500 2130
rect 2340 2080 2350 2120
rect 2390 2080 2430 2120
rect 2470 2090 2500 2120
rect 2540 2090 2560 2130
rect 2470 2080 2560 2090
rect 2340 2070 2560 2080
rect 2340 2060 2480 2070
rect -448 1780 -358 1790
rect -448 1730 -428 1780
rect -378 1730 -358 1780
rect -448 1720 -358 1730
rect 950 1780 1040 1790
rect 950 1730 970 1780
rect 1020 1730 1040 1780
rect 950 1720 1040 1730
rect -1720 1519 2300 1560
rect -1720 1496 -1580 1519
rect -1720 1462 -1681 1496
rect -1647 1485 -1580 1496
rect -1546 1485 -1490 1519
rect -1456 1485 -1400 1519
rect -1366 1485 -1310 1519
rect -1276 1485 -1220 1519
rect -1186 1485 -1130 1519
rect -1096 1485 -1040 1519
rect -1006 1485 -950 1519
rect -916 1485 -860 1519
rect -826 1485 -770 1519
rect -736 1485 -680 1519
rect -646 1485 -590 1519
rect -556 1496 -220 1519
rect -556 1485 -494 1496
rect -1647 1462 -494 1485
rect -460 1462 -321 1496
rect -287 1485 -220 1496
rect -186 1485 -130 1519
rect -96 1485 -40 1519
rect -6 1485 50 1519
rect 84 1485 140 1519
rect 174 1485 230 1519
rect 264 1485 320 1519
rect 354 1485 410 1519
rect 444 1485 500 1519
rect 534 1485 590 1519
rect 624 1485 680 1519
rect 714 1485 770 1519
rect 804 1496 1140 1519
rect 804 1485 866 1496
rect -287 1462 866 1485
rect 900 1462 1039 1496
rect 1073 1485 1140 1496
rect 1174 1485 1230 1519
rect 1264 1485 1320 1519
rect 1354 1485 1410 1519
rect 1444 1485 1500 1519
rect 1534 1485 1590 1519
rect 1624 1485 1680 1519
rect 1714 1485 1770 1519
rect 1804 1485 1860 1519
rect 1894 1485 1950 1519
rect 1984 1485 2040 1519
rect 2074 1485 2130 1519
rect 2164 1496 2300 1519
rect 2164 1485 2226 1496
rect 1073 1462 2226 1485
rect 2260 1462 2300 1496
rect -1720 1406 2300 1462
rect -1720 1372 -1681 1406
rect -1647 1372 -494 1406
rect -460 1372 -321 1406
rect -287 1372 866 1406
rect 900 1372 1039 1406
rect 1073 1372 2226 1406
rect 2260 1372 2300 1406
rect -1720 1338 -1474 1372
rect -1440 1338 -1384 1372
rect -1350 1338 -1294 1372
rect -1260 1338 -1204 1372
rect -1170 1338 -1114 1372
rect -1080 1338 -1024 1372
rect -990 1338 -934 1372
rect -900 1338 -844 1372
rect -810 1338 -754 1372
rect -720 1338 -114 1372
rect -80 1338 -24 1372
rect 10 1338 66 1372
rect 100 1338 156 1372
rect 190 1338 246 1372
rect 280 1338 336 1372
rect 370 1338 426 1372
rect 460 1338 516 1372
rect 550 1338 606 1372
rect 640 1338 1246 1372
rect 1280 1338 1336 1372
rect 1370 1338 1426 1372
rect 1460 1338 1516 1372
rect 1550 1338 1606 1372
rect 1640 1338 1696 1372
rect 1730 1338 1786 1372
rect 1820 1338 1876 1372
rect 1910 1338 1966 1372
rect 2000 1338 2300 1372
rect -1720 1316 2300 1338
rect -1720 1310 -1681 1316
rect -1714 1282 -1681 1310
rect -1647 1315 -494 1316
rect -1647 1310 -642 1315
rect -1647 1282 -1615 1310
rect -1714 1226 -1615 1282
rect -1714 1192 -1681 1226
rect -1647 1192 -1615 1226
rect -1714 1136 -1615 1192
rect -1714 1102 -1681 1136
rect -1647 1102 -1615 1136
rect -1714 1046 -1615 1102
rect -1714 1012 -1681 1046
rect -1647 1012 -1615 1046
rect -1714 956 -1615 1012
rect -1714 922 -1681 956
rect -1647 922 -1615 956
rect -1714 866 -1615 922
rect -1714 832 -1681 866
rect -1647 832 -1615 866
rect -1714 776 -1615 832
rect -1714 742 -1681 776
rect -1647 742 -1615 776
rect -1714 686 -1615 742
rect -1714 652 -1681 686
rect -1647 652 -1615 686
rect -1714 596 -1615 652
rect -1714 562 -1681 596
rect -1647 562 -1615 596
rect -1714 506 -1615 562
rect -1714 472 -1681 506
rect -1647 472 -1615 506
rect -1714 416 -1615 472
rect -1551 1296 -1479 1310
rect -1551 1262 -1532 1296
rect -1498 1262 -1479 1296
rect -1551 1206 -1479 1262
rect -661 1281 -642 1310
rect -608 1310 -494 1315
rect -608 1281 -589 1310
rect -1551 1172 -1532 1206
rect -1498 1172 -1479 1206
rect -1551 1116 -1479 1172
rect -1551 1082 -1532 1116
rect -1498 1082 -1479 1116
rect -1551 1026 -1479 1082
rect -1551 992 -1532 1026
rect -1498 992 -1479 1026
rect -1551 936 -1479 992
rect -1551 902 -1532 936
rect -1498 902 -1479 936
rect -1551 846 -1479 902
rect -1551 812 -1532 846
rect -1498 812 -1479 846
rect -1551 756 -1479 812
rect -1551 722 -1532 756
rect -1498 722 -1479 756
rect -1551 666 -1479 722
rect -1551 632 -1532 666
rect -1498 632 -1479 666
rect -1551 576 -1479 632
rect -1551 542 -1532 576
rect -1498 542 -1479 576
rect -1417 1198 -723 1257
rect -1417 1164 -1358 1198
rect -1324 1170 -1268 1198
rect -1296 1164 -1268 1170
rect -1234 1170 -1178 1198
rect -1234 1164 -1230 1170
rect -1417 1136 -1330 1164
rect -1296 1136 -1230 1164
rect -1196 1164 -1178 1170
rect -1144 1170 -1088 1198
rect -1144 1164 -1130 1170
rect -1196 1136 -1130 1164
rect -1096 1164 -1088 1170
rect -1054 1170 -998 1198
rect -964 1170 -908 1198
rect -874 1170 -818 1198
rect -1054 1164 -1030 1170
rect -964 1164 -930 1170
rect -874 1164 -830 1170
rect -784 1164 -723 1198
rect -1096 1136 -1030 1164
rect -996 1136 -930 1164
rect -896 1136 -830 1164
rect -796 1136 -723 1164
rect -1417 1108 -723 1136
rect -1417 1074 -1358 1108
rect -1324 1074 -1268 1108
rect -1234 1074 -1178 1108
rect -1144 1074 -1088 1108
rect -1054 1074 -998 1108
rect -964 1074 -908 1108
rect -874 1074 -818 1108
rect -784 1074 -723 1108
rect -1417 1070 -723 1074
rect -1417 1036 -1330 1070
rect -1296 1036 -1230 1070
rect -1196 1036 -1130 1070
rect -1096 1036 -1030 1070
rect -996 1036 -930 1070
rect -896 1036 -830 1070
rect -796 1036 -723 1070
rect -1417 1018 -723 1036
rect -1417 984 -1358 1018
rect -1324 984 -1268 1018
rect -1234 984 -1178 1018
rect -1144 984 -1088 1018
rect -1054 984 -998 1018
rect -964 984 -908 1018
rect -874 984 -818 1018
rect -784 984 -723 1018
rect -1417 970 -723 984
rect -1417 936 -1330 970
rect -1296 936 -1230 970
rect -1196 936 -1130 970
rect -1096 936 -1030 970
rect -996 936 -930 970
rect -896 936 -830 970
rect -796 936 -723 970
rect -1417 928 -723 936
rect -1417 894 -1358 928
rect -1324 894 -1268 928
rect -1234 894 -1178 928
rect -1144 894 -1088 928
rect -1054 894 -998 928
rect -964 894 -908 928
rect -874 894 -818 928
rect -784 894 -723 928
rect -1417 870 -723 894
rect -1417 838 -1330 870
rect -1296 838 -1230 870
rect -1417 804 -1358 838
rect -1296 836 -1268 838
rect -1324 804 -1268 836
rect -1234 836 -1230 838
rect -1196 838 -1130 870
rect -1196 836 -1178 838
rect -1234 804 -1178 836
rect -1144 836 -1130 838
rect -1096 838 -1030 870
rect -996 838 -930 870
rect -896 838 -830 870
rect -796 838 -723 870
rect -1096 836 -1088 838
rect -1144 804 -1088 836
rect -1054 836 -1030 838
rect -964 836 -930 838
rect -874 836 -830 838
rect -1054 804 -998 836
rect -964 804 -908 836
rect -874 804 -818 836
rect -784 804 -723 838
rect -1417 770 -723 804
rect -1417 748 -1330 770
rect -1296 748 -1230 770
rect -1417 714 -1358 748
rect -1296 736 -1268 748
rect -1324 714 -1268 736
rect -1234 736 -1230 748
rect -1196 748 -1130 770
rect -1196 736 -1178 748
rect -1234 714 -1178 736
rect -1144 736 -1130 748
rect -1096 748 -1030 770
rect -996 748 -930 770
rect -896 748 -830 770
rect -796 748 -723 770
rect -1096 736 -1088 748
rect -1144 714 -1088 736
rect -1054 736 -1030 748
rect -964 736 -930 748
rect -874 736 -830 748
rect -1054 714 -998 736
rect -964 714 -908 736
rect -874 714 -818 736
rect -784 714 -723 748
rect -1417 670 -723 714
rect -1417 658 -1330 670
rect -1296 658 -1230 670
rect -1417 624 -1358 658
rect -1296 636 -1268 658
rect -1324 624 -1268 636
rect -1234 636 -1230 658
rect -1196 658 -1130 670
rect -1196 636 -1178 658
rect -1234 624 -1178 636
rect -1144 636 -1130 658
rect -1096 658 -1030 670
rect -996 658 -930 670
rect -896 658 -830 670
rect -796 658 -723 670
rect -1096 636 -1088 658
rect -1144 624 -1088 636
rect -1054 636 -1030 658
rect -964 636 -930 658
rect -874 636 -830 658
rect -1054 624 -998 636
rect -964 624 -908 636
rect -874 624 -818 636
rect -784 624 -723 658
rect -1417 563 -723 624
rect -661 1225 -589 1281
rect -661 1191 -642 1225
rect -608 1191 -589 1225
rect -661 1135 -589 1191
rect -661 1101 -642 1135
rect -608 1101 -589 1135
rect -661 1045 -589 1101
rect -661 1011 -642 1045
rect -608 1011 -589 1045
rect -661 955 -589 1011
rect -661 921 -642 955
rect -608 921 -589 955
rect -661 865 -589 921
rect -661 831 -642 865
rect -608 831 -589 865
rect -661 775 -589 831
rect -661 741 -642 775
rect -608 741 -589 775
rect -661 685 -589 741
rect -661 651 -642 685
rect -608 651 -589 685
rect -661 595 -589 651
rect -1551 501 -1479 542
rect -661 561 -642 595
rect -608 561 -589 595
rect -661 501 -589 561
rect -1551 482 -589 501
rect -1551 448 -1440 482
rect -1406 448 -1350 482
rect -1316 448 -1260 482
rect -1226 448 -1170 482
rect -1136 448 -1080 482
rect -1046 448 -990 482
rect -956 448 -900 482
rect -866 448 -810 482
rect -776 448 -720 482
rect -686 448 -589 482
rect -1551 429 -589 448
rect -525 1282 -494 1310
rect -460 1282 -321 1316
rect -287 1315 866 1316
rect -287 1310 718 1315
rect -287 1282 -255 1310
rect -525 1226 -255 1282
rect -525 1192 -494 1226
rect -460 1192 -321 1226
rect -287 1192 -255 1226
rect -525 1136 -255 1192
rect -525 1102 -494 1136
rect -460 1102 -321 1136
rect -287 1102 -255 1136
rect -525 1046 -255 1102
rect -525 1012 -494 1046
rect -460 1012 -321 1046
rect -287 1012 -255 1046
rect -525 956 -255 1012
rect -525 922 -494 956
rect -460 922 -321 956
rect -287 922 -255 956
rect -525 866 -255 922
rect -525 832 -494 866
rect -460 832 -321 866
rect -287 832 -255 866
rect -525 776 -255 832
rect -525 742 -494 776
rect -460 742 -321 776
rect -287 742 -255 776
rect -525 686 -255 742
rect -525 652 -494 686
rect -460 652 -321 686
rect -287 652 -255 686
rect -525 596 -255 652
rect -525 562 -494 596
rect -460 562 -321 596
rect -287 562 -255 596
rect -525 506 -255 562
rect -525 472 -494 506
rect -460 472 -321 506
rect -287 472 -255 506
rect -1714 382 -1681 416
rect -1647 382 -1615 416
rect -1714 365 -1615 382
rect -525 416 -255 472
rect -191 1296 -119 1310
rect -191 1262 -172 1296
rect -138 1262 -119 1296
rect -191 1206 -119 1262
rect 699 1281 718 1310
rect 752 1310 866 1315
rect 752 1281 771 1310
rect -191 1172 -172 1206
rect -138 1172 -119 1206
rect -191 1116 -119 1172
rect -191 1082 -172 1116
rect -138 1082 -119 1116
rect -191 1026 -119 1082
rect -191 992 -172 1026
rect -138 992 -119 1026
rect -191 936 -119 992
rect -191 902 -172 936
rect -138 902 -119 936
rect -191 846 -119 902
rect -191 812 -172 846
rect -138 812 -119 846
rect -191 756 -119 812
rect -191 722 -172 756
rect -138 722 -119 756
rect -191 666 -119 722
rect -191 632 -172 666
rect -138 632 -119 666
rect -191 576 -119 632
rect -191 542 -172 576
rect -138 542 -119 576
rect -57 1198 637 1257
rect -57 1164 2 1198
rect 36 1170 92 1198
rect 64 1164 92 1170
rect 126 1170 182 1198
rect 126 1164 130 1170
rect -57 1136 30 1164
rect 64 1136 130 1164
rect 164 1164 182 1170
rect 216 1170 272 1198
rect 216 1164 230 1170
rect 164 1136 230 1164
rect 264 1164 272 1170
rect 306 1170 362 1198
rect 396 1170 452 1198
rect 486 1170 542 1198
rect 306 1164 330 1170
rect 396 1164 430 1170
rect 486 1164 530 1170
rect 576 1164 637 1198
rect 264 1136 330 1164
rect 364 1136 430 1164
rect 464 1136 530 1164
rect 564 1136 637 1164
rect -57 1108 637 1136
rect -57 1074 2 1108
rect 36 1074 92 1108
rect 126 1074 182 1108
rect 216 1074 272 1108
rect 306 1074 362 1108
rect 396 1074 452 1108
rect 486 1074 542 1108
rect 576 1074 637 1108
rect -57 1070 637 1074
rect -57 1036 30 1070
rect 64 1036 130 1070
rect 164 1036 230 1070
rect 264 1036 330 1070
rect 364 1036 430 1070
rect 464 1036 530 1070
rect 564 1036 637 1070
rect -57 1018 637 1036
rect -57 984 2 1018
rect 36 984 92 1018
rect 126 984 182 1018
rect 216 984 272 1018
rect 306 984 362 1018
rect 396 984 452 1018
rect 486 984 542 1018
rect 576 984 637 1018
rect -57 970 637 984
rect -57 936 30 970
rect 64 936 130 970
rect 164 936 230 970
rect 264 936 330 970
rect 364 936 430 970
rect 464 936 530 970
rect 564 936 637 970
rect -57 928 637 936
rect -57 894 2 928
rect 36 894 92 928
rect 126 894 182 928
rect 216 894 272 928
rect 306 894 362 928
rect 396 894 452 928
rect 486 894 542 928
rect 576 894 637 928
rect -57 870 637 894
rect -57 838 30 870
rect 64 838 130 870
rect -57 804 2 838
rect 64 836 92 838
rect 36 804 92 836
rect 126 836 130 838
rect 164 838 230 870
rect 164 836 182 838
rect 126 804 182 836
rect 216 836 230 838
rect 264 838 330 870
rect 364 838 430 870
rect 464 838 530 870
rect 564 838 637 870
rect 264 836 272 838
rect 216 804 272 836
rect 306 836 330 838
rect 396 836 430 838
rect 486 836 530 838
rect 306 804 362 836
rect 396 804 452 836
rect 486 804 542 836
rect 576 804 637 838
rect -57 770 637 804
rect -57 748 30 770
rect 64 748 130 770
rect -57 714 2 748
rect 64 736 92 748
rect 36 714 92 736
rect 126 736 130 748
rect 164 748 230 770
rect 164 736 182 748
rect 126 714 182 736
rect 216 736 230 748
rect 264 748 330 770
rect 364 748 430 770
rect 464 748 530 770
rect 564 748 637 770
rect 264 736 272 748
rect 216 714 272 736
rect 306 736 330 748
rect 396 736 430 748
rect 486 736 530 748
rect 306 714 362 736
rect 396 714 452 736
rect 486 714 542 736
rect 576 714 637 748
rect -57 670 637 714
rect -57 658 30 670
rect 64 658 130 670
rect -57 624 2 658
rect 64 636 92 658
rect 36 624 92 636
rect 126 636 130 658
rect 164 658 230 670
rect 164 636 182 658
rect 126 624 182 636
rect 216 636 230 658
rect 264 658 330 670
rect 364 658 430 670
rect 464 658 530 670
rect 564 658 637 670
rect 264 636 272 658
rect 216 624 272 636
rect 306 636 330 658
rect 396 636 430 658
rect 486 636 530 658
rect 306 624 362 636
rect 396 624 452 636
rect 486 624 542 636
rect 576 624 637 658
rect -57 563 637 624
rect 699 1225 771 1281
rect 699 1191 718 1225
rect 752 1191 771 1225
rect 699 1135 771 1191
rect 699 1101 718 1135
rect 752 1101 771 1135
rect 699 1045 771 1101
rect 699 1011 718 1045
rect 752 1011 771 1045
rect 699 955 771 1011
rect 699 921 718 955
rect 752 921 771 955
rect 699 865 771 921
rect 699 831 718 865
rect 752 831 771 865
rect 699 775 771 831
rect 699 741 718 775
rect 752 741 771 775
rect 699 685 771 741
rect 699 651 718 685
rect 752 651 771 685
rect 699 595 771 651
rect -191 501 -119 542
rect 699 561 718 595
rect 752 561 771 595
rect 699 501 771 561
rect -191 482 771 501
rect -191 448 -80 482
rect -46 448 10 482
rect 44 448 100 482
rect 134 448 190 482
rect 224 448 280 482
rect 314 448 370 482
rect 404 448 460 482
rect 494 448 550 482
rect 584 448 640 482
rect 674 448 771 482
rect -191 429 771 448
rect 835 1282 866 1310
rect 900 1282 1039 1316
rect 1073 1315 2226 1316
rect 1073 1310 2078 1315
rect 1073 1282 1105 1310
rect 835 1226 1105 1282
rect 835 1192 866 1226
rect 900 1192 1039 1226
rect 1073 1192 1105 1226
rect 835 1136 1105 1192
rect 835 1102 866 1136
rect 900 1102 1039 1136
rect 1073 1102 1105 1136
rect 835 1046 1105 1102
rect 835 1012 866 1046
rect 900 1012 1039 1046
rect 1073 1012 1105 1046
rect 835 956 1105 1012
rect 835 922 866 956
rect 900 922 1039 956
rect 1073 922 1105 956
rect 835 866 1105 922
rect 835 832 866 866
rect 900 832 1039 866
rect 1073 832 1105 866
rect 835 776 1105 832
rect 835 742 866 776
rect 900 742 1039 776
rect 1073 742 1105 776
rect 835 686 1105 742
rect 835 652 866 686
rect 900 652 1039 686
rect 1073 652 1105 686
rect 835 596 1105 652
rect 835 562 866 596
rect 900 562 1039 596
rect 1073 562 1105 596
rect 835 506 1105 562
rect 835 472 866 506
rect 900 472 1039 506
rect 1073 472 1105 506
rect -525 382 -494 416
rect -460 382 -321 416
rect -287 382 -255 416
rect -525 365 -255 382
rect 835 416 1105 472
rect 1169 1296 1241 1310
rect 1169 1262 1188 1296
rect 1222 1262 1241 1296
rect 1169 1206 1241 1262
rect 2059 1281 2078 1310
rect 2112 1310 2226 1315
rect 2112 1281 2131 1310
rect 1169 1172 1188 1206
rect 1222 1172 1241 1206
rect 1169 1116 1241 1172
rect 1169 1082 1188 1116
rect 1222 1082 1241 1116
rect 1169 1026 1241 1082
rect 1169 992 1188 1026
rect 1222 992 1241 1026
rect 1169 936 1241 992
rect 1169 902 1188 936
rect 1222 902 1241 936
rect 1169 846 1241 902
rect 1169 812 1188 846
rect 1222 812 1241 846
rect 1169 756 1241 812
rect 1169 722 1188 756
rect 1222 722 1241 756
rect 1169 666 1241 722
rect 1169 632 1188 666
rect 1222 632 1241 666
rect 1169 576 1241 632
rect 1169 542 1188 576
rect 1222 542 1241 576
rect 1303 1198 1997 1257
rect 1303 1164 1362 1198
rect 1396 1170 1452 1198
rect 1424 1164 1452 1170
rect 1486 1170 1542 1198
rect 1486 1164 1490 1170
rect 1303 1136 1390 1164
rect 1424 1136 1490 1164
rect 1524 1164 1542 1170
rect 1576 1170 1632 1198
rect 1576 1164 1590 1170
rect 1524 1136 1590 1164
rect 1624 1164 1632 1170
rect 1666 1170 1722 1198
rect 1756 1170 1812 1198
rect 1846 1170 1902 1198
rect 1666 1164 1690 1170
rect 1756 1164 1790 1170
rect 1846 1164 1890 1170
rect 1936 1164 1997 1198
rect 1624 1136 1690 1164
rect 1724 1136 1790 1164
rect 1824 1136 1890 1164
rect 1924 1136 1997 1164
rect 1303 1108 1997 1136
rect 1303 1074 1362 1108
rect 1396 1074 1452 1108
rect 1486 1074 1542 1108
rect 1576 1074 1632 1108
rect 1666 1074 1722 1108
rect 1756 1074 1812 1108
rect 1846 1074 1902 1108
rect 1936 1074 1997 1108
rect 1303 1070 1997 1074
rect 1303 1036 1390 1070
rect 1424 1036 1490 1070
rect 1524 1036 1590 1070
rect 1624 1036 1690 1070
rect 1724 1036 1790 1070
rect 1824 1036 1890 1070
rect 1924 1036 1997 1070
rect 1303 1018 1997 1036
rect 1303 984 1362 1018
rect 1396 984 1452 1018
rect 1486 984 1542 1018
rect 1576 984 1632 1018
rect 1666 984 1722 1018
rect 1756 984 1812 1018
rect 1846 984 1902 1018
rect 1936 984 1997 1018
rect 1303 970 1997 984
rect 1303 936 1390 970
rect 1424 936 1490 970
rect 1524 936 1590 970
rect 1624 936 1690 970
rect 1724 936 1790 970
rect 1824 936 1890 970
rect 1924 936 1997 970
rect 1303 928 1997 936
rect 1303 894 1362 928
rect 1396 894 1452 928
rect 1486 894 1542 928
rect 1576 894 1632 928
rect 1666 894 1722 928
rect 1756 894 1812 928
rect 1846 894 1902 928
rect 1936 894 1997 928
rect 1303 870 1997 894
rect 1303 838 1390 870
rect 1424 838 1490 870
rect 1303 804 1362 838
rect 1424 836 1452 838
rect 1396 804 1452 836
rect 1486 836 1490 838
rect 1524 838 1590 870
rect 1524 836 1542 838
rect 1486 804 1542 836
rect 1576 836 1590 838
rect 1624 838 1690 870
rect 1724 838 1790 870
rect 1824 838 1890 870
rect 1924 838 1997 870
rect 1624 836 1632 838
rect 1576 804 1632 836
rect 1666 836 1690 838
rect 1756 836 1790 838
rect 1846 836 1890 838
rect 1666 804 1722 836
rect 1756 804 1812 836
rect 1846 804 1902 836
rect 1936 804 1997 838
rect 1303 770 1997 804
rect 1303 748 1390 770
rect 1424 748 1490 770
rect 1303 714 1362 748
rect 1424 736 1452 748
rect 1396 714 1452 736
rect 1486 736 1490 748
rect 1524 748 1590 770
rect 1524 736 1542 748
rect 1486 714 1542 736
rect 1576 736 1590 748
rect 1624 748 1690 770
rect 1724 748 1790 770
rect 1824 748 1890 770
rect 1924 748 1997 770
rect 1624 736 1632 748
rect 1576 714 1632 736
rect 1666 736 1690 748
rect 1756 736 1790 748
rect 1846 736 1890 748
rect 1666 714 1722 736
rect 1756 714 1812 736
rect 1846 714 1902 736
rect 1936 714 1997 748
rect 1303 670 1997 714
rect 1303 658 1390 670
rect 1424 658 1490 670
rect 1303 624 1362 658
rect 1424 636 1452 658
rect 1396 624 1452 636
rect 1486 636 1490 658
rect 1524 658 1590 670
rect 1524 636 1542 658
rect 1486 624 1542 636
rect 1576 636 1590 658
rect 1624 658 1690 670
rect 1724 658 1790 670
rect 1824 658 1890 670
rect 1924 658 1997 670
rect 1624 636 1632 658
rect 1576 624 1632 636
rect 1666 636 1690 658
rect 1756 636 1790 658
rect 1846 636 1890 658
rect 1666 624 1722 636
rect 1756 624 1812 636
rect 1846 624 1902 636
rect 1936 624 1997 658
rect 1303 563 1997 624
rect 2059 1225 2131 1281
rect 2059 1191 2078 1225
rect 2112 1191 2131 1225
rect 2059 1135 2131 1191
rect 2059 1101 2078 1135
rect 2112 1101 2131 1135
rect 2059 1045 2131 1101
rect 2059 1011 2078 1045
rect 2112 1011 2131 1045
rect 2059 955 2131 1011
rect 2059 921 2078 955
rect 2112 921 2131 955
rect 2059 865 2131 921
rect 2059 831 2078 865
rect 2112 831 2131 865
rect 2059 775 2131 831
rect 2059 741 2078 775
rect 2112 741 2131 775
rect 2059 685 2131 741
rect 2059 651 2078 685
rect 2112 651 2131 685
rect 2059 595 2131 651
rect 1169 501 1241 542
rect 2059 561 2078 595
rect 2112 561 2131 595
rect 2059 501 2131 561
rect 1169 482 2131 501
rect 1169 448 1280 482
rect 1314 448 1370 482
rect 1404 448 1460 482
rect 1494 448 1550 482
rect 1584 448 1640 482
rect 1674 448 1730 482
rect 1764 448 1820 482
rect 1854 448 1910 482
rect 1944 448 2000 482
rect 2034 448 2131 482
rect 1169 429 2131 448
rect 2195 1282 2226 1310
rect 2260 1310 2300 1316
rect 2260 1282 2294 1310
rect 2195 1226 2294 1282
rect 2195 1192 2226 1226
rect 2260 1192 2294 1226
rect 2195 1136 2294 1192
rect 2195 1102 2226 1136
rect 2260 1102 2294 1136
rect 2195 1046 2294 1102
rect 2195 1012 2226 1046
rect 2260 1012 2294 1046
rect 2195 956 2294 1012
rect 2195 922 2226 956
rect 2260 922 2294 956
rect 2195 866 2294 922
rect 2195 832 2226 866
rect 2260 832 2294 866
rect 2195 776 2294 832
rect 2195 742 2226 776
rect 2260 742 2294 776
rect 2195 686 2294 742
rect 2195 652 2226 686
rect 2260 652 2294 686
rect 2195 596 2294 652
rect 2195 562 2226 596
rect 2260 562 2294 596
rect 2195 506 2294 562
rect 2195 472 2226 506
rect 2260 472 2294 506
rect 835 382 866 416
rect 900 382 1039 416
rect 1073 382 1105 416
rect 835 365 1105 382
rect 2195 416 2294 472
rect 2195 382 2226 416
rect 2260 382 2294 416
rect 2195 365 2294 382
rect -1714 332 2294 365
rect -1714 298 -1580 332
rect -1546 298 -1490 332
rect -1456 298 -1400 332
rect -1366 298 -1310 332
rect -1276 298 -1220 332
rect -1186 298 -1130 332
rect -1096 298 -1040 332
rect -1006 298 -950 332
rect -916 298 -860 332
rect -826 298 -770 332
rect -736 298 -680 332
rect -646 298 -590 332
rect -556 298 -220 332
rect -186 298 -130 332
rect -96 298 -40 332
rect -6 298 50 332
rect 84 298 140 332
rect 174 298 230 332
rect 264 298 320 332
rect 354 298 410 332
rect 444 298 500 332
rect 534 298 590 332
rect 624 298 680 332
rect 714 298 770 332
rect 804 298 1140 332
rect 1174 298 1230 332
rect 1264 298 1320 332
rect 1354 298 1410 332
rect 1444 298 1500 332
rect 1534 298 1590 332
rect 1624 298 1680 332
rect 1714 298 1770 332
rect 1804 298 1860 332
rect 1894 298 1950 332
rect 1984 298 2040 332
rect 2074 298 2130 332
rect 2164 298 2294 332
rect -1714 266 2294 298
rect -430 200 -350 266
rect 930 200 1010 266
rect -1720 159 2300 200
rect -1720 136 -1580 159
rect -1720 102 -1681 136
rect -1647 125 -1580 136
rect -1546 125 -1490 159
rect -1456 125 -1400 159
rect -1366 125 -1310 159
rect -1276 125 -1220 159
rect -1186 125 -1130 159
rect -1096 125 -1040 159
rect -1006 125 -950 159
rect -916 125 -860 159
rect -826 125 -770 159
rect -736 125 -680 159
rect -646 125 -590 159
rect -556 136 -220 159
rect -556 125 -494 136
rect -1647 102 -494 125
rect -460 102 -321 136
rect -287 125 -220 136
rect -186 125 -130 159
rect -96 125 -40 159
rect -6 125 50 159
rect 84 125 140 159
rect 174 125 230 159
rect 264 125 320 159
rect 354 125 410 159
rect 444 125 500 159
rect 534 125 590 159
rect 624 125 680 159
rect 714 125 770 159
rect 804 136 1140 159
rect 804 125 866 136
rect -287 102 866 125
rect 900 102 1039 136
rect 1073 125 1140 136
rect 1174 125 1230 159
rect 1264 125 1320 159
rect 1354 125 1410 159
rect 1444 125 1500 159
rect 1534 125 1590 159
rect 1624 125 1680 159
rect 1714 125 1770 159
rect 1804 125 1860 159
rect 1894 125 1950 159
rect 1984 125 2040 159
rect 2074 125 2130 159
rect 2164 136 2300 159
rect 2164 125 2226 136
rect 1073 102 2226 125
rect 2260 102 2300 136
rect -1720 46 2300 102
rect -1720 12 -1681 46
rect -1647 12 -494 46
rect -460 12 -321 46
rect -287 12 866 46
rect 900 12 1039 46
rect 1073 12 2226 46
rect 2260 12 2300 46
rect -2310 -20 -2240 0
rect -2310 -70 -2300 -20
rect -2250 -70 -2240 -20
rect -1720 -22 -1474 12
rect -1440 -22 -1384 12
rect -1350 -22 -1294 12
rect -1260 -22 -1204 12
rect -1170 -22 -1114 12
rect -1080 -22 -1024 12
rect -990 -22 -934 12
rect -900 -22 -844 12
rect -810 -22 -754 12
rect -720 -22 -114 12
rect -80 -22 -24 12
rect 10 -22 66 12
rect 100 -22 156 12
rect 190 -22 246 12
rect 280 -22 336 12
rect 370 -22 426 12
rect 460 -22 516 12
rect 550 -22 606 12
rect 640 -22 1246 12
rect 1280 -22 1336 12
rect 1370 -22 1426 12
rect 1460 -22 1516 12
rect 1550 -22 1606 12
rect 1640 -22 1696 12
rect 1730 -22 1786 12
rect 1820 -22 1876 12
rect 1910 -22 1966 12
rect 2000 -22 2300 12
rect -1720 -44 2300 -22
rect -1720 -50 -1681 -44
rect -2310 -90 -2240 -70
rect -1714 -78 -1681 -50
rect -1647 -45 -494 -44
rect -1647 -50 -642 -45
rect -1647 -78 -1615 -50
rect -2740 -400 -2670 -380
rect -2860 -450 -2790 -430
rect -2860 -500 -2850 -450
rect -2800 -500 -2790 -450
rect -2860 -522 -2790 -500
rect -2740 -450 -2730 -400
rect -2680 -450 -2670 -400
rect -2740 -470 -2670 -450
rect -2550 -540 -2500 -470
rect -2120 -160 -2070 -90
rect -1714 -134 -1615 -78
rect -1714 -168 -1681 -134
rect -1647 -168 -1615 -134
rect -1714 -224 -1615 -168
rect -1714 -258 -1681 -224
rect -1647 -258 -1615 -224
rect -1714 -314 -1615 -258
rect -1714 -348 -1681 -314
rect -1647 -348 -1615 -314
rect -1714 -404 -1615 -348
rect -1714 -438 -1681 -404
rect -1647 -438 -1615 -404
rect -1714 -494 -1615 -438
rect -1714 -528 -1681 -494
rect -1647 -528 -1615 -494
rect -1714 -584 -1615 -528
rect -1714 -618 -1681 -584
rect -1647 -618 -1615 -584
rect -1714 -674 -1615 -618
rect -1714 -708 -1681 -674
rect -1647 -708 -1615 -674
rect -1714 -764 -1615 -708
rect -1714 -798 -1681 -764
rect -1647 -798 -1615 -764
rect -1714 -854 -1615 -798
rect -1714 -888 -1681 -854
rect -1647 -888 -1615 -854
rect -1714 -944 -1615 -888
rect -1551 -64 -1479 -50
rect -1551 -98 -1532 -64
rect -1498 -98 -1479 -64
rect -1551 -154 -1479 -98
rect -661 -79 -642 -50
rect -608 -50 -494 -45
rect -608 -79 -589 -50
rect -1551 -188 -1532 -154
rect -1498 -188 -1479 -154
rect -1551 -244 -1479 -188
rect -1551 -278 -1532 -244
rect -1498 -278 -1479 -244
rect -1551 -334 -1479 -278
rect -1551 -368 -1532 -334
rect -1498 -368 -1479 -334
rect -1551 -424 -1479 -368
rect -1551 -458 -1532 -424
rect -1498 -458 -1479 -424
rect -1551 -514 -1479 -458
rect -1551 -548 -1532 -514
rect -1498 -548 -1479 -514
rect -1551 -604 -1479 -548
rect -1551 -638 -1532 -604
rect -1498 -638 -1479 -604
rect -1551 -694 -1479 -638
rect -1551 -728 -1532 -694
rect -1498 -728 -1479 -694
rect -1551 -784 -1479 -728
rect -1551 -818 -1532 -784
rect -1498 -818 -1479 -784
rect -1417 -162 -723 -103
rect -1417 -196 -1358 -162
rect -1324 -190 -1268 -162
rect -1296 -196 -1268 -190
rect -1234 -190 -1178 -162
rect -1234 -196 -1230 -190
rect -1417 -224 -1330 -196
rect -1296 -224 -1230 -196
rect -1196 -196 -1178 -190
rect -1144 -190 -1088 -162
rect -1144 -196 -1130 -190
rect -1196 -224 -1130 -196
rect -1096 -196 -1088 -190
rect -1054 -190 -998 -162
rect -964 -190 -908 -162
rect -874 -190 -818 -162
rect -1054 -196 -1030 -190
rect -964 -196 -930 -190
rect -874 -196 -830 -190
rect -784 -196 -723 -162
rect -1096 -224 -1030 -196
rect -996 -224 -930 -196
rect -896 -224 -830 -196
rect -796 -224 -723 -196
rect -1417 -252 -723 -224
rect -1417 -286 -1358 -252
rect -1324 -286 -1268 -252
rect -1234 -286 -1178 -252
rect -1144 -286 -1088 -252
rect -1054 -286 -998 -252
rect -964 -286 -908 -252
rect -874 -286 -818 -252
rect -784 -286 -723 -252
rect -1417 -290 -723 -286
rect -1417 -324 -1330 -290
rect -1296 -324 -1230 -290
rect -1196 -324 -1130 -290
rect -1096 -324 -1030 -290
rect -996 -324 -930 -290
rect -896 -324 -830 -290
rect -796 -324 -723 -290
rect -1417 -342 -723 -324
rect -1417 -376 -1358 -342
rect -1324 -376 -1268 -342
rect -1234 -376 -1178 -342
rect -1144 -376 -1088 -342
rect -1054 -376 -998 -342
rect -964 -376 -908 -342
rect -874 -376 -818 -342
rect -784 -376 -723 -342
rect -1417 -390 -723 -376
rect -1417 -424 -1330 -390
rect -1296 -424 -1230 -390
rect -1196 -424 -1130 -390
rect -1096 -424 -1030 -390
rect -996 -424 -930 -390
rect -896 -424 -830 -390
rect -796 -424 -723 -390
rect -1417 -432 -723 -424
rect -1417 -466 -1358 -432
rect -1324 -466 -1268 -432
rect -1234 -466 -1178 -432
rect -1144 -466 -1088 -432
rect -1054 -466 -998 -432
rect -964 -466 -908 -432
rect -874 -466 -818 -432
rect -784 -466 -723 -432
rect -1417 -490 -723 -466
rect -1417 -522 -1330 -490
rect -1296 -522 -1230 -490
rect -1417 -556 -1358 -522
rect -1296 -524 -1268 -522
rect -1324 -556 -1268 -524
rect -1234 -524 -1230 -522
rect -1196 -522 -1130 -490
rect -1196 -524 -1178 -522
rect -1234 -556 -1178 -524
rect -1144 -524 -1130 -522
rect -1096 -522 -1030 -490
rect -996 -522 -930 -490
rect -896 -522 -830 -490
rect -796 -522 -723 -490
rect -1096 -524 -1088 -522
rect -1144 -556 -1088 -524
rect -1054 -524 -1030 -522
rect -964 -524 -930 -522
rect -874 -524 -830 -522
rect -1054 -556 -998 -524
rect -964 -556 -908 -524
rect -874 -556 -818 -524
rect -784 -556 -723 -522
rect -1417 -590 -723 -556
rect -1417 -612 -1330 -590
rect -1296 -612 -1230 -590
rect -1417 -646 -1358 -612
rect -1296 -624 -1268 -612
rect -1324 -646 -1268 -624
rect -1234 -624 -1230 -612
rect -1196 -612 -1130 -590
rect -1196 -624 -1178 -612
rect -1234 -646 -1178 -624
rect -1144 -624 -1130 -612
rect -1096 -612 -1030 -590
rect -996 -612 -930 -590
rect -896 -612 -830 -590
rect -796 -612 -723 -590
rect -1096 -624 -1088 -612
rect -1144 -646 -1088 -624
rect -1054 -624 -1030 -612
rect -964 -624 -930 -612
rect -874 -624 -830 -612
rect -1054 -646 -998 -624
rect -964 -646 -908 -624
rect -874 -646 -818 -624
rect -784 -646 -723 -612
rect -1417 -690 -723 -646
rect -1417 -702 -1330 -690
rect -1296 -702 -1230 -690
rect -1417 -736 -1358 -702
rect -1296 -724 -1268 -702
rect -1324 -736 -1268 -724
rect -1234 -724 -1230 -702
rect -1196 -702 -1130 -690
rect -1196 -724 -1178 -702
rect -1234 -736 -1178 -724
rect -1144 -724 -1130 -702
rect -1096 -702 -1030 -690
rect -996 -702 -930 -690
rect -896 -702 -830 -690
rect -796 -702 -723 -690
rect -1096 -724 -1088 -702
rect -1144 -736 -1088 -724
rect -1054 -724 -1030 -702
rect -964 -724 -930 -702
rect -874 -724 -830 -702
rect -1054 -736 -998 -724
rect -964 -736 -908 -724
rect -874 -736 -818 -724
rect -784 -736 -723 -702
rect -1417 -797 -723 -736
rect -661 -135 -589 -79
rect -661 -169 -642 -135
rect -608 -169 -589 -135
rect -661 -225 -589 -169
rect -661 -259 -642 -225
rect -608 -259 -589 -225
rect -661 -315 -589 -259
rect -661 -349 -642 -315
rect -608 -349 -589 -315
rect -661 -405 -589 -349
rect -661 -439 -642 -405
rect -608 -439 -589 -405
rect -661 -495 -589 -439
rect -661 -529 -642 -495
rect -608 -529 -589 -495
rect -661 -585 -589 -529
rect -661 -619 -642 -585
rect -608 -619 -589 -585
rect -661 -675 -589 -619
rect -661 -709 -642 -675
rect -608 -709 -589 -675
rect -661 -765 -589 -709
rect -1551 -859 -1479 -818
rect -661 -799 -642 -765
rect -608 -799 -589 -765
rect -661 -859 -589 -799
rect -1551 -878 -589 -859
rect -1551 -912 -1440 -878
rect -1406 -912 -1350 -878
rect -1316 -912 -1260 -878
rect -1226 -912 -1170 -878
rect -1136 -912 -1080 -878
rect -1046 -912 -990 -878
rect -956 -912 -900 -878
rect -866 -912 -810 -878
rect -776 -912 -720 -878
rect -686 -912 -589 -878
rect -1551 -931 -589 -912
rect -525 -78 -494 -50
rect -460 -78 -321 -44
rect -287 -45 866 -44
rect -287 -50 718 -45
rect -287 -78 -255 -50
rect -525 -134 -255 -78
rect -525 -168 -494 -134
rect -460 -168 -321 -134
rect -287 -168 -255 -134
rect -525 -224 -255 -168
rect -525 -258 -494 -224
rect -460 -258 -321 -224
rect -287 -258 -255 -224
rect -525 -314 -255 -258
rect -525 -348 -494 -314
rect -460 -348 -321 -314
rect -287 -348 -255 -314
rect -525 -404 -255 -348
rect -525 -438 -494 -404
rect -460 -438 -321 -404
rect -287 -438 -255 -404
rect -525 -494 -255 -438
rect -525 -528 -494 -494
rect -460 -528 -321 -494
rect -287 -528 -255 -494
rect -525 -584 -255 -528
rect -525 -618 -494 -584
rect -460 -618 -321 -584
rect -287 -618 -255 -584
rect -525 -674 -255 -618
rect -525 -708 -494 -674
rect -460 -708 -321 -674
rect -287 -708 -255 -674
rect -525 -764 -255 -708
rect -525 -798 -494 -764
rect -460 -798 -321 -764
rect -287 -798 -255 -764
rect -525 -854 -255 -798
rect -525 -888 -494 -854
rect -460 -888 -321 -854
rect -287 -888 -255 -854
rect -1714 -978 -1681 -944
rect -1647 -978 -1615 -944
rect -1714 -995 -1615 -978
rect -525 -944 -255 -888
rect -191 -64 -119 -50
rect -191 -98 -172 -64
rect -138 -98 -119 -64
rect -191 -154 -119 -98
rect 699 -79 718 -50
rect 752 -50 866 -45
rect 752 -79 771 -50
rect -191 -188 -172 -154
rect -138 -188 -119 -154
rect -191 -244 -119 -188
rect -191 -278 -172 -244
rect -138 -278 -119 -244
rect -191 -334 -119 -278
rect -191 -368 -172 -334
rect -138 -368 -119 -334
rect -191 -424 -119 -368
rect -191 -458 -172 -424
rect -138 -458 -119 -424
rect -191 -514 -119 -458
rect -191 -548 -172 -514
rect -138 -548 -119 -514
rect -191 -604 -119 -548
rect -191 -638 -172 -604
rect -138 -638 -119 -604
rect -191 -694 -119 -638
rect -191 -728 -172 -694
rect -138 -728 -119 -694
rect -191 -784 -119 -728
rect -191 -818 -172 -784
rect -138 -818 -119 -784
rect -57 -162 637 -103
rect -57 -196 2 -162
rect 36 -190 92 -162
rect 64 -196 92 -190
rect 126 -190 182 -162
rect 126 -196 130 -190
rect -57 -224 30 -196
rect 64 -224 130 -196
rect 164 -196 182 -190
rect 216 -190 272 -162
rect 216 -196 230 -190
rect 164 -224 230 -196
rect 264 -196 272 -190
rect 306 -190 362 -162
rect 396 -190 452 -162
rect 486 -190 542 -162
rect 306 -196 330 -190
rect 396 -196 430 -190
rect 486 -196 530 -190
rect 576 -196 637 -162
rect 264 -224 330 -196
rect 364 -224 430 -196
rect 464 -224 530 -196
rect 564 -224 637 -196
rect -57 -252 637 -224
rect -57 -286 2 -252
rect 36 -286 92 -252
rect 126 -286 182 -252
rect 216 -286 272 -252
rect 306 -286 362 -252
rect 396 -286 452 -252
rect 486 -286 542 -252
rect 576 -286 637 -252
rect -57 -290 637 -286
rect -57 -324 30 -290
rect 64 -324 130 -290
rect 164 -324 230 -290
rect 264 -324 330 -290
rect 364 -324 430 -290
rect 464 -324 530 -290
rect 564 -324 637 -290
rect -57 -342 637 -324
rect -57 -376 2 -342
rect 36 -376 92 -342
rect 126 -376 182 -342
rect 216 -376 272 -342
rect 306 -376 362 -342
rect 396 -376 452 -342
rect 486 -376 542 -342
rect 576 -376 637 -342
rect -57 -390 637 -376
rect -57 -424 30 -390
rect 64 -424 130 -390
rect 164 -424 230 -390
rect 264 -424 330 -390
rect 364 -424 430 -390
rect 464 -424 530 -390
rect 564 -424 637 -390
rect -57 -432 637 -424
rect -57 -466 2 -432
rect 36 -466 92 -432
rect 126 -466 182 -432
rect 216 -466 272 -432
rect 306 -466 362 -432
rect 396 -466 452 -432
rect 486 -466 542 -432
rect 576 -466 637 -432
rect -57 -490 637 -466
rect -57 -522 30 -490
rect 64 -522 130 -490
rect -57 -556 2 -522
rect 64 -524 92 -522
rect 36 -556 92 -524
rect 126 -524 130 -522
rect 164 -522 230 -490
rect 164 -524 182 -522
rect 126 -556 182 -524
rect 216 -524 230 -522
rect 264 -522 330 -490
rect 364 -522 430 -490
rect 464 -522 530 -490
rect 564 -522 637 -490
rect 264 -524 272 -522
rect 216 -556 272 -524
rect 306 -524 330 -522
rect 396 -524 430 -522
rect 486 -524 530 -522
rect 306 -556 362 -524
rect 396 -556 452 -524
rect 486 -556 542 -524
rect 576 -556 637 -522
rect -57 -590 637 -556
rect -57 -612 30 -590
rect 64 -612 130 -590
rect -57 -646 2 -612
rect 64 -624 92 -612
rect 36 -646 92 -624
rect 126 -624 130 -612
rect 164 -612 230 -590
rect 164 -624 182 -612
rect 126 -646 182 -624
rect 216 -624 230 -612
rect 264 -612 330 -590
rect 364 -612 430 -590
rect 464 -612 530 -590
rect 564 -612 637 -590
rect 264 -624 272 -612
rect 216 -646 272 -624
rect 306 -624 330 -612
rect 396 -624 430 -612
rect 486 -624 530 -612
rect 306 -646 362 -624
rect 396 -646 452 -624
rect 486 -646 542 -624
rect 576 -646 637 -612
rect -57 -690 637 -646
rect -57 -702 30 -690
rect 64 -702 130 -690
rect -57 -736 2 -702
rect 64 -724 92 -702
rect 36 -736 92 -724
rect 126 -724 130 -702
rect 164 -702 230 -690
rect 164 -724 182 -702
rect 126 -736 182 -724
rect 216 -724 230 -702
rect 264 -702 330 -690
rect 364 -702 430 -690
rect 464 -702 530 -690
rect 564 -702 637 -690
rect 264 -724 272 -702
rect 216 -736 272 -724
rect 306 -724 330 -702
rect 396 -724 430 -702
rect 486 -724 530 -702
rect 306 -736 362 -724
rect 396 -736 452 -724
rect 486 -736 542 -724
rect 576 -736 637 -702
rect -57 -797 637 -736
rect 699 -135 771 -79
rect 699 -169 718 -135
rect 752 -169 771 -135
rect 699 -225 771 -169
rect 699 -259 718 -225
rect 752 -259 771 -225
rect 699 -315 771 -259
rect 699 -349 718 -315
rect 752 -349 771 -315
rect 699 -405 771 -349
rect 699 -439 718 -405
rect 752 -439 771 -405
rect 699 -495 771 -439
rect 699 -529 718 -495
rect 752 -529 771 -495
rect 699 -585 771 -529
rect 699 -619 718 -585
rect 752 -619 771 -585
rect 699 -675 771 -619
rect 699 -709 718 -675
rect 752 -709 771 -675
rect 699 -765 771 -709
rect -191 -859 -119 -818
rect 699 -799 718 -765
rect 752 -799 771 -765
rect 699 -859 771 -799
rect -191 -878 771 -859
rect -191 -912 -80 -878
rect -46 -912 10 -878
rect 44 -912 100 -878
rect 134 -912 190 -878
rect 224 -912 280 -878
rect 314 -912 370 -878
rect 404 -912 460 -878
rect 494 -912 550 -878
rect 584 -912 640 -878
rect 674 -912 771 -878
rect -191 -931 771 -912
rect 835 -78 866 -50
rect 900 -78 1039 -44
rect 1073 -45 2226 -44
rect 1073 -50 2078 -45
rect 1073 -78 1105 -50
rect 835 -134 1105 -78
rect 835 -168 866 -134
rect 900 -168 1039 -134
rect 1073 -168 1105 -134
rect 835 -224 1105 -168
rect 835 -258 866 -224
rect 900 -258 1039 -224
rect 1073 -258 1105 -224
rect 835 -314 1105 -258
rect 835 -348 866 -314
rect 900 -348 1039 -314
rect 1073 -348 1105 -314
rect 835 -404 1105 -348
rect 835 -438 866 -404
rect 900 -438 1039 -404
rect 1073 -438 1105 -404
rect 835 -494 1105 -438
rect 835 -528 866 -494
rect 900 -528 1039 -494
rect 1073 -528 1105 -494
rect 835 -584 1105 -528
rect 835 -618 866 -584
rect 900 -618 1039 -584
rect 1073 -618 1105 -584
rect 835 -674 1105 -618
rect 835 -708 866 -674
rect 900 -708 1039 -674
rect 1073 -708 1105 -674
rect 835 -764 1105 -708
rect 835 -798 866 -764
rect 900 -798 1039 -764
rect 1073 -798 1105 -764
rect 835 -854 1105 -798
rect 835 -888 866 -854
rect 900 -888 1039 -854
rect 1073 -888 1105 -854
rect -525 -978 -494 -944
rect -460 -978 -321 -944
rect -287 -978 -255 -944
rect -525 -995 -255 -978
rect 835 -944 1105 -888
rect 1169 -64 1241 -50
rect 1169 -98 1188 -64
rect 1222 -98 1241 -64
rect 1169 -154 1241 -98
rect 2059 -79 2078 -50
rect 2112 -50 2226 -45
rect 2112 -79 2131 -50
rect 1169 -188 1188 -154
rect 1222 -188 1241 -154
rect 1169 -244 1241 -188
rect 1169 -278 1188 -244
rect 1222 -278 1241 -244
rect 1169 -334 1241 -278
rect 1169 -368 1188 -334
rect 1222 -368 1241 -334
rect 1169 -424 1241 -368
rect 1169 -458 1188 -424
rect 1222 -458 1241 -424
rect 1169 -514 1241 -458
rect 1169 -548 1188 -514
rect 1222 -548 1241 -514
rect 1169 -604 1241 -548
rect 1169 -638 1188 -604
rect 1222 -638 1241 -604
rect 1169 -694 1241 -638
rect 1169 -728 1188 -694
rect 1222 -728 1241 -694
rect 1169 -784 1241 -728
rect 1169 -818 1188 -784
rect 1222 -818 1241 -784
rect 1303 -162 1997 -103
rect 1303 -196 1362 -162
rect 1396 -190 1452 -162
rect 1424 -196 1452 -190
rect 1486 -190 1542 -162
rect 1486 -196 1490 -190
rect 1303 -224 1390 -196
rect 1424 -224 1490 -196
rect 1524 -196 1542 -190
rect 1576 -190 1632 -162
rect 1576 -196 1590 -190
rect 1524 -224 1590 -196
rect 1624 -196 1632 -190
rect 1666 -190 1722 -162
rect 1756 -190 1812 -162
rect 1846 -190 1902 -162
rect 1666 -196 1690 -190
rect 1756 -196 1790 -190
rect 1846 -196 1890 -190
rect 1936 -196 1997 -162
rect 1624 -224 1690 -196
rect 1724 -224 1790 -196
rect 1824 -224 1890 -196
rect 1924 -224 1997 -196
rect 1303 -252 1997 -224
rect 1303 -286 1362 -252
rect 1396 -286 1452 -252
rect 1486 -286 1542 -252
rect 1576 -286 1632 -252
rect 1666 -286 1722 -252
rect 1756 -286 1812 -252
rect 1846 -286 1902 -252
rect 1936 -286 1997 -252
rect 1303 -290 1997 -286
rect 1303 -324 1390 -290
rect 1424 -324 1490 -290
rect 1524 -324 1590 -290
rect 1624 -324 1690 -290
rect 1724 -324 1790 -290
rect 1824 -324 1890 -290
rect 1924 -324 1997 -290
rect 1303 -342 1997 -324
rect 1303 -376 1362 -342
rect 1396 -376 1452 -342
rect 1486 -376 1542 -342
rect 1576 -376 1632 -342
rect 1666 -376 1722 -342
rect 1756 -376 1812 -342
rect 1846 -376 1902 -342
rect 1936 -376 1997 -342
rect 1303 -390 1997 -376
rect 1303 -424 1390 -390
rect 1424 -424 1490 -390
rect 1524 -424 1590 -390
rect 1624 -424 1690 -390
rect 1724 -424 1790 -390
rect 1824 -424 1890 -390
rect 1924 -424 1997 -390
rect 1303 -432 1997 -424
rect 1303 -466 1362 -432
rect 1396 -466 1452 -432
rect 1486 -466 1542 -432
rect 1576 -466 1632 -432
rect 1666 -466 1722 -432
rect 1756 -466 1812 -432
rect 1846 -466 1902 -432
rect 1936 -466 1997 -432
rect 1303 -490 1997 -466
rect 1303 -522 1390 -490
rect 1424 -522 1490 -490
rect 1303 -556 1362 -522
rect 1424 -524 1452 -522
rect 1396 -556 1452 -524
rect 1486 -524 1490 -522
rect 1524 -522 1590 -490
rect 1524 -524 1542 -522
rect 1486 -556 1542 -524
rect 1576 -524 1590 -522
rect 1624 -522 1690 -490
rect 1724 -522 1790 -490
rect 1824 -522 1890 -490
rect 1924 -522 1997 -490
rect 1624 -524 1632 -522
rect 1576 -556 1632 -524
rect 1666 -524 1690 -522
rect 1756 -524 1790 -522
rect 1846 -524 1890 -522
rect 1666 -556 1722 -524
rect 1756 -556 1812 -524
rect 1846 -556 1902 -524
rect 1936 -556 1997 -522
rect 1303 -590 1997 -556
rect 1303 -612 1390 -590
rect 1424 -612 1490 -590
rect 1303 -646 1362 -612
rect 1424 -624 1452 -612
rect 1396 -646 1452 -624
rect 1486 -624 1490 -612
rect 1524 -612 1590 -590
rect 1524 -624 1542 -612
rect 1486 -646 1542 -624
rect 1576 -624 1590 -612
rect 1624 -612 1690 -590
rect 1724 -612 1790 -590
rect 1824 -612 1890 -590
rect 1924 -612 1997 -590
rect 1624 -624 1632 -612
rect 1576 -646 1632 -624
rect 1666 -624 1690 -612
rect 1756 -624 1790 -612
rect 1846 -624 1890 -612
rect 1666 -646 1722 -624
rect 1756 -646 1812 -624
rect 1846 -646 1902 -624
rect 1936 -646 1997 -612
rect 1303 -690 1997 -646
rect 1303 -702 1390 -690
rect 1424 -702 1490 -690
rect 1303 -736 1362 -702
rect 1424 -724 1452 -702
rect 1396 -736 1452 -724
rect 1486 -724 1490 -702
rect 1524 -702 1590 -690
rect 1524 -724 1542 -702
rect 1486 -736 1542 -724
rect 1576 -724 1590 -702
rect 1624 -702 1690 -690
rect 1724 -702 1790 -690
rect 1824 -702 1890 -690
rect 1924 -702 1997 -690
rect 1624 -724 1632 -702
rect 1576 -736 1632 -724
rect 1666 -724 1690 -702
rect 1756 -724 1790 -702
rect 1846 -724 1890 -702
rect 1666 -736 1722 -724
rect 1756 -736 1812 -724
rect 1846 -736 1902 -724
rect 1936 -736 1997 -702
rect 1303 -797 1997 -736
rect 2059 -135 2131 -79
rect 2059 -169 2078 -135
rect 2112 -169 2131 -135
rect 2059 -225 2131 -169
rect 2059 -259 2078 -225
rect 2112 -259 2131 -225
rect 2059 -315 2131 -259
rect 2059 -349 2078 -315
rect 2112 -349 2131 -315
rect 2059 -405 2131 -349
rect 2059 -439 2078 -405
rect 2112 -439 2131 -405
rect 2059 -495 2131 -439
rect 2059 -529 2078 -495
rect 2112 -529 2131 -495
rect 2059 -585 2131 -529
rect 2059 -619 2078 -585
rect 2112 -619 2131 -585
rect 2059 -675 2131 -619
rect 2059 -709 2078 -675
rect 2112 -709 2131 -675
rect 2059 -765 2131 -709
rect 1169 -859 1241 -818
rect 2059 -799 2078 -765
rect 2112 -799 2131 -765
rect 2059 -859 2131 -799
rect 1169 -878 2131 -859
rect 1169 -912 1280 -878
rect 1314 -912 1370 -878
rect 1404 -912 1460 -878
rect 1494 -912 1550 -878
rect 1584 -912 1640 -878
rect 1674 -912 1730 -878
rect 1764 -912 1820 -878
rect 1854 -912 1910 -878
rect 1944 -912 2000 -878
rect 2034 -912 2131 -878
rect 1169 -931 2131 -912
rect 2195 -78 2226 -50
rect 2260 -50 2300 -44
rect 2700 -20 2770 0
rect 2260 -78 2294 -50
rect 2195 -134 2294 -78
rect 2700 -70 2710 -20
rect 2760 -70 2770 -20
rect 2700 -90 2770 -70
rect 2195 -168 2226 -134
rect 2260 -168 2294 -134
rect 2195 -224 2294 -168
rect 2195 -258 2226 -224
rect 2260 -258 2294 -224
rect 2195 -314 2294 -258
rect 2195 -348 2226 -314
rect 2260 -348 2294 -314
rect 2195 -404 2294 -348
rect 2195 -438 2226 -404
rect 2260 -438 2294 -404
rect 2195 -494 2294 -438
rect 2195 -528 2226 -494
rect 2260 -528 2294 -494
rect 2195 -584 2294 -528
rect 2530 -160 2580 -90
rect 2195 -618 2226 -584
rect 2260 -618 2294 -584
rect 2195 -674 2294 -618
rect 2195 -708 2226 -674
rect 2260 -708 2294 -674
rect 2195 -764 2294 -708
rect 2195 -798 2226 -764
rect 2260 -798 2294 -764
rect 2195 -854 2294 -798
rect 3480 -662 3550 -640
rect 3480 -712 3490 -662
rect 3540 -712 3550 -662
rect 3480 -732 3550 -712
rect 2195 -888 2226 -854
rect 2260 -888 2294 -854
rect 835 -978 866 -944
rect 900 -978 1039 -944
rect 1073 -978 1105 -944
rect 835 -995 1105 -978
rect 2195 -944 2294 -888
rect 2195 -978 2226 -944
rect 2260 -978 2294 -944
rect 2195 -995 2294 -978
rect -1714 -1028 2294 -995
rect -1714 -1062 -1580 -1028
rect -1546 -1062 -1490 -1028
rect -1456 -1062 -1400 -1028
rect -1366 -1062 -1310 -1028
rect -1276 -1062 -1220 -1028
rect -1186 -1062 -1130 -1028
rect -1096 -1062 -1040 -1028
rect -1006 -1062 -950 -1028
rect -916 -1062 -860 -1028
rect -826 -1062 -770 -1028
rect -736 -1062 -680 -1028
rect -646 -1062 -590 -1028
rect -556 -1062 -220 -1028
rect -186 -1062 -130 -1028
rect -96 -1062 -40 -1028
rect -6 -1062 50 -1028
rect 84 -1062 140 -1028
rect 174 -1062 230 -1028
rect 264 -1062 320 -1028
rect 354 -1062 410 -1028
rect 444 -1062 500 -1028
rect 534 -1062 590 -1028
rect 624 -1062 680 -1028
rect 714 -1062 770 -1028
rect 804 -1062 1140 -1028
rect 1174 -1062 1230 -1028
rect 1264 -1062 1320 -1028
rect 1354 -1062 1410 -1028
rect 1444 -1062 1500 -1028
rect 1534 -1062 1590 -1028
rect 1624 -1062 1680 -1028
rect 1714 -1062 1770 -1028
rect 1804 -1062 1860 -1028
rect 1894 -1062 1950 -1028
rect 1984 -1062 2040 -1028
rect 2074 -1062 2130 -1028
rect 2164 -1062 2294 -1028
rect -1714 -1094 2294 -1062
rect 2820 -870 2890 -850
rect 2820 -920 2830 -870
rect 2880 -920 2890 -870
rect 2820 -940 2890 -920
rect -430 -1160 -350 -1094
rect 930 -1160 1010 -1094
rect -1720 -1201 2300 -1160
rect -1720 -1224 -1580 -1201
rect -1720 -1258 -1681 -1224
rect -1647 -1235 -1580 -1224
rect -1546 -1235 -1490 -1201
rect -1456 -1235 -1400 -1201
rect -1366 -1235 -1310 -1201
rect -1276 -1235 -1220 -1201
rect -1186 -1235 -1130 -1201
rect -1096 -1235 -1040 -1201
rect -1006 -1235 -950 -1201
rect -916 -1235 -860 -1201
rect -826 -1235 -770 -1201
rect -736 -1235 -680 -1201
rect -646 -1235 -590 -1201
rect -556 -1224 -220 -1201
rect -556 -1235 -494 -1224
rect -1647 -1258 -494 -1235
rect -460 -1258 -321 -1224
rect -287 -1235 -220 -1224
rect -186 -1235 -130 -1201
rect -96 -1235 -40 -1201
rect -6 -1235 50 -1201
rect 84 -1235 140 -1201
rect 174 -1235 230 -1201
rect 264 -1235 320 -1201
rect 354 -1235 410 -1201
rect 444 -1235 500 -1201
rect 534 -1235 590 -1201
rect 624 -1235 680 -1201
rect 714 -1235 770 -1201
rect 804 -1224 1140 -1201
rect 804 -1235 866 -1224
rect -287 -1258 866 -1235
rect 900 -1258 1039 -1224
rect 1073 -1235 1140 -1224
rect 1174 -1235 1230 -1201
rect 1264 -1235 1320 -1201
rect 1354 -1235 1410 -1201
rect 1444 -1235 1500 -1201
rect 1534 -1235 1590 -1201
rect 1624 -1235 1680 -1201
rect 1714 -1235 1770 -1201
rect 1804 -1235 1860 -1201
rect 1894 -1235 1950 -1201
rect 1984 -1235 2040 -1201
rect 2074 -1235 2130 -1201
rect 2164 -1224 2300 -1201
rect 2164 -1235 2226 -1224
rect 1073 -1258 2226 -1235
rect 2260 -1258 2300 -1224
rect -1720 -1314 2300 -1258
rect -3030 -1390 -2970 -1370
rect -3030 -1430 -3020 -1390
rect -2980 -1430 -2970 -1390
rect -3030 -1450 -2970 -1430
rect -1720 -1348 -1681 -1314
rect -1647 -1348 -494 -1314
rect -460 -1348 -321 -1314
rect -287 -1348 866 -1314
rect 900 -1348 1039 -1314
rect 1073 -1348 2226 -1314
rect 2260 -1348 2300 -1314
rect -1720 -1382 -1474 -1348
rect -1440 -1382 -1384 -1348
rect -1350 -1382 -1294 -1348
rect -1260 -1382 -1204 -1348
rect -1170 -1382 -1114 -1348
rect -1080 -1382 -1024 -1348
rect -990 -1382 -934 -1348
rect -900 -1382 -844 -1348
rect -810 -1382 -754 -1348
rect -720 -1382 -114 -1348
rect -80 -1382 -24 -1348
rect 10 -1382 66 -1348
rect 100 -1382 156 -1348
rect 190 -1382 246 -1348
rect 280 -1382 336 -1348
rect 370 -1382 426 -1348
rect 460 -1382 516 -1348
rect 550 -1382 606 -1348
rect 640 -1382 1246 -1348
rect 1280 -1382 1336 -1348
rect 1370 -1382 1426 -1348
rect 1460 -1382 1516 -1348
rect 1550 -1382 1606 -1348
rect 1640 -1382 1696 -1348
rect 1730 -1382 1786 -1348
rect 1820 -1382 1876 -1348
rect 1910 -1382 1966 -1348
rect 2000 -1382 2300 -1348
rect -1720 -1404 2300 -1382
rect -1720 -1410 -1681 -1404
rect -1714 -1438 -1681 -1410
rect -1647 -1405 -494 -1404
rect -1647 -1410 -642 -1405
rect -1647 -1438 -1615 -1410
rect -1714 -1494 -1615 -1438
rect -1714 -1528 -1681 -1494
rect -1647 -1528 -1615 -1494
rect -2860 -1798 -2790 -1778
rect -2860 -1848 -2850 -1798
rect -2800 -1848 -2790 -1798
rect -2860 -1868 -2790 -1848
rect -2670 -1988 -2620 -1918
rect -1714 -1584 -1615 -1528
rect -1714 -1618 -1681 -1584
rect -1647 -1618 -1615 -1584
rect -1714 -1674 -1615 -1618
rect -2500 -2008 -2430 -1988
rect -2500 -2058 -2490 -2008
rect -2440 -2058 -2430 -2008
rect -2500 -2078 -2430 -2058
rect -2240 -2138 -2190 -2068
rect -2070 -2158 -2000 -2138
rect -2070 -2208 -2060 -2158
rect -2010 -2208 -2000 -2158
rect -2070 -2228 -2000 -2208
rect -1714 -1708 -1681 -1674
rect -1647 -1708 -1615 -1674
rect -1714 -1764 -1615 -1708
rect -1714 -1798 -1681 -1764
rect -1647 -1798 -1615 -1764
rect -1714 -1854 -1615 -1798
rect -1714 -1888 -1681 -1854
rect -1647 -1888 -1615 -1854
rect -1714 -1944 -1615 -1888
rect -1714 -1978 -1681 -1944
rect -1647 -1978 -1615 -1944
rect -1714 -2034 -1615 -1978
rect -1714 -2068 -1681 -2034
rect -1647 -2068 -1615 -2034
rect -1714 -2124 -1615 -2068
rect -1714 -2158 -1681 -2124
rect -1647 -2158 -1615 -2124
rect -1714 -2214 -1615 -2158
rect -1714 -2248 -1681 -2214
rect -1647 -2248 -1615 -2214
rect -1714 -2304 -1615 -2248
rect -1551 -1424 -1479 -1410
rect -1551 -1458 -1532 -1424
rect -1498 -1458 -1479 -1424
rect -1551 -1514 -1479 -1458
rect -661 -1439 -642 -1410
rect -608 -1410 -494 -1405
rect -608 -1439 -589 -1410
rect -1551 -1548 -1532 -1514
rect -1498 -1548 -1479 -1514
rect -1551 -1604 -1479 -1548
rect -1551 -1638 -1532 -1604
rect -1498 -1638 -1479 -1604
rect -1551 -1694 -1479 -1638
rect -1551 -1728 -1532 -1694
rect -1498 -1728 -1479 -1694
rect -1551 -1784 -1479 -1728
rect -1551 -1818 -1532 -1784
rect -1498 -1818 -1479 -1784
rect -1551 -1874 -1479 -1818
rect -1551 -1908 -1532 -1874
rect -1498 -1908 -1479 -1874
rect -1551 -1964 -1479 -1908
rect -1551 -1998 -1532 -1964
rect -1498 -1998 -1479 -1964
rect -1551 -2054 -1479 -1998
rect -1551 -2088 -1532 -2054
rect -1498 -2088 -1479 -2054
rect -1551 -2144 -1479 -2088
rect -1551 -2178 -1532 -2144
rect -1498 -2178 -1479 -2144
rect -1417 -1522 -723 -1463
rect -1417 -1556 -1358 -1522
rect -1324 -1550 -1268 -1522
rect -1296 -1556 -1268 -1550
rect -1234 -1550 -1178 -1522
rect -1234 -1556 -1230 -1550
rect -1417 -1584 -1330 -1556
rect -1296 -1584 -1230 -1556
rect -1196 -1556 -1178 -1550
rect -1144 -1550 -1088 -1522
rect -1144 -1556 -1130 -1550
rect -1196 -1584 -1130 -1556
rect -1096 -1556 -1088 -1550
rect -1054 -1550 -998 -1522
rect -964 -1550 -908 -1522
rect -874 -1550 -818 -1522
rect -1054 -1556 -1030 -1550
rect -964 -1556 -930 -1550
rect -874 -1556 -830 -1550
rect -784 -1556 -723 -1522
rect -1096 -1584 -1030 -1556
rect -996 -1584 -930 -1556
rect -896 -1584 -830 -1556
rect -796 -1584 -723 -1556
rect -1417 -1612 -723 -1584
rect -1417 -1646 -1358 -1612
rect -1324 -1646 -1268 -1612
rect -1234 -1646 -1178 -1612
rect -1144 -1646 -1088 -1612
rect -1054 -1646 -998 -1612
rect -964 -1646 -908 -1612
rect -874 -1646 -818 -1612
rect -784 -1646 -723 -1612
rect -1417 -1650 -723 -1646
rect -1417 -1684 -1330 -1650
rect -1296 -1684 -1230 -1650
rect -1196 -1684 -1130 -1650
rect -1096 -1684 -1030 -1650
rect -996 -1684 -930 -1650
rect -896 -1684 -830 -1650
rect -796 -1684 -723 -1650
rect -1417 -1702 -723 -1684
rect -1417 -1736 -1358 -1702
rect -1324 -1736 -1268 -1702
rect -1234 -1736 -1178 -1702
rect -1144 -1736 -1088 -1702
rect -1054 -1736 -998 -1702
rect -964 -1736 -908 -1702
rect -874 -1736 -818 -1702
rect -784 -1736 -723 -1702
rect -1417 -1750 -723 -1736
rect -1417 -1784 -1330 -1750
rect -1296 -1784 -1230 -1750
rect -1196 -1784 -1130 -1750
rect -1096 -1784 -1030 -1750
rect -996 -1784 -930 -1750
rect -896 -1784 -830 -1750
rect -796 -1784 -723 -1750
rect -1417 -1792 -723 -1784
rect -1417 -1826 -1358 -1792
rect -1324 -1826 -1268 -1792
rect -1234 -1826 -1178 -1792
rect -1144 -1826 -1088 -1792
rect -1054 -1826 -998 -1792
rect -964 -1826 -908 -1792
rect -874 -1826 -818 -1792
rect -784 -1826 -723 -1792
rect -1417 -1850 -723 -1826
rect -1417 -1882 -1330 -1850
rect -1296 -1882 -1230 -1850
rect -1417 -1916 -1358 -1882
rect -1296 -1884 -1268 -1882
rect -1324 -1916 -1268 -1884
rect -1234 -1884 -1230 -1882
rect -1196 -1882 -1130 -1850
rect -1196 -1884 -1178 -1882
rect -1234 -1916 -1178 -1884
rect -1144 -1884 -1130 -1882
rect -1096 -1882 -1030 -1850
rect -996 -1882 -930 -1850
rect -896 -1882 -830 -1850
rect -796 -1882 -723 -1850
rect -1096 -1884 -1088 -1882
rect -1144 -1916 -1088 -1884
rect -1054 -1884 -1030 -1882
rect -964 -1884 -930 -1882
rect -874 -1884 -830 -1882
rect -1054 -1916 -998 -1884
rect -964 -1916 -908 -1884
rect -874 -1916 -818 -1884
rect -784 -1916 -723 -1882
rect -1417 -1950 -723 -1916
rect -1417 -1972 -1330 -1950
rect -1296 -1972 -1230 -1950
rect -1417 -2006 -1358 -1972
rect -1296 -1984 -1268 -1972
rect -1324 -2006 -1268 -1984
rect -1234 -1984 -1230 -1972
rect -1196 -1972 -1130 -1950
rect -1196 -1984 -1178 -1972
rect -1234 -2006 -1178 -1984
rect -1144 -1984 -1130 -1972
rect -1096 -1972 -1030 -1950
rect -996 -1972 -930 -1950
rect -896 -1972 -830 -1950
rect -796 -1972 -723 -1950
rect -1096 -1984 -1088 -1972
rect -1144 -2006 -1088 -1984
rect -1054 -1984 -1030 -1972
rect -964 -1984 -930 -1972
rect -874 -1984 -830 -1972
rect -1054 -2006 -998 -1984
rect -964 -2006 -908 -1984
rect -874 -2006 -818 -1984
rect -784 -2006 -723 -1972
rect -1417 -2050 -723 -2006
rect -1417 -2062 -1330 -2050
rect -1296 -2062 -1230 -2050
rect -1417 -2096 -1358 -2062
rect -1296 -2084 -1268 -2062
rect -1324 -2096 -1268 -2084
rect -1234 -2084 -1230 -2062
rect -1196 -2062 -1130 -2050
rect -1196 -2084 -1178 -2062
rect -1234 -2096 -1178 -2084
rect -1144 -2084 -1130 -2062
rect -1096 -2062 -1030 -2050
rect -996 -2062 -930 -2050
rect -896 -2062 -830 -2050
rect -796 -2062 -723 -2050
rect -1096 -2084 -1088 -2062
rect -1144 -2096 -1088 -2084
rect -1054 -2084 -1030 -2062
rect -964 -2084 -930 -2062
rect -874 -2084 -830 -2062
rect -1054 -2096 -998 -2084
rect -964 -2096 -908 -2084
rect -874 -2096 -818 -2084
rect -784 -2096 -723 -2062
rect -1417 -2157 -723 -2096
rect -661 -1495 -589 -1439
rect -661 -1529 -642 -1495
rect -608 -1529 -589 -1495
rect -661 -1585 -589 -1529
rect -661 -1619 -642 -1585
rect -608 -1619 -589 -1585
rect -661 -1675 -589 -1619
rect -661 -1709 -642 -1675
rect -608 -1709 -589 -1675
rect -661 -1765 -589 -1709
rect -661 -1799 -642 -1765
rect -608 -1799 -589 -1765
rect -661 -1855 -589 -1799
rect -661 -1889 -642 -1855
rect -608 -1889 -589 -1855
rect -661 -1945 -589 -1889
rect -661 -1979 -642 -1945
rect -608 -1979 -589 -1945
rect -661 -2035 -589 -1979
rect -661 -2069 -642 -2035
rect -608 -2069 -589 -2035
rect -661 -2125 -589 -2069
rect -1551 -2219 -1479 -2178
rect -661 -2159 -642 -2125
rect -608 -2159 -589 -2125
rect -661 -2219 -589 -2159
rect -1551 -2238 -589 -2219
rect -1551 -2272 -1440 -2238
rect -1406 -2272 -1350 -2238
rect -1316 -2272 -1260 -2238
rect -1226 -2272 -1170 -2238
rect -1136 -2272 -1080 -2238
rect -1046 -2272 -990 -2238
rect -956 -2272 -900 -2238
rect -866 -2272 -810 -2238
rect -776 -2272 -720 -2238
rect -686 -2272 -589 -2238
rect -1551 -2291 -589 -2272
rect -525 -1438 -494 -1410
rect -460 -1438 -321 -1404
rect -287 -1405 866 -1404
rect -287 -1410 718 -1405
rect -287 -1438 -255 -1410
rect -525 -1494 -255 -1438
rect -525 -1528 -494 -1494
rect -460 -1528 -321 -1494
rect -287 -1528 -255 -1494
rect -525 -1584 -255 -1528
rect -525 -1618 -494 -1584
rect -460 -1618 -321 -1584
rect -287 -1618 -255 -1584
rect -525 -1674 -255 -1618
rect -525 -1708 -494 -1674
rect -460 -1708 -321 -1674
rect -287 -1708 -255 -1674
rect -525 -1764 -255 -1708
rect -525 -1798 -494 -1764
rect -460 -1798 -321 -1764
rect -287 -1798 -255 -1764
rect -525 -1854 -255 -1798
rect -525 -1888 -494 -1854
rect -460 -1888 -321 -1854
rect -287 -1888 -255 -1854
rect -525 -1944 -255 -1888
rect -525 -1978 -494 -1944
rect -460 -1978 -321 -1944
rect -287 -1978 -255 -1944
rect -525 -2034 -255 -1978
rect -525 -2068 -494 -2034
rect -460 -2068 -321 -2034
rect -287 -2068 -255 -2034
rect -525 -2124 -255 -2068
rect -525 -2158 -494 -2124
rect -460 -2158 -321 -2124
rect -287 -2158 -255 -2124
rect -525 -2214 -255 -2158
rect -525 -2248 -494 -2214
rect -460 -2248 -321 -2214
rect -287 -2248 -255 -2214
rect -1714 -2338 -1681 -2304
rect -1647 -2338 -1615 -2304
rect -1714 -2355 -1615 -2338
rect -525 -2304 -255 -2248
rect -191 -1424 -119 -1410
rect -191 -1458 -172 -1424
rect -138 -1458 -119 -1424
rect -191 -1514 -119 -1458
rect 699 -1439 718 -1410
rect 752 -1410 866 -1405
rect 752 -1439 771 -1410
rect -191 -1548 -172 -1514
rect -138 -1548 -119 -1514
rect -191 -1604 -119 -1548
rect -191 -1638 -172 -1604
rect -138 -1638 -119 -1604
rect -191 -1694 -119 -1638
rect -191 -1728 -172 -1694
rect -138 -1728 -119 -1694
rect -191 -1784 -119 -1728
rect -191 -1818 -172 -1784
rect -138 -1818 -119 -1784
rect -191 -1874 -119 -1818
rect -191 -1908 -172 -1874
rect -138 -1908 -119 -1874
rect -191 -1964 -119 -1908
rect -191 -1998 -172 -1964
rect -138 -1998 -119 -1964
rect -191 -2054 -119 -1998
rect -191 -2088 -172 -2054
rect -138 -2088 -119 -2054
rect -191 -2144 -119 -2088
rect -191 -2178 -172 -2144
rect -138 -2178 -119 -2144
rect -57 -1522 637 -1463
rect -57 -1556 2 -1522
rect 36 -1550 92 -1522
rect 64 -1556 92 -1550
rect 126 -1550 182 -1522
rect 126 -1556 130 -1550
rect -57 -1584 30 -1556
rect 64 -1584 130 -1556
rect 164 -1556 182 -1550
rect 216 -1550 272 -1522
rect 216 -1556 230 -1550
rect 164 -1584 230 -1556
rect 264 -1556 272 -1550
rect 306 -1550 362 -1522
rect 396 -1550 452 -1522
rect 486 -1550 542 -1522
rect 306 -1556 330 -1550
rect 396 -1556 430 -1550
rect 486 -1556 530 -1550
rect 576 -1556 637 -1522
rect 264 -1584 330 -1556
rect 364 -1584 430 -1556
rect 464 -1584 530 -1556
rect 564 -1584 637 -1556
rect -57 -1612 637 -1584
rect -57 -1646 2 -1612
rect 36 -1646 92 -1612
rect 126 -1646 182 -1612
rect 216 -1646 272 -1612
rect 306 -1646 362 -1612
rect 396 -1646 452 -1612
rect 486 -1646 542 -1612
rect 576 -1646 637 -1612
rect -57 -1650 637 -1646
rect -57 -1684 30 -1650
rect 64 -1684 130 -1650
rect 164 -1684 230 -1650
rect 264 -1684 330 -1650
rect 364 -1684 430 -1650
rect 464 -1684 530 -1650
rect 564 -1684 637 -1650
rect -57 -1702 637 -1684
rect -57 -1736 2 -1702
rect 36 -1736 92 -1702
rect 126 -1736 182 -1702
rect 216 -1736 272 -1702
rect 306 -1736 362 -1702
rect 396 -1736 452 -1702
rect 486 -1736 542 -1702
rect 576 -1736 637 -1702
rect -57 -1750 637 -1736
rect -57 -1784 30 -1750
rect 64 -1784 130 -1750
rect 164 -1784 230 -1750
rect 264 -1784 330 -1750
rect 364 -1784 430 -1750
rect 464 -1784 530 -1750
rect 564 -1784 637 -1750
rect -57 -1792 637 -1784
rect -57 -1826 2 -1792
rect 36 -1826 92 -1792
rect 126 -1826 182 -1792
rect 216 -1826 272 -1792
rect 306 -1826 362 -1792
rect 396 -1826 452 -1792
rect 486 -1826 542 -1792
rect 576 -1826 637 -1792
rect -57 -1850 637 -1826
rect -57 -1882 30 -1850
rect 64 -1882 130 -1850
rect -57 -1916 2 -1882
rect 64 -1884 92 -1882
rect 36 -1916 92 -1884
rect 126 -1884 130 -1882
rect 164 -1882 230 -1850
rect 164 -1884 182 -1882
rect 126 -1916 182 -1884
rect 216 -1884 230 -1882
rect 264 -1882 330 -1850
rect 364 -1882 430 -1850
rect 464 -1882 530 -1850
rect 564 -1882 637 -1850
rect 264 -1884 272 -1882
rect 216 -1916 272 -1884
rect 306 -1884 330 -1882
rect 396 -1884 430 -1882
rect 486 -1884 530 -1882
rect 306 -1916 362 -1884
rect 396 -1916 452 -1884
rect 486 -1916 542 -1884
rect 576 -1916 637 -1882
rect -57 -1950 637 -1916
rect -57 -1972 30 -1950
rect 64 -1972 130 -1950
rect -57 -2006 2 -1972
rect 64 -1984 92 -1972
rect 36 -2006 92 -1984
rect 126 -1984 130 -1972
rect 164 -1972 230 -1950
rect 164 -1984 182 -1972
rect 126 -2006 182 -1984
rect 216 -1984 230 -1972
rect 264 -1972 330 -1950
rect 364 -1972 430 -1950
rect 464 -1972 530 -1950
rect 564 -1972 637 -1950
rect 264 -1984 272 -1972
rect 216 -2006 272 -1984
rect 306 -1984 330 -1972
rect 396 -1984 430 -1972
rect 486 -1984 530 -1972
rect 306 -2006 362 -1984
rect 396 -2006 452 -1984
rect 486 -2006 542 -1984
rect 576 -2006 637 -1972
rect -57 -2050 637 -2006
rect -57 -2062 30 -2050
rect 64 -2062 130 -2050
rect -57 -2096 2 -2062
rect 64 -2084 92 -2062
rect 36 -2096 92 -2084
rect 126 -2084 130 -2062
rect 164 -2062 230 -2050
rect 164 -2084 182 -2062
rect 126 -2096 182 -2084
rect 216 -2084 230 -2062
rect 264 -2062 330 -2050
rect 364 -2062 430 -2050
rect 464 -2062 530 -2050
rect 564 -2062 637 -2050
rect 264 -2084 272 -2062
rect 216 -2096 272 -2084
rect 306 -2084 330 -2062
rect 396 -2084 430 -2062
rect 486 -2084 530 -2062
rect 306 -2096 362 -2084
rect 396 -2096 452 -2084
rect 486 -2096 542 -2084
rect 576 -2096 637 -2062
rect -57 -2157 637 -2096
rect 699 -1495 771 -1439
rect 699 -1529 718 -1495
rect 752 -1529 771 -1495
rect 699 -1585 771 -1529
rect 699 -1619 718 -1585
rect 752 -1619 771 -1585
rect 699 -1675 771 -1619
rect 699 -1709 718 -1675
rect 752 -1709 771 -1675
rect 699 -1765 771 -1709
rect 699 -1799 718 -1765
rect 752 -1799 771 -1765
rect 699 -1855 771 -1799
rect 699 -1889 718 -1855
rect 752 -1889 771 -1855
rect 699 -1945 771 -1889
rect 699 -1979 718 -1945
rect 752 -1979 771 -1945
rect 699 -2035 771 -1979
rect 699 -2069 718 -2035
rect 752 -2069 771 -2035
rect 699 -2125 771 -2069
rect -191 -2219 -119 -2178
rect 699 -2159 718 -2125
rect 752 -2159 771 -2125
rect 699 -2219 771 -2159
rect -191 -2238 771 -2219
rect -191 -2272 -80 -2238
rect -46 -2272 10 -2238
rect 44 -2272 100 -2238
rect 134 -2272 190 -2238
rect 224 -2272 280 -2238
rect 314 -2272 370 -2238
rect 404 -2272 460 -2238
rect 494 -2272 550 -2238
rect 584 -2272 640 -2238
rect 674 -2272 771 -2238
rect -191 -2291 771 -2272
rect 835 -1438 866 -1410
rect 900 -1438 1039 -1404
rect 1073 -1405 2226 -1404
rect 1073 -1410 2078 -1405
rect 1073 -1438 1105 -1410
rect 835 -1494 1105 -1438
rect 835 -1528 866 -1494
rect 900 -1528 1039 -1494
rect 1073 -1528 1105 -1494
rect 835 -1584 1105 -1528
rect 835 -1618 866 -1584
rect 900 -1618 1039 -1584
rect 1073 -1618 1105 -1584
rect 835 -1674 1105 -1618
rect 835 -1708 866 -1674
rect 900 -1708 1039 -1674
rect 1073 -1708 1105 -1674
rect 835 -1764 1105 -1708
rect 835 -1798 866 -1764
rect 900 -1798 1039 -1764
rect 1073 -1798 1105 -1764
rect 835 -1854 1105 -1798
rect 835 -1888 866 -1854
rect 900 -1888 1039 -1854
rect 1073 -1888 1105 -1854
rect 835 -1944 1105 -1888
rect 835 -1978 866 -1944
rect 900 -1978 1039 -1944
rect 1073 -1978 1105 -1944
rect 835 -2034 1105 -1978
rect 835 -2068 866 -2034
rect 900 -2068 1039 -2034
rect 1073 -2068 1105 -2034
rect 835 -2124 1105 -2068
rect 835 -2158 866 -2124
rect 900 -2158 1039 -2124
rect 1073 -2158 1105 -2124
rect 835 -2214 1105 -2158
rect 835 -2248 866 -2214
rect 900 -2248 1039 -2214
rect 1073 -2248 1105 -2214
rect -525 -2338 -494 -2304
rect -460 -2338 -321 -2304
rect -287 -2338 -255 -2304
rect -525 -2355 -255 -2338
rect 835 -2304 1105 -2248
rect 1169 -1424 1241 -1410
rect 1169 -1458 1188 -1424
rect 1222 -1458 1241 -1424
rect 1169 -1514 1241 -1458
rect 2059 -1439 2078 -1410
rect 2112 -1410 2226 -1405
rect 2112 -1439 2131 -1410
rect 1169 -1548 1188 -1514
rect 1222 -1548 1241 -1514
rect 1169 -1604 1241 -1548
rect 1169 -1638 1188 -1604
rect 1222 -1638 1241 -1604
rect 1169 -1694 1241 -1638
rect 1169 -1728 1188 -1694
rect 1222 -1728 1241 -1694
rect 1169 -1784 1241 -1728
rect 1169 -1818 1188 -1784
rect 1222 -1818 1241 -1784
rect 1169 -1874 1241 -1818
rect 1169 -1908 1188 -1874
rect 1222 -1908 1241 -1874
rect 1169 -1964 1241 -1908
rect 1169 -1998 1188 -1964
rect 1222 -1998 1241 -1964
rect 1169 -2054 1241 -1998
rect 1169 -2088 1188 -2054
rect 1222 -2088 1241 -2054
rect 1169 -2144 1241 -2088
rect 1169 -2178 1188 -2144
rect 1222 -2178 1241 -2144
rect 1303 -1522 1997 -1463
rect 1303 -1556 1362 -1522
rect 1396 -1550 1452 -1522
rect 1424 -1556 1452 -1550
rect 1486 -1550 1542 -1522
rect 1486 -1556 1490 -1550
rect 1303 -1584 1390 -1556
rect 1424 -1584 1490 -1556
rect 1524 -1556 1542 -1550
rect 1576 -1550 1632 -1522
rect 1576 -1556 1590 -1550
rect 1524 -1584 1590 -1556
rect 1624 -1556 1632 -1550
rect 1666 -1550 1722 -1522
rect 1756 -1550 1812 -1522
rect 1846 -1550 1902 -1522
rect 1666 -1556 1690 -1550
rect 1756 -1556 1790 -1550
rect 1846 -1556 1890 -1550
rect 1936 -1556 1997 -1522
rect 1624 -1584 1690 -1556
rect 1724 -1584 1790 -1556
rect 1824 -1584 1890 -1556
rect 1924 -1584 1997 -1556
rect 1303 -1612 1997 -1584
rect 1303 -1646 1362 -1612
rect 1396 -1646 1452 -1612
rect 1486 -1646 1542 -1612
rect 1576 -1646 1632 -1612
rect 1666 -1646 1722 -1612
rect 1756 -1646 1812 -1612
rect 1846 -1646 1902 -1612
rect 1936 -1646 1997 -1612
rect 1303 -1650 1997 -1646
rect 1303 -1684 1390 -1650
rect 1424 -1684 1490 -1650
rect 1524 -1684 1590 -1650
rect 1624 -1684 1690 -1650
rect 1724 -1684 1790 -1650
rect 1824 -1684 1890 -1650
rect 1924 -1684 1997 -1650
rect 1303 -1702 1997 -1684
rect 1303 -1736 1362 -1702
rect 1396 -1736 1452 -1702
rect 1486 -1736 1542 -1702
rect 1576 -1736 1632 -1702
rect 1666 -1736 1722 -1702
rect 1756 -1736 1812 -1702
rect 1846 -1736 1902 -1702
rect 1936 -1736 1997 -1702
rect 1303 -1750 1997 -1736
rect 1303 -1784 1390 -1750
rect 1424 -1784 1490 -1750
rect 1524 -1784 1590 -1750
rect 1624 -1784 1690 -1750
rect 1724 -1784 1790 -1750
rect 1824 -1784 1890 -1750
rect 1924 -1784 1997 -1750
rect 1303 -1792 1997 -1784
rect 1303 -1826 1362 -1792
rect 1396 -1826 1452 -1792
rect 1486 -1826 1542 -1792
rect 1576 -1826 1632 -1792
rect 1666 -1826 1722 -1792
rect 1756 -1826 1812 -1792
rect 1846 -1826 1902 -1792
rect 1936 -1826 1997 -1792
rect 1303 -1850 1997 -1826
rect 1303 -1882 1390 -1850
rect 1424 -1882 1490 -1850
rect 1303 -1916 1362 -1882
rect 1424 -1884 1452 -1882
rect 1396 -1916 1452 -1884
rect 1486 -1884 1490 -1882
rect 1524 -1882 1590 -1850
rect 1524 -1884 1542 -1882
rect 1486 -1916 1542 -1884
rect 1576 -1884 1590 -1882
rect 1624 -1882 1690 -1850
rect 1724 -1882 1790 -1850
rect 1824 -1882 1890 -1850
rect 1924 -1882 1997 -1850
rect 1624 -1884 1632 -1882
rect 1576 -1916 1632 -1884
rect 1666 -1884 1690 -1882
rect 1756 -1884 1790 -1882
rect 1846 -1884 1890 -1882
rect 1666 -1916 1722 -1884
rect 1756 -1916 1812 -1884
rect 1846 -1916 1902 -1884
rect 1936 -1916 1997 -1882
rect 1303 -1950 1997 -1916
rect 1303 -1972 1390 -1950
rect 1424 -1972 1490 -1950
rect 1303 -2006 1362 -1972
rect 1424 -1984 1452 -1972
rect 1396 -2006 1452 -1984
rect 1486 -1984 1490 -1972
rect 1524 -1972 1590 -1950
rect 1524 -1984 1542 -1972
rect 1486 -2006 1542 -1984
rect 1576 -1984 1590 -1972
rect 1624 -1972 1690 -1950
rect 1724 -1972 1790 -1950
rect 1824 -1972 1890 -1950
rect 1924 -1972 1997 -1950
rect 1624 -1984 1632 -1972
rect 1576 -2006 1632 -1984
rect 1666 -1984 1690 -1972
rect 1756 -1984 1790 -1972
rect 1846 -1984 1890 -1972
rect 1666 -2006 1722 -1984
rect 1756 -2006 1812 -1984
rect 1846 -2006 1902 -1984
rect 1936 -2006 1997 -1972
rect 1303 -2050 1997 -2006
rect 1303 -2062 1390 -2050
rect 1424 -2062 1490 -2050
rect 1303 -2096 1362 -2062
rect 1424 -2084 1452 -2062
rect 1396 -2096 1452 -2084
rect 1486 -2084 1490 -2062
rect 1524 -2062 1590 -2050
rect 1524 -2084 1542 -2062
rect 1486 -2096 1542 -2084
rect 1576 -2084 1590 -2062
rect 1624 -2062 1690 -2050
rect 1724 -2062 1790 -2050
rect 1824 -2062 1890 -2050
rect 1924 -2062 1997 -2050
rect 1624 -2084 1632 -2062
rect 1576 -2096 1632 -2084
rect 1666 -2084 1690 -2062
rect 1756 -2084 1790 -2062
rect 1846 -2084 1890 -2062
rect 1666 -2096 1722 -2084
rect 1756 -2096 1812 -2084
rect 1846 -2096 1902 -2084
rect 1936 -2096 1997 -2062
rect 1303 -2157 1997 -2096
rect 2059 -1495 2131 -1439
rect 2059 -1529 2078 -1495
rect 2112 -1529 2131 -1495
rect 2059 -1585 2131 -1529
rect 2059 -1619 2078 -1585
rect 2112 -1619 2131 -1585
rect 2059 -1675 2131 -1619
rect 2059 -1709 2078 -1675
rect 2112 -1709 2131 -1675
rect 2059 -1765 2131 -1709
rect 2059 -1799 2078 -1765
rect 2112 -1799 2131 -1765
rect 2059 -1855 2131 -1799
rect 2059 -1889 2078 -1855
rect 2112 -1889 2131 -1855
rect 2059 -1945 2131 -1889
rect 2059 -1979 2078 -1945
rect 2112 -1979 2131 -1945
rect 2059 -2035 2131 -1979
rect 2059 -2069 2078 -2035
rect 2112 -2069 2131 -2035
rect 2059 -2125 2131 -2069
rect 1169 -2219 1241 -2178
rect 2059 -2159 2078 -2125
rect 2112 -2159 2131 -2125
rect 2059 -2219 2131 -2159
rect 1169 -2238 2131 -2219
rect 1169 -2272 1280 -2238
rect 1314 -2272 1370 -2238
rect 1404 -2272 1460 -2238
rect 1494 -2272 1550 -2238
rect 1584 -2272 1640 -2238
rect 1674 -2272 1730 -2238
rect 1764 -2272 1820 -2238
rect 1854 -2272 1910 -2238
rect 1944 -2272 2000 -2238
rect 2034 -2272 2131 -2238
rect 1169 -2291 2131 -2272
rect 2195 -1438 2226 -1410
rect 2260 -1410 2300 -1404
rect 2260 -1438 2294 -1410
rect 2195 -1494 2294 -1438
rect 2195 -1528 2226 -1494
rect 2260 -1528 2294 -1494
rect 3000 -1450 3060 -1430
rect 3000 -1490 3010 -1450
rect 3050 -1490 3060 -1450
rect 3000 -1510 3060 -1490
rect 2195 -1584 2294 -1528
rect 2195 -1618 2226 -1584
rect 2260 -1618 2294 -1584
rect 2195 -1674 2294 -1618
rect 2195 -1708 2226 -1674
rect 2260 -1708 2294 -1674
rect 2195 -1764 2294 -1708
rect 2195 -1798 2226 -1764
rect 2260 -1798 2294 -1764
rect 2195 -1854 2294 -1798
rect 2195 -1888 2226 -1854
rect 2260 -1888 2294 -1854
rect 2195 -1944 2294 -1888
rect 2195 -1978 2226 -1944
rect 2260 -1978 2294 -1944
rect 2195 -2034 2294 -1978
rect 2195 -2068 2226 -2034
rect 2260 -2068 2294 -2034
rect 2195 -2124 2294 -2068
rect 2195 -2158 2226 -2124
rect 2260 -2158 2294 -2124
rect 2195 -2214 2294 -2158
rect 2195 -2248 2226 -2214
rect 2260 -2248 2294 -2214
rect 2650 -2138 2700 -2068
rect 2820 -2008 2890 -1988
rect 2820 -2058 2830 -2008
rect 2880 -2058 2890 -2008
rect 2820 -2078 2890 -2058
rect 3480 -2008 3550 -1988
rect 3480 -2058 3490 -2008
rect 3540 -2058 3550 -2008
rect 3480 -2078 3550 -2058
rect 2460 -2158 2530 -2138
rect 2460 -2208 2470 -2158
rect 2520 -2208 2530 -2158
rect 2460 -2228 2530 -2208
rect 835 -2338 866 -2304
rect 900 -2338 1039 -2304
rect 1073 -2338 1105 -2304
rect 835 -2355 1105 -2338
rect 2195 -2304 2294 -2248
rect 2195 -2338 2226 -2304
rect 2260 -2338 2294 -2304
rect 2195 -2355 2294 -2338
rect -1714 -2388 2294 -2355
rect -1714 -2422 -1580 -2388
rect -1546 -2422 -1490 -2388
rect -1456 -2422 -1400 -2388
rect -1366 -2422 -1310 -2388
rect -1276 -2422 -1220 -2388
rect -1186 -2422 -1130 -2388
rect -1096 -2422 -1040 -2388
rect -1006 -2422 -950 -2388
rect -916 -2422 -860 -2388
rect -826 -2422 -770 -2388
rect -736 -2422 -680 -2388
rect -646 -2422 -590 -2388
rect -556 -2422 -220 -2388
rect -186 -2422 -130 -2388
rect -96 -2422 -40 -2388
rect -6 -2422 50 -2388
rect 84 -2422 140 -2388
rect 174 -2422 230 -2388
rect 264 -2422 320 -2388
rect 354 -2422 410 -2388
rect 444 -2422 500 -2388
rect 534 -2422 590 -2388
rect 624 -2422 680 -2388
rect 714 -2422 770 -2388
rect 804 -2422 1140 -2388
rect 1174 -2422 1230 -2388
rect 1264 -2422 1320 -2388
rect 1354 -2422 1410 -2388
rect 1444 -2422 1500 -2388
rect 1534 -2422 1590 -2388
rect 1624 -2422 1680 -2388
rect 1714 -2422 1770 -2388
rect 1804 -2422 1860 -2388
rect 1894 -2422 1950 -2388
rect 1984 -2422 2040 -2388
rect 2074 -2422 2130 -2388
rect 2164 -2422 2294 -2388
rect -1714 -2454 2294 -2422
rect -430 -2460 -350 -2454
rect 250 -2540 330 -2454
rect 930 -2460 1010 -2454
rect 250 -2580 270 -2540
rect 310 -2580 330 -2540
rect 250 -2620 330 -2580
rect 250 -2660 270 -2620
rect 310 -2660 330 -2620
rect 250 -2700 330 -2660
rect 250 -2740 270 -2700
rect 310 -2740 330 -2700
rect 250 -2760 330 -2740
rect 2890 -2910 2970 -2900
rect 5340 -2910 5420 -2900
rect 2890 -2920 2978 -2910
rect 2890 -2960 2910 -2920
rect 2950 -2960 2978 -2920
rect 2890 -2980 2978 -2960
rect 5330 -2920 5420 -2910
rect 5330 -2960 5360 -2920
rect 5400 -2960 5420 -2920
rect 5330 -2980 5420 -2960
<< viali >>
rect 9430 13850 9470 13890
rect 9950 13850 9990 13890
rect 10470 13850 10510 13890
rect 10960 13850 11000 13890
rect 9320 13720 9360 13760
rect 9320 13620 9360 13660
rect 9430 13720 9470 13760
rect 9430 13620 9470 13660
rect 9840 13720 9880 13760
rect 9840 13620 9880 13660
rect 9950 13720 9990 13760
rect 9950 13620 9990 13660
rect 10360 13720 10400 13760
rect 10360 13620 10400 13660
rect 10470 13720 10510 13760
rect 10470 13620 10510 13660
rect 10960 13720 11000 13760
rect 10960 13620 11000 13660
rect 11070 13720 11110 13760
rect 11070 13620 11110 13660
rect 9378 13508 9412 13542
rect 9898 13508 9932 13542
rect 10418 13508 10452 13542
rect 10986 13508 11020 13542
rect 9320 13340 9360 13380
rect 9320 13240 9360 13280
rect 9430 13340 9470 13380
rect 9430 13240 9470 13280
rect 9840 13340 9880 13380
rect 9840 13240 9880 13280
rect 9950 13340 9990 13380
rect 9950 13240 9990 13280
rect 10360 13340 10400 13380
rect 10360 13240 10400 13280
rect 10470 13340 10510 13380
rect 10470 13240 10510 13280
rect -1330 13000 -1290 13040
rect -1110 13000 -1070 13040
rect -640 13000 -600 13040
rect -300 13000 -260 13040
rect -80 13000 -40 13040
rect 360 13000 400 13040
rect 1040 13000 1080 13040
rect 1260 13000 1300 13040
rect 1730 13000 1770 13040
rect 2190 13000 2230 13040
rect 2540 13000 2580 13040
rect 2790 13000 2830 13040
rect 3010 13000 3050 13040
rect 3340 13000 3380 13040
rect 4000 13000 4040 13040
rect 4220 13000 4260 13040
rect 4790 13000 4830 13040
rect 5050 13000 5090 13040
rect 5300 13000 5340 13040
rect 5520 13000 5560 13040
rect 6070 13000 6110 13040
rect 6350 13000 6390 13040
rect 6600 13000 6640 13040
rect 6820 13000 6860 13040
rect 7370 13000 7410 13040
rect 7650 13000 7690 13040
rect 7900 13000 7940 13040
rect 8120 13000 8160 13040
rect 8670 13000 8710 13040
rect -1490 12890 -1450 12930
rect -540 12870 -500 12910
rect -410 12880 -370 12920
rect 530 12880 570 12920
rect 2090 12880 2130 12920
rect 4694 12890 4734 12930
rect -1550 12620 -1510 12660
rect 120 12650 160 12690
rect 640 12650 680 12690
rect 860 12450 900 12490
rect 2360 12640 2400 12680
rect 9392 13128 9426 13162
rect 9912 13128 9946 13162
rect 10432 13128 10466 13162
rect 9320 12960 9360 13000
rect 9430 12960 9470 13000
rect 9840 12960 9880 13000
rect 9950 12960 9990 13000
rect 10360 12960 10400 13000
rect 10470 12960 10510 13000
rect 9364 12848 9398 12882
rect 9884 12848 9918 12882
rect 10404 12848 10438 12882
rect 8874 12628 8908 12662
rect -850 12330 -810 12370
rect -660 12330 -620 12370
rect -540 12350 -500 12390
rect 270 12330 310 12370
rect 400 12330 440 12370
rect 1530 12330 1570 12370
rect 1750 12330 1790 12370
rect 2880 12320 2920 12360
rect 3290 12320 3330 12360
rect 5240 12330 5280 12370
rect 5820 12330 5860 12370
rect 6540 12330 6580 12370
rect 7120 12330 7160 12370
rect 7840 12330 7880 12370
rect 8420 12330 8460 12370
rect -1170 12220 -1130 12260
rect -750 12220 -710 12260
rect -80 12220 -40 12260
rect 490 12220 530 12260
rect 1200 12220 1240 12260
rect 1630 12220 1670 12260
rect 2070 12220 2110 12260
rect 2320 12220 2360 12260
rect 2540 12220 2580 12260
rect 3010 12220 3050 12260
rect 3450 12220 3490 12260
rect 4070 12220 4110 12260
rect 4410 12220 4450 12260
rect 4770 12220 4810 12260
rect 5370 12220 5410 12260
rect 5710 12220 5750 12260
rect 6070 12220 6110 12260
rect 6670 12220 6710 12260
rect 7010 12220 7050 12260
rect 7370 12220 7410 12260
rect 7970 12220 8010 12260
rect 8310 12220 8350 12260
rect 8670 12220 8710 12260
rect 9364 12418 9398 12452
rect 9884 12418 9918 12452
rect 10404 12418 10438 12452
rect 9320 12300 9360 12340
rect 9320 12200 9360 12240
rect 9430 12300 9470 12340
rect 9430 12200 9470 12240
rect 9840 12300 9880 12340
rect 9840 12200 9880 12240
rect 9950 12300 9990 12340
rect 9950 12200 9990 12240
rect 10360 12300 10400 12340
rect 10360 12200 10400 12240
rect 10470 12300 10510 12340
rect 10470 12200 10510 12240
rect 9392 12038 9426 12072
rect 9912 12038 9946 12072
rect 10432 12038 10466 12072
rect 9320 11920 9360 11960
rect 9320 11820 9360 11860
rect 9320 11720 9360 11760
rect 9320 11620 9360 11660
rect 9430 11920 9470 11960
rect 9430 11820 9470 11860
rect 9430 11720 9470 11760
rect 9430 11620 9470 11660
rect 9840 11920 9880 11960
rect 9840 11820 9880 11860
rect 9840 11720 9880 11760
rect 9840 11620 9880 11660
rect 9950 11920 9990 11960
rect 9950 11820 9990 11860
rect 9950 11720 9990 11760
rect 9950 11620 9990 11660
rect 10360 11920 10400 11960
rect 10360 11820 10400 11860
rect 10360 11720 10400 11760
rect 10360 11620 10400 11660
rect 10470 11920 10510 11960
rect 10470 11820 10510 11860
rect 10470 11720 10510 11760
rect 10470 11620 10510 11660
rect 9510 11350 9550 11390
rect 10030 11350 10070 11390
rect 10550 11350 10590 11390
rect 11070 11350 11110 11390
rect 9320 11230 9360 11270
rect 9320 11130 9360 11170
rect 9320 11030 9360 11070
rect 9320 10930 9360 10970
rect 9700 11230 9740 11270
rect 9700 11130 9740 11170
rect 9700 11030 9740 11070
rect 9700 10930 9740 10970
rect 9840 11230 9880 11270
rect 9840 11130 9880 11170
rect 9840 11030 9880 11070
rect 9840 10930 9880 10970
rect 10220 11230 10260 11270
rect 10220 11130 10260 11170
rect 10220 11030 10260 11070
rect 10220 10930 10260 10970
rect 10360 11230 10400 11270
rect 10360 11130 10400 11170
rect 10360 11030 10400 11070
rect 10360 10930 10400 10970
rect 10740 11230 10780 11270
rect 10740 11130 10780 11170
rect 10740 11030 10780 11070
rect 10740 10930 10780 10970
rect 10880 11230 10920 11270
rect 10880 11130 10920 11170
rect 10880 11030 10920 11070
rect 10880 10930 10920 10970
rect 11260 11230 11300 11270
rect 11260 11130 11300 11170
rect 11260 11030 11300 11070
rect 11260 10930 11300 10970
rect 9700 10800 9740 10840
rect 10220 10800 10260 10840
rect 10740 10800 10780 10840
rect 11260 10800 11300 10840
rect -620 10400 -580 10440
rect -400 10400 -360 10440
rect -100 10400 -60 10440
rect 120 10400 160 10440
rect 280 10400 320 10440
rect 500 10400 540 10440
rect 800 10400 840 10440
rect 1020 10400 1060 10440
rect 1320 10400 1360 10440
rect 1760 10400 1800 10440
rect 2090 10400 2130 10440
rect 2520 10400 2560 10440
rect 2910 10400 2950 10440
rect 3300 10400 3340 10440
rect 9110 10450 9180 10520
rect -210 10290 -170 10330
rect -740 9910 -700 9950
rect 1510 10290 1550 10330
rect 3590 10290 3630 10330
rect 1160 9940 1200 9980
rect 2250 9900 2290 9940
rect 2380 9930 2420 9970
rect 4130 9950 4170 9990
rect 3820 9870 3860 9910
rect 5670 9840 5710 9880
rect 8510 9840 8550 9880
rect 5670 9720 5710 9760
rect 5670 9620 5710 9660
rect 5670 9520 5710 9560
rect 1380 9330 1420 9370
rect 5670 9420 5710 9460
rect 5890 9720 5930 9760
rect 5890 9620 5930 9660
rect 5890 9520 5930 9560
rect 5890 9420 5930 9460
rect 6110 9720 6150 9760
rect 6110 9620 6150 9660
rect 6110 9520 6150 9560
rect 6110 9420 6150 9460
rect 6330 9720 6370 9760
rect 6330 9620 6370 9660
rect 6330 9520 6370 9560
rect 6330 9420 6370 9460
rect 6550 9720 6590 9760
rect 6550 9620 6590 9660
rect 6550 9520 6590 9560
rect 6550 9420 6590 9460
rect 6770 9720 6810 9760
rect 6770 9620 6810 9660
rect 6770 9520 6810 9560
rect 6770 9420 6810 9460
rect 6990 9720 7030 9760
rect 7090 9720 7130 9760
rect 7190 9720 7230 9760
rect 6990 9620 7030 9660
rect 7090 9620 7130 9660
rect 7190 9620 7230 9660
rect 6990 9520 7030 9560
rect 7090 9520 7130 9560
rect 7190 9520 7230 9560
rect 6990 9420 7030 9460
rect 7090 9420 7130 9460
rect 7190 9420 7230 9460
rect 7410 9720 7450 9760
rect 7410 9620 7450 9660
rect 7410 9520 7450 9560
rect 7410 9420 7450 9460
rect 7630 9720 7670 9760
rect 7630 9620 7670 9660
rect 7630 9520 7670 9560
rect 7630 9420 7670 9460
rect 7850 9720 7890 9760
rect 7850 9620 7890 9660
rect 7850 9520 7890 9560
rect 7850 9420 7890 9460
rect 8070 9720 8110 9760
rect 8070 9620 8110 9660
rect 8070 9520 8110 9560
rect 8070 9420 8110 9460
rect 8290 9720 8330 9760
rect 8290 9620 8330 9660
rect 8290 9520 8330 9560
rect 8290 9420 8330 9460
rect 8510 9720 8550 9760
rect 8510 9620 8550 9660
rect 8510 9520 8550 9560
rect 8510 9420 8550 9460
rect 6330 9300 6370 9340
rect -620 9220 -580 9260
rect 120 9220 160 9260
rect 280 9220 320 9260
rect 1020 9220 1060 9260
rect 1270 9220 1310 9260
rect 1460 9220 1500 9260
rect 1540 9220 1580 9260
rect 1750 9220 1790 9260
rect 2080 9220 2120 9260
rect 2520 9220 2560 9260
rect 2910 9220 2950 9260
rect 3300 9220 3340 9260
rect 3980 9220 4020 9260
rect 7500 9270 7540 9310
rect 8200 9270 8240 9310
rect 8870 9270 8940 9340
rect -170 9110 -130 9150
rect 2950 9110 2990 9150
rect 3590 9110 3630 9150
rect -740 8530 -700 8570
rect 5910 8730 5950 8770
rect 1180 8540 1220 8580
rect 2210 8540 2250 8580
rect 2360 8530 2400 8570
rect 5470 8620 5510 8660
rect 4130 8490 4170 8530
rect 5470 8520 5510 8560
rect 5470 8420 5510 8460
rect 5470 8320 5510 8360
rect 5690 8620 5730 8660
rect 5690 8520 5730 8560
rect 5690 8420 5730 8460
rect 5690 8320 5730 8360
rect 7940 8770 7980 8810
rect 8200 8770 8240 8810
rect 8870 8740 8940 8810
rect 5910 8620 5950 8660
rect 5910 8520 5950 8560
rect 5910 8420 5950 8460
rect 5910 8320 5950 8360
rect 6130 8620 6170 8660
rect 6130 8520 6170 8560
rect 6130 8420 6170 8460
rect 6130 8320 6170 8360
rect 6350 8620 6390 8660
rect 6450 8620 6490 8660
rect 6550 8620 6590 8660
rect 6350 8520 6390 8560
rect 6450 8520 6490 8560
rect 6550 8520 6590 8560
rect 6350 8420 6390 8460
rect 6450 8420 6490 8460
rect 6550 8420 6590 8460
rect 6350 8320 6390 8360
rect 6450 8320 6490 8360
rect 6550 8320 6590 8360
rect 6770 8620 6810 8660
rect 6770 8520 6810 8560
rect 6770 8420 6810 8460
rect 6770 8320 6810 8360
rect 6990 8620 7030 8660
rect 6990 8520 7030 8560
rect 6990 8420 7030 8460
rect 6990 8320 7030 8360
rect 7210 8620 7250 8660
rect 7210 8520 7250 8560
rect 7210 8420 7250 8460
rect 7210 8320 7250 8360
rect 7430 8620 7470 8660
rect 7530 8620 7570 8660
rect 7630 8620 7670 8660
rect 7430 8520 7470 8560
rect 7530 8520 7570 8560
rect 7630 8520 7670 8560
rect 7430 8420 7470 8460
rect 7530 8420 7570 8460
rect 7630 8420 7670 8460
rect 7430 8320 7470 8360
rect 7530 8320 7570 8360
rect 7630 8320 7670 8360
rect 7850 8620 7890 8660
rect 7850 8520 7890 8560
rect 7850 8420 7890 8460
rect 7850 8320 7890 8360
rect 8070 8620 8110 8660
rect 8070 8520 8110 8560
rect 8070 8420 8110 8460
rect 8070 8320 8110 8360
rect 8290 8620 8330 8660
rect 8290 8520 8330 8560
rect 8290 8420 8330 8460
rect 8290 8320 8330 8360
rect 8510 8620 8550 8660
rect 8510 8520 8550 8560
rect 8510 8420 8550 8460
rect 8510 8320 8550 8360
rect 3030 8150 3070 8190
rect 3660 8150 3700 8190
rect 5470 8200 5510 8240
rect 8510 8200 8550 8240
rect -620 8040 -580 8080
rect -400 8040 -360 8080
rect -100 8040 -60 8080
rect 130 8040 170 8080
rect 280 8040 320 8080
rect 500 8040 540 8080
rect 800 8040 840 8080
rect 1020 8040 1060 8080
rect 1420 8040 1460 8080
rect 1750 8040 1790 8080
rect 2080 8040 2120 8080
rect 2520 8040 2560 8080
rect 3300 8040 3340 8080
rect 3980 8040 4020 8080
rect 9220 7950 9290 8020
rect 9340 7200 9400 7260
rect -1340 6920 -1300 6960
rect -20 6920 20 6960
rect 560 6920 600 6960
rect 1880 6920 1920 6960
rect -1420 6800 -1380 6840
rect -1340 6800 -1300 6840
rect -1420 6700 -1380 6740
rect -1340 6700 -1300 6740
rect -1230 6800 -1190 6840
rect -1230 6700 -1190 6740
rect -1120 6800 -1080 6840
rect -1120 6700 -1080 6740
rect -1010 6800 -970 6840
rect -1010 6700 -970 6740
rect -900 6800 -860 6840
rect -900 6700 -860 6740
rect -790 6800 -750 6840
rect -790 6700 -750 6740
rect -680 6800 -640 6840
rect -680 6700 -640 6740
rect -570 6800 -530 6840
rect -570 6700 -530 6740
rect -460 6800 -420 6840
rect -460 6700 -420 6740
rect -350 6800 -310 6840
rect -350 6700 -310 6740
rect -240 6800 -200 6840
rect -240 6700 -200 6740
rect -130 6800 -90 6840
rect -130 6700 -90 6740
rect -20 6800 20 6840
rect 60 6800 100 6840
rect -20 6700 20 6740
rect 60 6700 100 6740
rect 480 6800 520 6840
rect 560 6800 600 6840
rect 480 6700 520 6740
rect 560 6700 600 6740
rect 670 6800 710 6840
rect 670 6700 710 6740
rect 780 6800 820 6840
rect 780 6700 820 6740
rect 890 6800 930 6840
rect 890 6700 930 6740
rect 1000 6800 1040 6840
rect 1000 6700 1040 6740
rect 1110 6800 1150 6840
rect 1110 6700 1150 6740
rect 1220 6800 1260 6840
rect 1220 6700 1260 6740
rect 1330 6800 1370 6840
rect 1330 6700 1370 6740
rect 1440 6800 1480 6840
rect 1440 6700 1480 6740
rect 1550 6800 1590 6840
rect 1550 6700 1590 6740
rect 1660 6800 1700 6840
rect 1660 6700 1700 6740
rect 1770 6800 1810 6840
rect 1770 6700 1810 6740
rect 1880 6800 1920 6840
rect 1960 6800 2000 6840
rect 1880 6700 1920 6740
rect 1960 6700 2000 6740
rect 9140 6690 9180 6730
rect -1172 6588 -1138 6622
rect -1062 6588 -1028 6622
rect -952 6588 -918 6622
rect -842 6588 -808 6622
rect -732 6588 -698 6622
rect -622 6588 -588 6622
rect -512 6588 -478 6622
rect -402 6588 -368 6622
rect -292 6588 -258 6622
rect -182 6588 -148 6622
rect 728 6588 762 6622
rect 838 6588 872 6622
rect 948 6588 982 6622
rect 1058 6588 1092 6622
rect 1168 6588 1202 6622
rect 1278 6588 1312 6622
rect 1388 6588 1422 6622
rect 1498 6588 1532 6622
rect 1608 6588 1642 6622
rect 1718 6588 1752 6622
rect -1350 6320 -1310 6360
rect -990 6320 -950 6360
rect -630 6320 -590 6360
rect -270 6320 -230 6360
rect 90 6320 130 6360
rect 450 6320 490 6360
rect 810 6320 850 6360
rect 1170 6320 1210 6360
rect 1530 6320 1570 6360
rect 1890 6320 1930 6360
rect 5270 6300 5310 6340
rect -1350 6200 -1310 6240
rect -1350 6100 -1310 6140
rect -1350 6000 -1310 6040
rect -1350 5900 -1310 5940
rect -1350 5800 -1310 5840
rect -1350 5700 -1310 5740
rect -1170 6200 -1130 6240
rect -1170 6100 -1130 6140
rect -1170 6000 -1130 6040
rect -1170 5900 -1130 5940
rect -1170 5800 -1130 5840
rect -1170 5700 -1130 5740
rect -990 6200 -950 6240
rect -990 6100 -950 6140
rect -990 6000 -950 6040
rect -990 5900 -950 5940
rect -990 5800 -950 5840
rect -990 5700 -950 5740
rect -810 6200 -770 6240
rect -810 6100 -770 6140
rect -810 6000 -770 6040
rect -810 5900 -770 5940
rect -810 5800 -770 5840
rect -810 5700 -770 5740
rect -630 6200 -590 6240
rect -630 6100 -590 6140
rect -630 6000 -590 6040
rect -630 5900 -590 5940
rect -630 5800 -590 5840
rect -630 5700 -590 5740
rect -450 6200 -410 6240
rect -450 6100 -410 6140
rect -450 6000 -410 6040
rect -450 5900 -410 5940
rect -450 5800 -410 5840
rect -450 5700 -410 5740
rect -270 6200 -230 6240
rect -270 6100 -230 6140
rect -270 6000 -230 6040
rect -270 5900 -230 5940
rect -270 5800 -230 5840
rect -270 5700 -230 5740
rect -90 6200 -50 6240
rect -90 6100 -50 6140
rect -90 6000 -50 6040
rect -90 5900 -50 5940
rect -90 5800 -50 5840
rect -90 5700 -50 5740
rect 90 6200 130 6240
rect 90 6100 130 6140
rect 90 6000 130 6040
rect 90 5900 130 5940
rect 90 5800 130 5840
rect 90 5700 130 5740
rect 270 6200 310 6240
rect 270 6100 310 6140
rect 270 6000 310 6040
rect 270 5900 310 5940
rect 270 5800 310 5840
rect 270 5700 310 5740
rect 450 6200 490 6240
rect 450 6100 490 6140
rect 450 6000 490 6040
rect 450 5900 490 5940
rect 450 5800 490 5840
rect 450 5700 490 5740
rect 630 6200 670 6240
rect 630 6100 670 6140
rect 630 6000 670 6040
rect 630 5900 670 5940
rect 630 5800 670 5840
rect 630 5700 670 5740
rect 810 6200 850 6240
rect 810 6100 850 6140
rect 810 6000 850 6040
rect 810 5900 850 5940
rect 810 5800 850 5840
rect 810 5700 850 5740
rect 990 6200 1030 6240
rect 990 6100 1030 6140
rect 990 6000 1030 6040
rect 990 5900 1030 5940
rect 990 5800 1030 5840
rect 990 5700 1030 5740
rect 1170 6200 1210 6240
rect 1170 6100 1210 6140
rect 1170 6000 1210 6040
rect 1170 5900 1210 5940
rect 1170 5800 1210 5840
rect 1170 5700 1210 5740
rect 1350 6200 1390 6240
rect 1350 6100 1390 6140
rect 1350 6000 1390 6040
rect 1350 5900 1390 5940
rect 1350 5800 1390 5840
rect 1350 5700 1390 5740
rect 1530 6200 1570 6240
rect 1530 6100 1570 6140
rect 1530 6000 1570 6040
rect 1530 5900 1570 5940
rect 1530 5800 1570 5840
rect 1530 5700 1570 5740
rect 1710 6200 1750 6240
rect 1710 6100 1750 6140
rect 1710 6000 1750 6040
rect 1710 5900 1750 5940
rect 1710 5800 1750 5840
rect 1710 5700 1750 5740
rect 1890 6200 1930 6240
rect 1890 6100 1930 6140
rect 2520 6120 2560 6160
rect 2740 6120 2780 6160
rect 2960 6120 3000 6160
rect 1890 6000 1930 6040
rect 1890 5900 1930 5940
rect 2520 6000 2560 6040
rect 2520 5900 2560 5940
rect 2630 6000 2670 6040
rect 2630 5900 2670 5940
rect 2740 6000 2780 6040
rect 2740 5900 2780 5940
rect 2850 6000 2890 6040
rect 2850 5900 2890 5940
rect 2960 6000 3000 6040
rect 2960 5900 3000 5940
rect 1890 5800 1930 5840
rect 2620 5780 2660 5820
rect 2740 5780 2780 5820
rect 5730 5980 5770 6030
rect 5730 5840 5770 5890
rect 6130 5980 6170 6030
rect 6130 5840 6170 5890
rect 6530 5980 6570 6030
rect 6530 5840 6570 5890
rect 6930 5980 6970 6030
rect 6930 5840 6970 5890
rect 7330 5980 7370 6030
rect 7330 5840 7370 5890
rect 2860 5780 2900 5820
rect 1890 5700 1930 5740
rect 5530 5720 5570 5760
rect 7110 5680 7150 5720
rect 7530 5720 7570 5760
rect -1080 5580 -1040 5620
rect -900 5580 -860 5620
rect -720 5580 -680 5620
rect -540 5580 -500 5620
rect -360 5580 -320 5620
rect -180 5580 -140 5620
rect 0 5580 40 5620
rect 180 5580 220 5620
rect 360 5580 400 5620
rect 540 5580 580 5620
rect 720 5580 760 5620
rect 900 5580 940 5620
rect 1080 5580 1120 5620
rect 1260 5580 1300 5620
rect 1440 5580 1480 5620
rect 1620 5580 1660 5620
rect 5970 5570 6010 5610
rect 8250 5570 8290 5610
rect 7110 5460 7150 5500
rect 5580 5300 5620 5340
rect 5710 5300 5750 5340
rect 5840 5300 5880 5340
rect 5970 5300 6010 5340
rect 6100 5300 6140 5340
rect 6230 5300 6270 5340
rect 6360 5300 6400 5340
rect 6720 5300 6760 5340
rect 6850 5300 6890 5340
rect 6980 5300 7020 5340
rect 7110 5300 7150 5340
rect 7240 5300 7280 5340
rect 7370 5300 7410 5340
rect 7500 5300 7540 5340
rect 5840 5180 5880 5220
rect 6890 5180 6930 5220
rect 7330 5180 7370 5220
rect 9570 5260 9640 5330
rect 8870 5180 8910 5220
rect 8030 5060 8070 5100
rect 9740 5010 9780 5050
rect 5750 4840 5790 4880
rect 6190 4840 6230 4880
rect 6980 4850 7020 4890
rect 8030 4840 8070 4880
rect -2450 4760 -2410 4800
rect -50 4760 -10 4800
rect 590 4760 630 4800
rect 2990 4760 3030 4800
rect 8870 4840 8910 4880
rect 5580 4720 5620 4760
rect -2450 4640 -2410 4680
rect -2450 4540 -2410 4580
rect -2330 4640 -2290 4680
rect -2330 4540 -2290 4580
rect -2210 4640 -2170 4680
rect -2210 4540 -2170 4580
rect -2090 4640 -2050 4680
rect -2090 4540 -2050 4580
rect -1970 4640 -1930 4680
rect -1970 4540 -1930 4580
rect -1850 4640 -1810 4680
rect -1850 4540 -1810 4580
rect -1730 4640 -1690 4680
rect -1730 4540 -1690 4580
rect -1610 4640 -1570 4680
rect -1610 4540 -1570 4580
rect -1490 4640 -1450 4680
rect -1490 4540 -1450 4580
rect -1370 4640 -1330 4680
rect -1370 4540 -1330 4580
rect -1250 4640 -1210 4680
rect -1250 4540 -1210 4580
rect -1130 4640 -1090 4680
rect -1130 4540 -1090 4580
rect -1010 4640 -970 4680
rect -1010 4540 -970 4580
rect -890 4640 -850 4680
rect -890 4540 -850 4580
rect -770 4640 -730 4680
rect -770 4540 -730 4580
rect -650 4640 -610 4680
rect -650 4540 -610 4580
rect -530 4640 -490 4680
rect -530 4540 -490 4580
rect -410 4640 -370 4680
rect -410 4540 -370 4580
rect -290 4640 -250 4680
rect -290 4540 -250 4580
rect -170 4640 -130 4680
rect -170 4540 -130 4580
rect -50 4640 -10 4680
rect -50 4540 -10 4580
rect 590 4640 630 4680
rect 590 4540 630 4580
rect 710 4640 750 4680
rect 710 4540 750 4580
rect 830 4640 870 4680
rect 830 4540 870 4580
rect 950 4640 990 4680
rect 950 4540 990 4580
rect 1070 4640 1110 4680
rect 1070 4540 1110 4580
rect 1190 4640 1230 4680
rect 1190 4540 1230 4580
rect 1310 4640 1350 4680
rect 1310 4540 1350 4580
rect 1430 4640 1470 4680
rect 1430 4540 1470 4580
rect 1550 4640 1590 4680
rect 1550 4540 1590 4580
rect 1670 4640 1710 4680
rect 1670 4540 1710 4580
rect 1790 4640 1830 4680
rect 1790 4540 1830 4580
rect 1910 4640 1950 4680
rect 1910 4540 1950 4580
rect 2030 4640 2070 4680
rect 2030 4540 2070 4580
rect 2150 4640 2190 4680
rect 2150 4540 2190 4580
rect 2270 4640 2310 4680
rect 2270 4540 2310 4580
rect 2390 4640 2430 4680
rect 2390 4540 2430 4580
rect 2510 4640 2550 4680
rect 2510 4540 2550 4580
rect 2630 4640 2670 4680
rect 2630 4540 2670 4580
rect 2750 4640 2790 4680
rect 2750 4540 2790 4580
rect 2870 4640 2910 4680
rect 2870 4540 2910 4580
rect 2990 4640 3030 4680
rect 5580 4620 5620 4660
rect 5710 4720 5750 4760
rect 5710 4620 5750 4660
rect 5840 4720 5880 4760
rect 5840 4620 5880 4660
rect 5970 4720 6010 4760
rect 5970 4620 6010 4660
rect 6100 4720 6140 4760
rect 6100 4620 6140 4660
rect 6230 4720 6270 4760
rect 6230 4620 6270 4660
rect 6360 4720 6400 4760
rect 6360 4620 6400 4660
rect 6720 4720 6760 4760
rect 6720 4620 6760 4660
rect 6850 4720 6890 4760
rect 6850 4620 6890 4660
rect 6980 4720 7020 4760
rect 6980 4620 7020 4660
rect 7110 4720 7150 4760
rect 7110 4620 7150 4660
rect 7240 4720 7280 4760
rect 7240 4620 7280 4660
rect 7370 4720 7410 4760
rect 7370 4620 7410 4660
rect 7500 4720 7540 4760
rect 7500 4620 7540 4660
rect 9570 4750 9640 4820
rect 2990 4540 3030 4580
rect -2270 4410 -2230 4450
rect -2090 4420 -2050 4460
rect -1610 4420 -1570 4460
rect -1370 4420 -1330 4460
rect -890 4420 -850 4460
rect -650 4420 -610 4460
rect -230 4420 -190 4460
rect 770 4420 810 4460
rect 1190 4420 1230 4460
rect 1430 4420 1470 4460
rect 1910 4420 1950 4460
rect 2150 4420 2190 4460
rect 2630 4420 2670 4460
rect 2810 4410 2850 4450
rect 6050 4460 6090 4500
rect 7130 4350 7170 4390
rect 8250 4350 8290 4390
rect 5650 4190 5690 4230
rect 7650 4190 7690 4230
rect 5650 4070 5690 4110
rect 5650 3970 5690 4010
rect 5650 3870 5690 3910
rect -1446 3818 -1412 3852
rect -1288 3818 -1254 3852
rect -964 3818 -930 3852
rect -810 3818 -776 3852
rect -486 3818 -452 3852
rect -170 3770 -130 3810
rect -1610 3700 -1570 3740
rect -1490 3700 -1450 3740
rect -1370 3700 -1330 3740
rect -1250 3700 -1210 3740
rect -1130 3700 -1090 3740
rect -1010 3700 -970 3740
rect -890 3700 -850 3740
rect -770 3700 -730 3740
rect -650 3700 -610 3740
rect -530 3700 -490 3740
rect -410 3700 -370 3740
rect -170 3690 -130 3730
rect -1547 3588 -1513 3622
rect -1187 3588 -1153 3622
rect -1067 3588 -1033 3622
rect -707 3588 -673 3622
rect -587 3588 -553 3622
rect -170 3610 -130 3650
rect 710 3770 750 3810
rect 1032 3818 1066 3852
rect 1356 3818 1390 3852
rect 1510 3818 1544 3852
rect 1834 3818 1868 3852
rect 1992 3818 2026 3852
rect 5650 3770 5690 3810
rect 710 3690 750 3730
rect 950 3700 990 3740
rect 1070 3700 1110 3740
rect 1190 3700 1230 3740
rect 1310 3700 1350 3740
rect 1430 3700 1470 3740
rect 1550 3700 1590 3740
rect 1670 3700 1710 3740
rect 1790 3700 1830 3740
rect 1910 3700 1950 3740
rect 2030 3700 2070 3740
rect 2150 3700 2190 3740
rect 5650 3670 5690 3710
rect 5850 4070 5890 4110
rect 5850 3970 5890 4010
rect 5850 3870 5890 3910
rect 5850 3770 5890 3810
rect 5850 3670 5890 3710
rect 6050 4070 6090 4110
rect 6050 3970 6090 4010
rect 6050 3870 6090 3910
rect 6050 3770 6090 3810
rect 6050 3670 6090 3710
rect 6250 4070 6290 4110
rect 6250 3970 6290 4010
rect 6250 3870 6290 3910
rect 6250 3770 6290 3810
rect 6250 3670 6290 3710
rect 6450 4070 6490 4110
rect 6450 3970 6490 4010
rect 6450 3870 6490 3910
rect 6450 3770 6490 3810
rect 6450 3670 6490 3710
rect 6650 4070 6690 4110
rect 6650 3970 6690 4010
rect 6650 3870 6690 3910
rect 6650 3770 6690 3810
rect 6650 3670 6690 3710
rect 6850 4070 6890 4110
rect 6850 3970 6890 4010
rect 6850 3870 6890 3910
rect 6850 3770 6890 3810
rect 6850 3670 6890 3710
rect 7050 4070 7090 4110
rect 7050 3970 7090 4010
rect 7050 3870 7090 3910
rect 7050 3770 7090 3810
rect 7050 3670 7090 3710
rect 7250 4070 7290 4110
rect 7250 3970 7290 4010
rect 7250 3870 7290 3910
rect 7250 3770 7290 3810
rect 7250 3670 7290 3710
rect 7450 4070 7490 4110
rect 7450 3970 7490 4010
rect 7450 3870 7490 3910
rect 7450 3770 7490 3810
rect 7450 3670 7490 3710
rect 7650 4070 7690 4110
rect 7650 3970 7690 4010
rect 7650 3870 7690 3910
rect 7650 3770 7690 3810
rect 7650 3670 7690 3710
rect 710 3610 750 3650
rect 1133 3588 1167 3622
rect 1253 3588 1287 3622
rect 1613 3588 1647 3622
rect 1733 3588 1767 3622
rect 2093 3588 2127 3622
rect 6450 3550 6490 3590
rect 6850 3550 6890 3590
rect -2230 3170 -2190 3210
rect -2050 3210 -2010 3250
rect -1810 3210 -1770 3250
rect -1570 3210 -1530 3250
rect -1330 3210 -1290 3250
rect -690 3210 -650 3250
rect -450 3210 -410 3250
rect -210 3210 -170 3250
rect 90 3180 130 3220
rect 450 3180 490 3220
rect 750 3210 790 3250
rect 990 3210 1030 3250
rect 1230 3210 1270 3250
rect 1870 3210 1910 3250
rect 2110 3210 2150 3250
rect 2350 3210 2390 3250
rect 2590 3210 2630 3250
rect 9140 3160 9180 3200
rect 2770 3090 2810 3130
rect 2770 2990 2810 3030
rect 2770 2890 2810 2930
rect 2770 2790 2810 2830
rect 9340 2820 9400 2880
rect 2770 2690 2810 2730
rect -1070 2570 -1030 2610
rect 1610 2570 1650 2610
rect -1810 2300 -1770 2340
rect -1650 2300 -1610 2340
rect -1490 2300 -1450 2340
rect -1330 2300 -1290 2340
rect -1170 2300 -1130 2340
rect -1010 2300 -970 2340
rect -850 2300 -810 2340
rect -690 2300 -650 2340
rect -530 2300 -490 2340
rect -370 2300 -330 2340
rect -210 2300 -170 2340
rect -50 2300 -10 2340
rect 110 2300 150 2340
rect 270 2300 310 2340
rect 430 2300 470 2340
rect 590 2300 630 2340
rect 750 2300 790 2340
rect 910 2300 950 2340
rect 1070 2300 1110 2340
rect 1230 2300 1270 2340
rect 1390 2300 1430 2340
rect 1550 2300 1590 2340
rect 1710 2300 1750 2340
rect 1870 2300 1910 2340
rect 2030 2300 2070 2340
rect 2190 2300 2230 2340
rect -1890 2130 -1850 2170
rect 2500 2170 2540 2210
rect 2500 2090 2540 2130
rect -428 1730 -378 1780
rect 970 1730 1020 1780
rect -1330 1164 -1324 1170
rect -1324 1164 -1296 1170
rect -1330 1136 -1296 1164
rect -1230 1136 -1196 1170
rect -1130 1136 -1096 1170
rect -1030 1164 -998 1170
rect -998 1164 -996 1170
rect -930 1164 -908 1170
rect -908 1164 -896 1170
rect -830 1164 -818 1170
rect -818 1164 -796 1170
rect -1030 1136 -996 1164
rect -930 1136 -896 1164
rect -830 1136 -796 1164
rect -1330 1036 -1296 1070
rect -1230 1036 -1196 1070
rect -1130 1036 -1096 1070
rect -1030 1036 -996 1070
rect -930 1036 -896 1070
rect -830 1036 -796 1070
rect -1330 936 -1296 970
rect -1230 936 -1196 970
rect -1130 936 -1096 970
rect -1030 936 -996 970
rect -930 936 -896 970
rect -830 936 -796 970
rect -1330 838 -1296 870
rect -1330 836 -1324 838
rect -1324 836 -1296 838
rect -1230 836 -1196 870
rect -1130 836 -1096 870
rect -1030 838 -996 870
rect -930 838 -896 870
rect -830 838 -796 870
rect -1030 836 -998 838
rect -998 836 -996 838
rect -930 836 -908 838
rect -908 836 -896 838
rect -830 836 -818 838
rect -818 836 -796 838
rect -1330 748 -1296 770
rect -1330 736 -1324 748
rect -1324 736 -1296 748
rect -1230 736 -1196 770
rect -1130 736 -1096 770
rect -1030 748 -996 770
rect -930 748 -896 770
rect -830 748 -796 770
rect -1030 736 -998 748
rect -998 736 -996 748
rect -930 736 -908 748
rect -908 736 -896 748
rect -830 736 -818 748
rect -818 736 -796 748
rect -1330 658 -1296 670
rect -1330 636 -1324 658
rect -1324 636 -1296 658
rect -1230 636 -1196 670
rect -1130 636 -1096 670
rect -1030 658 -996 670
rect -930 658 -896 670
rect -830 658 -796 670
rect -1030 636 -998 658
rect -998 636 -996 658
rect -930 636 -908 658
rect -908 636 -896 658
rect -830 636 -818 658
rect -818 636 -796 658
rect 30 1164 36 1170
rect 36 1164 64 1170
rect 30 1136 64 1164
rect 130 1136 164 1170
rect 230 1136 264 1170
rect 330 1164 362 1170
rect 362 1164 364 1170
rect 430 1164 452 1170
rect 452 1164 464 1170
rect 530 1164 542 1170
rect 542 1164 564 1170
rect 330 1136 364 1164
rect 430 1136 464 1164
rect 530 1136 564 1164
rect 30 1036 64 1070
rect 130 1036 164 1070
rect 230 1036 264 1070
rect 330 1036 364 1070
rect 430 1036 464 1070
rect 530 1036 564 1070
rect 30 936 64 970
rect 130 936 164 970
rect 230 936 264 970
rect 330 936 364 970
rect 430 936 464 970
rect 530 936 564 970
rect 30 838 64 870
rect 30 836 36 838
rect 36 836 64 838
rect 130 836 164 870
rect 230 836 264 870
rect 330 838 364 870
rect 430 838 464 870
rect 530 838 564 870
rect 330 836 362 838
rect 362 836 364 838
rect 430 836 452 838
rect 452 836 464 838
rect 530 836 542 838
rect 542 836 564 838
rect 30 748 64 770
rect 30 736 36 748
rect 36 736 64 748
rect 130 736 164 770
rect 230 736 264 770
rect 330 748 364 770
rect 430 748 464 770
rect 530 748 564 770
rect 330 736 362 748
rect 362 736 364 748
rect 430 736 452 748
rect 452 736 464 748
rect 530 736 542 748
rect 542 736 564 748
rect 30 658 64 670
rect 30 636 36 658
rect 36 636 64 658
rect 130 636 164 670
rect 230 636 264 670
rect 330 658 364 670
rect 430 658 464 670
rect 530 658 564 670
rect 330 636 362 658
rect 362 636 364 658
rect 430 636 452 658
rect 452 636 464 658
rect 530 636 542 658
rect 542 636 564 658
rect 1390 1164 1396 1170
rect 1396 1164 1424 1170
rect 1390 1136 1424 1164
rect 1490 1136 1524 1170
rect 1590 1136 1624 1170
rect 1690 1164 1722 1170
rect 1722 1164 1724 1170
rect 1790 1164 1812 1170
rect 1812 1164 1824 1170
rect 1890 1164 1902 1170
rect 1902 1164 1924 1170
rect 1690 1136 1724 1164
rect 1790 1136 1824 1164
rect 1890 1136 1924 1164
rect 1390 1036 1424 1070
rect 1490 1036 1524 1070
rect 1590 1036 1624 1070
rect 1690 1036 1724 1070
rect 1790 1036 1824 1070
rect 1890 1036 1924 1070
rect 1390 936 1424 970
rect 1490 936 1524 970
rect 1590 936 1624 970
rect 1690 936 1724 970
rect 1790 936 1824 970
rect 1890 936 1924 970
rect 1390 838 1424 870
rect 1390 836 1396 838
rect 1396 836 1424 838
rect 1490 836 1524 870
rect 1590 836 1624 870
rect 1690 838 1724 870
rect 1790 838 1824 870
rect 1890 838 1924 870
rect 1690 836 1722 838
rect 1722 836 1724 838
rect 1790 836 1812 838
rect 1812 836 1824 838
rect 1890 836 1902 838
rect 1902 836 1924 838
rect 1390 748 1424 770
rect 1390 736 1396 748
rect 1396 736 1424 748
rect 1490 736 1524 770
rect 1590 736 1624 770
rect 1690 748 1724 770
rect 1790 748 1824 770
rect 1890 748 1924 770
rect 1690 736 1722 748
rect 1722 736 1724 748
rect 1790 736 1812 748
rect 1812 736 1824 748
rect 1890 736 1902 748
rect 1902 736 1924 748
rect 1390 658 1424 670
rect 1390 636 1396 658
rect 1396 636 1424 658
rect 1490 636 1524 670
rect 1590 636 1624 670
rect 1690 658 1724 670
rect 1790 658 1824 670
rect 1890 658 1924 670
rect 1690 636 1722 658
rect 1722 636 1724 658
rect 1790 636 1812 658
rect 1812 636 1824 658
rect 1890 636 1902 658
rect 1902 636 1924 658
rect -2300 -70 -2250 -20
rect -2850 -500 -2800 -450
rect -2730 -450 -2680 -400
rect -1330 -196 -1324 -190
rect -1324 -196 -1296 -190
rect -1330 -224 -1296 -196
rect -1230 -224 -1196 -190
rect -1130 -224 -1096 -190
rect -1030 -196 -998 -190
rect -998 -196 -996 -190
rect -930 -196 -908 -190
rect -908 -196 -896 -190
rect -830 -196 -818 -190
rect -818 -196 -796 -190
rect -1030 -224 -996 -196
rect -930 -224 -896 -196
rect -830 -224 -796 -196
rect -1330 -324 -1296 -290
rect -1230 -324 -1196 -290
rect -1130 -324 -1096 -290
rect -1030 -324 -996 -290
rect -930 -324 -896 -290
rect -830 -324 -796 -290
rect -1330 -424 -1296 -390
rect -1230 -424 -1196 -390
rect -1130 -424 -1096 -390
rect -1030 -424 -996 -390
rect -930 -424 -896 -390
rect -830 -424 -796 -390
rect -1330 -522 -1296 -490
rect -1330 -524 -1324 -522
rect -1324 -524 -1296 -522
rect -1230 -524 -1196 -490
rect -1130 -524 -1096 -490
rect -1030 -522 -996 -490
rect -930 -522 -896 -490
rect -830 -522 -796 -490
rect -1030 -524 -998 -522
rect -998 -524 -996 -522
rect -930 -524 -908 -522
rect -908 -524 -896 -522
rect -830 -524 -818 -522
rect -818 -524 -796 -522
rect -1330 -612 -1296 -590
rect -1330 -624 -1324 -612
rect -1324 -624 -1296 -612
rect -1230 -624 -1196 -590
rect -1130 -624 -1096 -590
rect -1030 -612 -996 -590
rect -930 -612 -896 -590
rect -830 -612 -796 -590
rect -1030 -624 -998 -612
rect -998 -624 -996 -612
rect -930 -624 -908 -612
rect -908 -624 -896 -612
rect -830 -624 -818 -612
rect -818 -624 -796 -612
rect -1330 -702 -1296 -690
rect -1330 -724 -1324 -702
rect -1324 -724 -1296 -702
rect -1230 -724 -1196 -690
rect -1130 -724 -1096 -690
rect -1030 -702 -996 -690
rect -930 -702 -896 -690
rect -830 -702 -796 -690
rect -1030 -724 -998 -702
rect -998 -724 -996 -702
rect -930 -724 -908 -702
rect -908 -724 -896 -702
rect -830 -724 -818 -702
rect -818 -724 -796 -702
rect 30 -196 36 -190
rect 36 -196 64 -190
rect 30 -224 64 -196
rect 130 -224 164 -190
rect 230 -224 264 -190
rect 330 -196 362 -190
rect 362 -196 364 -190
rect 430 -196 452 -190
rect 452 -196 464 -190
rect 530 -196 542 -190
rect 542 -196 564 -190
rect 330 -224 364 -196
rect 430 -224 464 -196
rect 530 -224 564 -196
rect 30 -324 64 -290
rect 130 -324 164 -290
rect 230 -324 264 -290
rect 330 -324 364 -290
rect 430 -324 464 -290
rect 530 -324 564 -290
rect 30 -424 64 -390
rect 130 -424 164 -390
rect 230 -424 264 -390
rect 330 -424 364 -390
rect 430 -424 464 -390
rect 530 -424 564 -390
rect 30 -522 64 -490
rect 30 -524 36 -522
rect 36 -524 64 -522
rect 130 -524 164 -490
rect 230 -524 264 -490
rect 330 -522 364 -490
rect 430 -522 464 -490
rect 530 -522 564 -490
rect 330 -524 362 -522
rect 362 -524 364 -522
rect 430 -524 452 -522
rect 452 -524 464 -522
rect 530 -524 542 -522
rect 542 -524 564 -522
rect 30 -612 64 -590
rect 30 -624 36 -612
rect 36 -624 64 -612
rect 130 -624 164 -590
rect 230 -624 264 -590
rect 330 -612 364 -590
rect 430 -612 464 -590
rect 530 -612 564 -590
rect 330 -624 362 -612
rect 362 -624 364 -612
rect 430 -624 452 -612
rect 452 -624 464 -612
rect 530 -624 542 -612
rect 542 -624 564 -612
rect 30 -702 64 -690
rect 30 -724 36 -702
rect 36 -724 64 -702
rect 130 -724 164 -690
rect 230 -724 264 -690
rect 330 -702 364 -690
rect 430 -702 464 -690
rect 530 -702 564 -690
rect 330 -724 362 -702
rect 362 -724 364 -702
rect 430 -724 452 -702
rect 452 -724 464 -702
rect 530 -724 542 -702
rect 542 -724 564 -702
rect 1390 -196 1396 -190
rect 1396 -196 1424 -190
rect 1390 -224 1424 -196
rect 1490 -224 1524 -190
rect 1590 -224 1624 -190
rect 1690 -196 1722 -190
rect 1722 -196 1724 -190
rect 1790 -196 1812 -190
rect 1812 -196 1824 -190
rect 1890 -196 1902 -190
rect 1902 -196 1924 -190
rect 1690 -224 1724 -196
rect 1790 -224 1824 -196
rect 1890 -224 1924 -196
rect 1390 -324 1424 -290
rect 1490 -324 1524 -290
rect 1590 -324 1624 -290
rect 1690 -324 1724 -290
rect 1790 -324 1824 -290
rect 1890 -324 1924 -290
rect 1390 -424 1424 -390
rect 1490 -424 1524 -390
rect 1590 -424 1624 -390
rect 1690 -424 1724 -390
rect 1790 -424 1824 -390
rect 1890 -424 1924 -390
rect 1390 -522 1424 -490
rect 1390 -524 1396 -522
rect 1396 -524 1424 -522
rect 1490 -524 1524 -490
rect 1590 -524 1624 -490
rect 1690 -522 1724 -490
rect 1790 -522 1824 -490
rect 1890 -522 1924 -490
rect 1690 -524 1722 -522
rect 1722 -524 1724 -522
rect 1790 -524 1812 -522
rect 1812 -524 1824 -522
rect 1890 -524 1902 -522
rect 1902 -524 1924 -522
rect 1390 -612 1424 -590
rect 1390 -624 1396 -612
rect 1396 -624 1424 -612
rect 1490 -624 1524 -590
rect 1590 -624 1624 -590
rect 1690 -612 1724 -590
rect 1790 -612 1824 -590
rect 1890 -612 1924 -590
rect 1690 -624 1722 -612
rect 1722 -624 1724 -612
rect 1790 -624 1812 -612
rect 1812 -624 1824 -612
rect 1890 -624 1902 -612
rect 1902 -624 1924 -612
rect 1390 -702 1424 -690
rect 1390 -724 1396 -702
rect 1396 -724 1424 -702
rect 1490 -724 1524 -690
rect 1590 -724 1624 -690
rect 1690 -702 1724 -690
rect 1790 -702 1824 -690
rect 1890 -702 1924 -690
rect 1690 -724 1722 -702
rect 1722 -724 1724 -702
rect 1790 -724 1812 -702
rect 1812 -724 1824 -702
rect 1890 -724 1902 -702
rect 1902 -724 1924 -702
rect 2710 -70 2760 -20
rect 3490 -712 3540 -662
rect 2830 -920 2880 -870
rect -3020 -1430 -2980 -1390
rect -2850 -1848 -2800 -1798
rect -2490 -2058 -2440 -2008
rect -2060 -2208 -2010 -2158
rect -1330 -1556 -1324 -1550
rect -1324 -1556 -1296 -1550
rect -1330 -1584 -1296 -1556
rect -1230 -1584 -1196 -1550
rect -1130 -1584 -1096 -1550
rect -1030 -1556 -998 -1550
rect -998 -1556 -996 -1550
rect -930 -1556 -908 -1550
rect -908 -1556 -896 -1550
rect -830 -1556 -818 -1550
rect -818 -1556 -796 -1550
rect -1030 -1584 -996 -1556
rect -930 -1584 -896 -1556
rect -830 -1584 -796 -1556
rect -1330 -1684 -1296 -1650
rect -1230 -1684 -1196 -1650
rect -1130 -1684 -1096 -1650
rect -1030 -1684 -996 -1650
rect -930 -1684 -896 -1650
rect -830 -1684 -796 -1650
rect -1330 -1784 -1296 -1750
rect -1230 -1784 -1196 -1750
rect -1130 -1784 -1096 -1750
rect -1030 -1784 -996 -1750
rect -930 -1784 -896 -1750
rect -830 -1784 -796 -1750
rect -1330 -1882 -1296 -1850
rect -1330 -1884 -1324 -1882
rect -1324 -1884 -1296 -1882
rect -1230 -1884 -1196 -1850
rect -1130 -1884 -1096 -1850
rect -1030 -1882 -996 -1850
rect -930 -1882 -896 -1850
rect -830 -1882 -796 -1850
rect -1030 -1884 -998 -1882
rect -998 -1884 -996 -1882
rect -930 -1884 -908 -1882
rect -908 -1884 -896 -1882
rect -830 -1884 -818 -1882
rect -818 -1884 -796 -1882
rect -1330 -1972 -1296 -1950
rect -1330 -1984 -1324 -1972
rect -1324 -1984 -1296 -1972
rect -1230 -1984 -1196 -1950
rect -1130 -1984 -1096 -1950
rect -1030 -1972 -996 -1950
rect -930 -1972 -896 -1950
rect -830 -1972 -796 -1950
rect -1030 -1984 -998 -1972
rect -998 -1984 -996 -1972
rect -930 -1984 -908 -1972
rect -908 -1984 -896 -1972
rect -830 -1984 -818 -1972
rect -818 -1984 -796 -1972
rect -1330 -2062 -1296 -2050
rect -1330 -2084 -1324 -2062
rect -1324 -2084 -1296 -2062
rect -1230 -2084 -1196 -2050
rect -1130 -2084 -1096 -2050
rect -1030 -2062 -996 -2050
rect -930 -2062 -896 -2050
rect -830 -2062 -796 -2050
rect -1030 -2084 -998 -2062
rect -998 -2084 -996 -2062
rect -930 -2084 -908 -2062
rect -908 -2084 -896 -2062
rect -830 -2084 -818 -2062
rect -818 -2084 -796 -2062
rect 30 -1556 36 -1550
rect 36 -1556 64 -1550
rect 30 -1584 64 -1556
rect 130 -1584 164 -1550
rect 230 -1584 264 -1550
rect 330 -1556 362 -1550
rect 362 -1556 364 -1550
rect 430 -1556 452 -1550
rect 452 -1556 464 -1550
rect 530 -1556 542 -1550
rect 542 -1556 564 -1550
rect 330 -1584 364 -1556
rect 430 -1584 464 -1556
rect 530 -1584 564 -1556
rect 30 -1684 64 -1650
rect 130 -1684 164 -1650
rect 230 -1684 264 -1650
rect 330 -1684 364 -1650
rect 430 -1684 464 -1650
rect 530 -1684 564 -1650
rect 30 -1784 64 -1750
rect 130 -1784 164 -1750
rect 230 -1784 264 -1750
rect 330 -1784 364 -1750
rect 430 -1784 464 -1750
rect 530 -1784 564 -1750
rect 30 -1882 64 -1850
rect 30 -1884 36 -1882
rect 36 -1884 64 -1882
rect 130 -1884 164 -1850
rect 230 -1884 264 -1850
rect 330 -1882 364 -1850
rect 430 -1882 464 -1850
rect 530 -1882 564 -1850
rect 330 -1884 362 -1882
rect 362 -1884 364 -1882
rect 430 -1884 452 -1882
rect 452 -1884 464 -1882
rect 530 -1884 542 -1882
rect 542 -1884 564 -1882
rect 30 -1972 64 -1950
rect 30 -1984 36 -1972
rect 36 -1984 64 -1972
rect 130 -1984 164 -1950
rect 230 -1984 264 -1950
rect 330 -1972 364 -1950
rect 430 -1972 464 -1950
rect 530 -1972 564 -1950
rect 330 -1984 362 -1972
rect 362 -1984 364 -1972
rect 430 -1984 452 -1972
rect 452 -1984 464 -1972
rect 530 -1984 542 -1972
rect 542 -1984 564 -1972
rect 30 -2062 64 -2050
rect 30 -2084 36 -2062
rect 36 -2084 64 -2062
rect 130 -2084 164 -2050
rect 230 -2084 264 -2050
rect 330 -2062 364 -2050
rect 430 -2062 464 -2050
rect 530 -2062 564 -2050
rect 330 -2084 362 -2062
rect 362 -2084 364 -2062
rect 430 -2084 452 -2062
rect 452 -2084 464 -2062
rect 530 -2084 542 -2062
rect 542 -2084 564 -2062
rect 1390 -1556 1396 -1550
rect 1396 -1556 1424 -1550
rect 1390 -1584 1424 -1556
rect 1490 -1584 1524 -1550
rect 1590 -1584 1624 -1550
rect 1690 -1556 1722 -1550
rect 1722 -1556 1724 -1550
rect 1790 -1556 1812 -1550
rect 1812 -1556 1824 -1550
rect 1890 -1556 1902 -1550
rect 1902 -1556 1924 -1550
rect 1690 -1584 1724 -1556
rect 1790 -1584 1824 -1556
rect 1890 -1584 1924 -1556
rect 1390 -1684 1424 -1650
rect 1490 -1684 1524 -1650
rect 1590 -1684 1624 -1650
rect 1690 -1684 1724 -1650
rect 1790 -1684 1824 -1650
rect 1890 -1684 1924 -1650
rect 1390 -1784 1424 -1750
rect 1490 -1784 1524 -1750
rect 1590 -1784 1624 -1750
rect 1690 -1784 1724 -1750
rect 1790 -1784 1824 -1750
rect 1890 -1784 1924 -1750
rect 1390 -1882 1424 -1850
rect 1390 -1884 1396 -1882
rect 1396 -1884 1424 -1882
rect 1490 -1884 1524 -1850
rect 1590 -1884 1624 -1850
rect 1690 -1882 1724 -1850
rect 1790 -1882 1824 -1850
rect 1890 -1882 1924 -1850
rect 1690 -1884 1722 -1882
rect 1722 -1884 1724 -1882
rect 1790 -1884 1812 -1882
rect 1812 -1884 1824 -1882
rect 1890 -1884 1902 -1882
rect 1902 -1884 1924 -1882
rect 1390 -1972 1424 -1950
rect 1390 -1984 1396 -1972
rect 1396 -1984 1424 -1972
rect 1490 -1984 1524 -1950
rect 1590 -1984 1624 -1950
rect 1690 -1972 1724 -1950
rect 1790 -1972 1824 -1950
rect 1890 -1972 1924 -1950
rect 1690 -1984 1722 -1972
rect 1722 -1984 1724 -1972
rect 1790 -1984 1812 -1972
rect 1812 -1984 1824 -1972
rect 1890 -1984 1902 -1972
rect 1902 -1984 1924 -1972
rect 1390 -2062 1424 -2050
rect 1390 -2084 1396 -2062
rect 1396 -2084 1424 -2062
rect 1490 -2084 1524 -2050
rect 1590 -2084 1624 -2050
rect 1690 -2062 1724 -2050
rect 1790 -2062 1824 -2050
rect 1890 -2062 1924 -2050
rect 1690 -2084 1722 -2062
rect 1722 -2084 1724 -2062
rect 1790 -2084 1812 -2062
rect 1812 -2084 1824 -2062
rect 1890 -2084 1902 -2062
rect 1902 -2084 1924 -2062
rect 3010 -1490 3050 -1450
rect 2830 -2058 2880 -2008
rect 3490 -2058 3540 -2008
rect 2470 -2208 2520 -2158
rect 270 -2580 310 -2540
rect 270 -2660 310 -2620
rect 270 -2740 310 -2700
rect 2910 -2960 2950 -2920
rect 5360 -2960 5400 -2920
<< metal1 >>
rect 9410 14270 9490 14280
rect 9410 14210 9420 14270
rect 9480 14210 9490 14270
rect 8920 14160 9160 14170
rect 8920 14100 8930 14160
rect 8990 14100 9010 14160
rect 9070 14100 9090 14160
rect 9150 14100 9160 14160
rect 8920 14080 9160 14100
rect 8920 14020 8930 14080
rect 8990 14020 9010 14080
rect 9070 14020 9090 14080
rect 9150 14020 9160 14080
rect 8920 14000 9160 14020
rect 8920 13940 8930 14000
rect 8990 13940 9010 14000
rect 9070 13940 9090 14000
rect 9150 13940 9160 14000
rect -1350 13050 -1270 13060
rect -1350 12990 -1340 13050
rect -1280 12990 -1270 13050
rect -1350 12980 -1270 12990
rect -1130 13050 -1050 13060
rect -1130 12990 -1120 13050
rect -1060 12990 -1050 13050
rect -1130 12980 -1050 12990
rect -660 13050 -580 13060
rect -660 12990 -650 13050
rect -590 12990 -580 13050
rect -660 12980 -580 12990
rect -320 13050 -240 13060
rect -320 12990 -310 13050
rect -250 12990 -240 13050
rect -320 12980 -240 12990
rect -100 13050 -20 13060
rect -100 12990 -90 13050
rect -30 12990 -20 13050
rect -100 12980 -20 12990
rect 340 13050 420 13060
rect 340 12990 350 13050
rect 410 12990 420 13050
rect 340 12980 420 12990
rect 1020 13050 1100 13060
rect 1020 12990 1030 13050
rect 1090 12990 1100 13050
rect 1020 12980 1100 12990
rect 1240 13050 1320 13060
rect 1240 12990 1250 13050
rect 1310 12990 1320 13050
rect 1240 12980 1320 12990
rect 1710 13050 1790 13060
rect 1710 12990 1720 13050
rect 1780 12990 1790 13050
rect 1710 12980 1790 12990
rect 2170 13050 2250 13060
rect 2170 12990 2180 13050
rect 2240 12990 2250 13050
rect 2170 12980 2250 12990
rect 2520 13050 2600 13060
rect 2520 12990 2530 13050
rect 2590 12990 2600 13050
rect 2520 12980 2600 12990
rect 2770 13050 2850 13060
rect 2770 12990 2780 13050
rect 2840 12990 2850 13050
rect 2770 12980 2850 12990
rect 2990 13050 3070 13060
rect 2990 12990 3000 13050
rect 3060 12990 3070 13050
rect 2990 12980 3070 12990
rect 3320 13050 3400 13060
rect 3320 12990 3330 13050
rect 3390 12990 3400 13050
rect 3320 12980 3400 12990
rect 3980 13050 4060 13060
rect 3980 12990 3990 13050
rect 4050 12990 4060 13050
rect 3980 12980 4060 12990
rect 4200 13050 4280 13060
rect 4200 12990 4210 13050
rect 4270 12990 4280 13050
rect 4200 12980 4280 12990
rect 4770 13050 4850 13060
rect 4770 12990 4780 13050
rect 4840 12990 4850 13050
rect 4770 12980 4850 12990
rect 5030 13050 5110 13060
rect 5030 12990 5040 13050
rect 5100 12990 5110 13050
rect 5030 12980 5110 12990
rect 5280 13050 5360 13060
rect 5280 12990 5290 13050
rect 5350 12990 5360 13050
rect 5280 12980 5360 12990
rect 5500 13050 5580 13060
rect 5500 12990 5510 13050
rect 5570 12990 5580 13050
rect 5500 12980 5580 12990
rect 6050 13050 6130 13060
rect 6050 12990 6060 13050
rect 6120 12990 6130 13050
rect 6050 12980 6130 12990
rect 6330 13050 6410 13060
rect 6330 12990 6340 13050
rect 6400 12990 6410 13050
rect 6330 12980 6410 12990
rect 6580 13050 6660 13060
rect 6580 12990 6590 13050
rect 6650 12990 6660 13050
rect 6580 12980 6660 12990
rect 6800 13050 6880 13060
rect 6800 12990 6810 13050
rect 6870 12990 6880 13050
rect 6800 12980 6880 12990
rect 7350 13050 7430 13060
rect 7350 12990 7360 13050
rect 7420 12990 7430 13050
rect 7350 12980 7430 12990
rect 7630 13050 7710 13060
rect 7630 12990 7640 13050
rect 7700 12990 7710 13050
rect 7630 12980 7710 12990
rect 7880 13050 7960 13060
rect 7880 12990 7890 13050
rect 7950 12990 7960 13050
rect 7880 12980 7960 12990
rect 8100 13050 8180 13060
rect 8100 12990 8110 13050
rect 8170 12990 8180 13050
rect 8100 12980 8180 12990
rect 8650 13050 8730 13060
rect 8650 12990 8660 13050
rect 8720 12990 8730 13050
rect 8650 12980 8730 12990
rect -1510 12930 -1430 12950
rect -1510 12890 -1490 12930
rect -1450 12910 -480 12930
rect -1450 12890 -540 12910
rect -1510 12870 -1430 12890
rect -560 12870 -540 12890
rect -500 12870 -480 12910
rect -430 12920 2150 12940
rect -430 12880 -410 12920
rect -370 12900 530 12920
rect -370 12880 -350 12900
rect -430 12870 -350 12880
rect 510 12880 530 12900
rect 570 12900 2090 12920
rect 570 12880 590 12900
rect 510 12870 590 12880
rect 2070 12880 2090 12900
rect 2130 12880 2150 12920
rect 4684 12930 4750 12950
rect 4684 12910 4694 12930
rect 2070 12870 2150 12880
rect 2340 12890 4694 12910
rect 4734 12890 4750 12930
rect 2340 12870 4750 12890
rect -560 12850 -480 12870
rect 100 12690 180 12710
rect -1780 12670 -1700 12680
rect -1780 12610 -1770 12670
rect -1710 12610 -1700 12670
rect -1780 8580 -1700 12610
rect -1570 12670 -1490 12680
rect -1570 12610 -1560 12670
rect -1500 12610 -1490 12670
rect 100 12650 120 12690
rect 160 12680 180 12690
rect 620 12690 700 12710
rect 620 12680 640 12690
rect 160 12650 640 12680
rect 680 12650 700 12690
rect 100 12640 700 12650
rect 2340 12700 2380 12870
rect 8920 12760 9160 13940
rect 9410 13890 9490 14210
rect 9410 13850 9430 13890
rect 9470 13850 9490 13890
rect 9410 13830 9490 13850
rect 9930 14270 10010 14280
rect 9930 14210 9940 14270
rect 10000 14210 10010 14270
rect 9930 13890 10010 14210
rect 9930 13850 9950 13890
rect 9990 13850 10010 13890
rect 9930 13830 10010 13850
rect 10450 14270 10530 14280
rect 10450 14210 10460 14270
rect 10520 14210 10530 14270
rect 10450 13890 10530 14210
rect 10450 13850 10470 13890
rect 10510 13850 10530 13890
rect 10450 13830 10530 13850
rect 10940 14270 11020 14280
rect 10940 14210 10950 14270
rect 11010 14210 11020 14270
rect 10940 13890 11020 14210
rect 10940 13850 10960 13890
rect 11000 13850 11020 13890
rect 10940 13830 11020 13850
rect 11270 14160 11510 14170
rect 11270 14100 11280 14160
rect 11340 14100 11360 14160
rect 11420 14100 11440 14160
rect 11500 14100 11510 14160
rect 11270 14080 11510 14100
rect 11270 14020 11280 14080
rect 11340 14020 11360 14080
rect 11420 14020 11440 14080
rect 11500 14020 11510 14080
rect 11270 14000 11510 14020
rect 11270 13940 11280 14000
rect 11340 13940 11360 14000
rect 11420 13940 11440 14000
rect 11500 13940 11510 14000
rect 9420 13780 9480 13830
rect 9940 13780 10000 13830
rect 10460 13780 10520 13830
rect 9270 13760 9370 13780
rect 9270 13720 9320 13760
rect 9360 13720 9370 13760
rect 9270 13660 9370 13720
rect 9270 13620 9320 13660
rect 9360 13620 9370 13660
rect 9270 13600 9370 13620
rect 9420 13760 9520 13780
rect 9420 13720 9430 13760
rect 9470 13720 9520 13760
rect 9420 13660 9520 13720
rect 9420 13620 9430 13660
rect 9470 13620 9520 13660
rect 9420 13600 9520 13620
rect 9270 13400 9310 13600
rect 9366 13552 9424 13560
rect 9366 13500 9370 13552
rect 9422 13500 9424 13552
rect 9366 13490 9424 13500
rect 9480 13400 9520 13600
rect 9790 13760 9890 13780
rect 9790 13720 9840 13760
rect 9880 13720 9890 13760
rect 9790 13660 9890 13720
rect 9790 13620 9840 13660
rect 9880 13620 9890 13660
rect 9790 13600 9890 13620
rect 9940 13760 10040 13780
rect 9940 13720 9950 13760
rect 9990 13720 10040 13760
rect 9940 13660 10040 13720
rect 9940 13620 9950 13660
rect 9990 13620 10040 13660
rect 9940 13600 10040 13620
rect 9790 13400 9830 13600
rect 9886 13552 9944 13560
rect 9886 13500 9890 13552
rect 9942 13500 9944 13552
rect 9886 13490 9944 13500
rect 10000 13400 10040 13600
rect 10310 13760 10410 13780
rect 10310 13720 10360 13760
rect 10400 13720 10410 13760
rect 10310 13660 10410 13720
rect 10310 13620 10360 13660
rect 10400 13620 10410 13660
rect 10310 13600 10410 13620
rect 10460 13760 10560 13780
rect 10460 13720 10470 13760
rect 10510 13720 10560 13760
rect 10460 13660 10560 13720
rect 10460 13620 10470 13660
rect 10510 13620 10560 13660
rect 10460 13600 10560 13620
rect 10950 13760 11010 13830
rect 10950 13720 10960 13760
rect 11000 13720 11010 13760
rect 10950 13660 11010 13720
rect 10950 13620 10960 13660
rect 11000 13620 11010 13660
rect 10950 13600 11010 13620
rect 11060 13760 11120 13780
rect 11060 13720 11070 13760
rect 11110 13720 11120 13760
rect 11060 13660 11120 13720
rect 11060 13620 11070 13660
rect 11110 13620 11120 13660
rect 10310 13400 10350 13600
rect 10406 13552 10464 13560
rect 10406 13500 10410 13552
rect 10462 13500 10464 13552
rect 10406 13490 10464 13500
rect 10520 13400 10560 13600
rect 10974 13552 11032 13560
rect 10974 13500 10976 13552
rect 11028 13500 11032 13552
rect 10974 13490 11032 13500
rect 9270 13380 9370 13400
rect 9270 13340 9320 13380
rect 9360 13340 9370 13380
rect 9270 13280 9370 13340
rect 9270 13240 9320 13280
rect 9360 13240 9370 13280
rect 9270 13220 9370 13240
rect 9420 13390 9520 13400
rect 9480 13330 9520 13390
rect 9420 13290 9520 13330
rect 9480 13230 9520 13290
rect 9420 13220 9520 13230
rect 9620 13390 9700 13400
rect 9620 13330 9630 13390
rect 9690 13330 9700 13390
rect 9620 13290 9700 13330
rect 9620 13230 9630 13290
rect 9690 13230 9700 13290
rect 9270 13020 9310 13220
rect 9380 13172 9438 13180
rect 9380 13120 9384 13172
rect 9436 13120 9438 13172
rect 9380 13110 9438 13120
rect 9510 13170 9590 13180
rect 9510 13110 9520 13170
rect 9580 13110 9590 13170
rect 9510 13100 9590 13110
rect 9270 13000 9370 13020
rect 9270 12960 9320 13000
rect 9360 12960 9370 13000
rect 9270 12940 9370 12960
rect 9420 13000 9480 13020
rect 9420 12960 9430 13000
rect 9470 12960 9480 13000
rect 9420 12940 9480 12960
rect 9352 12882 9410 12900
rect 9352 12848 9364 12882
rect 9398 12848 9410 12882
rect 9352 12830 9410 12848
rect 9360 12770 9410 12830
rect 8920 12700 8930 12760
rect 8990 12700 9010 12760
rect 9070 12700 9090 12760
rect 9150 12700 9160 12760
rect 2340 12680 2420 12700
rect 8920 12690 9160 12700
rect 2340 12640 2360 12680
rect 2400 12640 2420 12680
rect 2340 12620 2420 12640
rect 8862 12680 9160 12690
rect 8862 12672 8930 12680
rect 8862 12620 8866 12672
rect 8918 12620 8930 12672
rect 8990 12620 9010 12680
rect 9070 12620 9090 12680
rect 9150 12620 9160 12680
rect 8862 12610 9160 12620
rect -1570 12600 -1490 12610
rect 8920 12600 9160 12610
rect 8920 12540 8930 12600
rect 8990 12540 9010 12600
rect 9070 12540 9090 12600
rect 9150 12540 9160 12600
rect 8920 12530 9160 12540
rect 9350 12760 9410 12770
rect 9350 12680 9410 12700
rect 9350 12600 9410 12620
rect 9350 12530 9410 12540
rect 840 12490 920 12510
rect 840 12450 860 12490
rect 900 12450 920 12490
rect 9360 12470 9410 12530
rect 840 12430 920 12450
rect 9352 12452 9410 12470
rect -560 12390 -480 12410
rect 840 12390 880 12430
rect 5260 12390 5300 12430
rect 6560 12390 6600 12430
rect 7860 12390 7900 12430
rect 9352 12418 9364 12452
rect 9398 12418 9410 12452
rect 9352 12400 9410 12418
rect 9440 12770 9480 12940
rect 9440 12760 9500 12770
rect 9440 12680 9500 12700
rect 9440 12600 9500 12620
rect 9440 12530 9500 12540
rect -870 12370 -600 12390
rect -870 12330 -850 12370
rect -810 12350 -660 12370
rect -810 12330 -790 12350
rect -870 12310 -790 12330
rect -670 12330 -660 12350
rect -620 12330 -600 12370
rect -560 12350 -540 12390
rect -500 12370 330 12390
rect -500 12350 270 12370
rect -560 12330 -480 12350
rect 250 12330 270 12350
rect 310 12330 330 12370
rect -670 12310 -600 12330
rect 250 12310 330 12330
rect 390 12370 880 12390
rect 390 12330 400 12370
rect 440 12350 880 12370
rect 1510 12370 1810 12390
rect 440 12330 450 12350
rect 390 12310 450 12330
rect 1510 12330 1530 12370
rect 1570 12350 1750 12370
rect 1570 12330 1590 12350
rect 1510 12310 1590 12330
rect 1730 12330 1750 12350
rect 1790 12330 1810 12370
rect 1730 12310 1810 12330
rect 2860 12360 3350 12380
rect 2860 12320 2880 12360
rect 2920 12340 3290 12360
rect 2920 12320 2940 12340
rect 2860 12310 2940 12320
rect 3270 12320 3290 12340
rect 3330 12320 3350 12360
rect 3270 12310 3350 12320
rect 5220 12370 5880 12390
rect 5220 12330 5240 12370
rect 5280 12350 5820 12370
rect 5280 12330 5300 12350
rect 5220 12310 5300 12330
rect 5800 12330 5820 12350
rect 5860 12330 5880 12370
rect 5800 12310 5880 12330
rect 6520 12370 7180 12390
rect 6520 12330 6540 12370
rect 6580 12350 7120 12370
rect 6580 12330 6600 12350
rect 6520 12310 6600 12330
rect 7100 12330 7120 12350
rect 7160 12330 7180 12370
rect 7100 12310 7180 12330
rect 7820 12370 8480 12390
rect 9440 12370 9480 12530
rect 7820 12330 7840 12370
rect 7880 12350 8420 12370
rect 7880 12330 7900 12350
rect 7820 12310 7900 12330
rect 8400 12330 8420 12350
rect 8460 12330 8480 12370
rect 8400 12310 8480 12330
rect 9310 12340 9370 12360
rect 9310 12300 9320 12340
rect 9360 12300 9370 12340
rect -1190 12270 -1110 12280
rect -1190 12210 -1180 12270
rect -1120 12210 -1110 12270
rect -1190 12200 -1110 12210
rect -770 12270 -690 12280
rect -770 12210 -760 12270
rect -700 12210 -690 12270
rect -770 12200 -690 12210
rect -100 12270 -20 12280
rect -100 12210 -90 12270
rect -30 12210 -20 12270
rect -100 12200 -20 12210
rect 470 12270 550 12280
rect 470 12210 480 12270
rect 540 12210 550 12270
rect 470 12200 550 12210
rect 1180 12270 1260 12280
rect 1180 12210 1190 12270
rect 1250 12210 1260 12270
rect 1180 12200 1260 12210
rect 1610 12270 1690 12280
rect 1610 12210 1620 12270
rect 1680 12210 1690 12270
rect 1610 12200 1690 12210
rect 2050 12270 2130 12280
rect 2050 12210 2060 12270
rect 2120 12210 2130 12270
rect 2050 12200 2130 12210
rect 2300 12270 2380 12280
rect 2300 12210 2310 12270
rect 2370 12210 2380 12270
rect 2300 12200 2380 12210
rect 2520 12270 2600 12280
rect 2520 12210 2530 12270
rect 2590 12210 2600 12270
rect 2520 12200 2600 12210
rect 2990 12270 3070 12280
rect 2990 12210 3000 12270
rect 3060 12210 3070 12270
rect 2990 12200 3070 12210
rect 3430 12270 3510 12280
rect 3430 12210 3440 12270
rect 3500 12210 3510 12270
rect 3430 12200 3510 12210
rect 4050 12270 4130 12280
rect 4050 12210 4060 12270
rect 4120 12210 4130 12270
rect 4050 12200 4130 12210
rect 4390 12270 4470 12280
rect 4390 12210 4400 12270
rect 4460 12210 4470 12270
rect 4390 12200 4470 12210
rect 4750 12270 4830 12280
rect 4750 12210 4760 12270
rect 4820 12210 4830 12270
rect 4750 12200 4830 12210
rect 5350 12270 5430 12280
rect 5350 12210 5360 12270
rect 5420 12210 5430 12270
rect 5350 12200 5430 12210
rect 5690 12270 5770 12280
rect 5690 12210 5700 12270
rect 5760 12210 5770 12270
rect 5690 12200 5770 12210
rect 6050 12270 6130 12280
rect 6050 12210 6060 12270
rect 6120 12210 6130 12270
rect 6050 12200 6130 12210
rect 6650 12270 6730 12280
rect 6650 12210 6660 12270
rect 6720 12210 6730 12270
rect 6650 12200 6730 12210
rect 6990 12270 7070 12280
rect 6990 12210 7000 12270
rect 7060 12210 7070 12270
rect 6990 12200 7070 12210
rect 7350 12270 7430 12280
rect 7350 12210 7360 12270
rect 7420 12210 7430 12270
rect 7350 12200 7430 12210
rect 7950 12270 8030 12280
rect 7950 12210 7960 12270
rect 8020 12210 8030 12270
rect 7950 12200 8030 12210
rect 8290 12270 8370 12280
rect 8290 12210 8300 12270
rect 8360 12210 8370 12270
rect 8290 12200 8370 12210
rect 8650 12270 8730 12280
rect 8650 12210 8660 12270
rect 8720 12210 8730 12270
rect 8650 12200 8730 12210
rect 9310 12240 9370 12300
rect 9310 12200 9320 12240
rect 9360 12200 9370 12240
rect 9310 12180 9370 12200
rect 9420 12340 9480 12370
rect 9420 12300 9430 12340
rect 9470 12300 9480 12340
rect 9420 12240 9480 12300
rect 9420 12200 9430 12240
rect 9470 12200 9480 12240
rect 9420 12180 9480 12200
rect 9310 11980 9350 12180
rect 9380 12082 9438 12090
rect 9380 12030 9384 12082
rect 9436 12030 9438 12082
rect 9380 12020 9438 12030
rect 9530 11980 9590 13100
rect 9620 12090 9700 13230
rect 9790 13380 9890 13400
rect 9790 13340 9840 13380
rect 9880 13340 9890 13380
rect 9790 13280 9890 13340
rect 9790 13240 9840 13280
rect 9880 13240 9890 13280
rect 9790 13220 9890 13240
rect 9940 13390 10040 13400
rect 10000 13330 10040 13390
rect 9940 13290 10040 13330
rect 10000 13230 10040 13290
rect 9940 13220 10040 13230
rect 10140 13390 10220 13400
rect 10140 13330 10150 13390
rect 10210 13330 10220 13390
rect 10140 13290 10220 13330
rect 10140 13230 10150 13290
rect 10210 13230 10220 13290
rect 9790 13020 9830 13220
rect 9900 13172 9958 13180
rect 9900 13120 9904 13172
rect 9956 13120 9958 13172
rect 9900 13110 9958 13120
rect 10030 13170 10110 13180
rect 10030 13110 10040 13170
rect 10100 13110 10110 13170
rect 10030 13100 10110 13110
rect 9790 13000 9890 13020
rect 9790 12960 9840 13000
rect 9880 12960 9890 13000
rect 9790 12940 9890 12960
rect 9940 13000 10000 13020
rect 9940 12960 9950 13000
rect 9990 12960 10000 13000
rect 9940 12940 10000 12960
rect 9872 12882 9930 12900
rect 9872 12848 9884 12882
rect 9918 12848 9930 12882
rect 9872 12830 9930 12848
rect 9880 12770 9930 12830
rect 9870 12760 9930 12770
rect 9870 12680 9930 12700
rect 9870 12600 9930 12620
rect 9870 12530 9930 12540
rect 9880 12470 9930 12530
rect 9872 12452 9930 12470
rect 9872 12418 9884 12452
rect 9918 12418 9930 12452
rect 9872 12400 9930 12418
rect 9960 12770 10000 12940
rect 9960 12760 10020 12770
rect 9960 12680 10020 12700
rect 9960 12600 10020 12620
rect 9960 12530 10020 12540
rect 9960 12370 10000 12530
rect 9620 12030 9630 12090
rect 9690 12030 9700 12090
rect 9620 12020 9700 12030
rect 9830 12340 9890 12360
rect 9830 12300 9840 12340
rect 9880 12300 9890 12340
rect 9830 12240 9890 12300
rect 9830 12200 9840 12240
rect 9880 12200 9890 12240
rect 9830 12180 9890 12200
rect 9940 12340 10000 12370
rect 9940 12300 9950 12340
rect 9990 12300 10000 12340
rect 9940 12240 10000 12300
rect 9940 12200 9950 12240
rect 9990 12200 10000 12240
rect 9940 12180 10000 12200
rect 9310 11960 9370 11980
rect 9310 11920 9320 11960
rect 9360 11920 9370 11960
rect 9310 11860 9370 11920
rect 9310 11820 9320 11860
rect 9360 11820 9370 11860
rect 9310 11760 9370 11820
rect 9310 11720 9320 11760
rect 9360 11720 9370 11760
rect 9310 11660 9370 11720
rect 9310 11620 9320 11660
rect 9360 11620 9370 11660
rect 9310 11270 9370 11620
rect 9420 11970 9480 11980
rect 9420 11860 9480 11910
rect 9510 11970 9590 11980
rect 9510 11910 9520 11970
rect 9580 11910 9590 11970
rect 9510 11900 9590 11910
rect 9830 11980 9870 12180
rect 9900 12082 9958 12090
rect 9900 12030 9904 12082
rect 9956 12030 9958 12082
rect 9900 12020 9958 12030
rect 10050 11980 10110 13100
rect 10140 12090 10220 13230
rect 10310 13380 10410 13400
rect 10310 13340 10360 13380
rect 10400 13340 10410 13380
rect 10310 13280 10410 13340
rect 10310 13240 10360 13280
rect 10400 13240 10410 13280
rect 10310 13220 10410 13240
rect 10460 13390 10560 13400
rect 10520 13330 10560 13390
rect 10460 13290 10560 13330
rect 10520 13230 10560 13290
rect 10460 13220 10560 13230
rect 10660 13390 10740 13400
rect 10660 13330 10670 13390
rect 10730 13330 10740 13390
rect 10660 13290 10740 13330
rect 10660 13230 10670 13290
rect 10730 13230 10740 13290
rect 10310 13020 10350 13220
rect 10420 13172 10478 13180
rect 10420 13120 10424 13172
rect 10476 13120 10478 13172
rect 10420 13110 10478 13120
rect 10550 13170 10630 13180
rect 10550 13110 10560 13170
rect 10620 13110 10630 13170
rect 10550 13100 10630 13110
rect 10310 13000 10410 13020
rect 10310 12960 10360 13000
rect 10400 12960 10410 13000
rect 10310 12940 10410 12960
rect 10460 13000 10520 13020
rect 10460 12960 10470 13000
rect 10510 12960 10520 13000
rect 10460 12940 10520 12960
rect 10392 12882 10450 12900
rect 10392 12848 10404 12882
rect 10438 12848 10450 12882
rect 10392 12830 10450 12848
rect 10400 12770 10450 12830
rect 10390 12760 10450 12770
rect 10390 12680 10450 12700
rect 10390 12600 10450 12620
rect 10390 12530 10450 12540
rect 10400 12470 10450 12530
rect 10392 12452 10450 12470
rect 10392 12418 10404 12452
rect 10438 12418 10450 12452
rect 10392 12400 10450 12418
rect 10480 12770 10520 12940
rect 10480 12760 10540 12770
rect 10480 12680 10540 12700
rect 10480 12600 10540 12620
rect 10480 12530 10540 12540
rect 10480 12370 10520 12530
rect 10140 12030 10150 12090
rect 10210 12030 10220 12090
rect 10140 12020 10220 12030
rect 10350 12340 10410 12360
rect 10350 12300 10360 12340
rect 10400 12300 10410 12340
rect 10350 12240 10410 12300
rect 10350 12200 10360 12240
rect 10400 12200 10410 12240
rect 10350 12180 10410 12200
rect 10460 12340 10520 12370
rect 10460 12300 10470 12340
rect 10510 12300 10520 12340
rect 10460 12240 10520 12300
rect 10460 12200 10470 12240
rect 10510 12200 10520 12240
rect 10460 12180 10520 12200
rect 9830 11960 9890 11980
rect 9830 11920 9840 11960
rect 9880 11920 9890 11960
rect 9420 11820 9430 11860
rect 9470 11820 9480 11860
rect 9420 11760 9480 11820
rect 9420 11720 9430 11760
rect 9470 11720 9480 11760
rect 9420 11660 9480 11720
rect 9420 11620 9430 11660
rect 9470 11620 9480 11660
rect 9420 11590 9480 11620
rect 9830 11860 9890 11920
rect 9830 11820 9840 11860
rect 9880 11820 9890 11860
rect 9830 11760 9890 11820
rect 9830 11720 9840 11760
rect 9880 11720 9890 11760
rect 9830 11660 9890 11720
rect 9830 11620 9840 11660
rect 9880 11620 9890 11660
rect 9410 11580 9490 11590
rect 9410 11520 9420 11580
rect 9480 11520 9490 11580
rect 9410 11510 9490 11520
rect 9680 11580 9760 11590
rect 9680 11520 9690 11580
rect 9750 11520 9760 11580
rect 9680 11510 9760 11520
rect 9490 11400 9570 11410
rect 9490 11340 9500 11400
rect 9560 11340 9570 11400
rect 9490 11330 9570 11340
rect 9310 11230 9320 11270
rect 9360 11230 9370 11270
rect 9310 11170 9370 11230
rect 9310 11130 9320 11170
rect 9360 11130 9370 11170
rect 9310 11070 9370 11130
rect 9310 11030 9320 11070
rect 9360 11030 9370 11070
rect 9310 10970 9370 11030
rect 9310 10930 9320 10970
rect 9360 10930 9370 10970
rect 9310 10910 9370 10930
rect 9690 11270 9750 11510
rect 9690 11230 9700 11270
rect 9740 11230 9750 11270
rect 9690 11170 9750 11230
rect 9690 11130 9700 11170
rect 9740 11130 9750 11170
rect 9690 11070 9750 11130
rect 9690 11030 9700 11070
rect 9740 11030 9750 11070
rect 9690 10970 9750 11030
rect 9690 10930 9700 10970
rect 9740 10930 9750 10970
rect 9690 10860 9750 10930
rect 9830 11270 9890 11620
rect 9940 11970 10000 11980
rect 9940 11860 10000 11910
rect 10030 11970 10110 11980
rect 10030 11910 10040 11970
rect 10100 11910 10110 11970
rect 10030 11900 10110 11910
rect 10350 11980 10390 12180
rect 10420 12082 10478 12090
rect 10420 12030 10424 12082
rect 10476 12030 10478 12082
rect 10420 12020 10478 12030
rect 10570 11980 10630 13100
rect 10660 12090 10740 13230
rect 10660 12030 10670 12090
rect 10730 12030 10740 12090
rect 10660 12020 10740 12030
rect 10350 11960 10410 11980
rect 10350 11920 10360 11960
rect 10400 11920 10410 11960
rect 9940 11820 9950 11860
rect 9990 11820 10000 11860
rect 9940 11760 10000 11820
rect 9940 11720 9950 11760
rect 9990 11720 10000 11760
rect 9940 11660 10000 11720
rect 9940 11620 9950 11660
rect 9990 11620 10000 11660
rect 9940 11590 10000 11620
rect 10350 11860 10410 11920
rect 10350 11820 10360 11860
rect 10400 11820 10410 11860
rect 10350 11760 10410 11820
rect 10350 11720 10360 11760
rect 10400 11720 10410 11760
rect 10350 11660 10410 11720
rect 10350 11620 10360 11660
rect 10400 11620 10410 11660
rect 9930 11580 10010 11590
rect 9930 11520 9940 11580
rect 10000 11520 10010 11580
rect 9930 11510 10010 11520
rect 10200 11580 10280 11590
rect 10200 11520 10210 11580
rect 10270 11520 10280 11580
rect 10200 11510 10280 11520
rect 10010 11400 10090 11410
rect 10010 11340 10020 11400
rect 10080 11340 10090 11400
rect 10010 11330 10090 11340
rect 9830 11230 9840 11270
rect 9880 11230 9890 11270
rect 9830 11170 9890 11230
rect 9830 11130 9840 11170
rect 9880 11130 9890 11170
rect 9830 11070 9890 11130
rect 9830 11030 9840 11070
rect 9880 11030 9890 11070
rect 9830 10970 9890 11030
rect 9830 10930 9840 10970
rect 9880 10930 9890 10970
rect 9830 10910 9890 10930
rect 10210 11270 10270 11510
rect 10210 11230 10220 11270
rect 10260 11230 10270 11270
rect 10210 11170 10270 11230
rect 10210 11130 10220 11170
rect 10260 11130 10270 11170
rect 10210 11070 10270 11130
rect 10210 11030 10220 11070
rect 10260 11030 10270 11070
rect 10210 10970 10270 11030
rect 10210 10930 10220 10970
rect 10260 10930 10270 10970
rect 10210 10860 10270 10930
rect 10350 11270 10410 11620
rect 10460 11970 10520 11980
rect 10460 11860 10520 11910
rect 10550 11970 10630 11980
rect 10550 11910 10560 11970
rect 10620 11910 10630 11970
rect 10550 11900 10630 11910
rect 10460 11820 10470 11860
rect 10510 11820 10520 11860
rect 10460 11760 10520 11820
rect 10460 11720 10470 11760
rect 10510 11720 10520 11760
rect 10460 11660 10520 11720
rect 10460 11620 10470 11660
rect 10510 11620 10520 11660
rect 10460 11590 10520 11620
rect 10450 11580 10530 11590
rect 10450 11520 10460 11580
rect 10520 11520 10530 11580
rect 10450 11510 10530 11520
rect 10720 11580 10800 11590
rect 10720 11520 10730 11580
rect 10790 11520 10800 11580
rect 10720 11510 10800 11520
rect 10530 11400 10610 11410
rect 10530 11340 10540 11400
rect 10600 11340 10610 11400
rect 10530 11330 10610 11340
rect 10350 11230 10360 11270
rect 10400 11230 10410 11270
rect 10350 11170 10410 11230
rect 10350 11130 10360 11170
rect 10400 11130 10410 11170
rect 10350 11070 10410 11130
rect 10350 11030 10360 11070
rect 10400 11030 10410 11070
rect 10350 10970 10410 11030
rect 10350 10930 10360 10970
rect 10400 10930 10410 10970
rect 10350 10910 10410 10930
rect 10730 11270 10790 11510
rect 10730 11230 10740 11270
rect 10780 11230 10790 11270
rect 10730 11170 10790 11230
rect 10730 11130 10740 11170
rect 10780 11130 10790 11170
rect 10730 11070 10790 11130
rect 10730 11030 10740 11070
rect 10780 11030 10790 11070
rect 10730 10970 10790 11030
rect 10730 10930 10740 10970
rect 10780 10930 10790 10970
rect 10730 10860 10790 10930
rect 10870 11400 10930 11410
rect 10870 11270 10930 11340
rect 11060 11400 11120 13620
rect 11270 12760 11510 13940
rect 11270 12700 11280 12760
rect 11340 12700 11360 12760
rect 11420 12700 11440 12760
rect 11500 12700 11510 12760
rect 11270 12680 11510 12700
rect 11270 12620 11280 12680
rect 11340 12620 11360 12680
rect 11420 12620 11440 12680
rect 11500 12620 11510 12680
rect 11270 12600 11510 12620
rect 11270 12540 11280 12600
rect 11340 12540 11360 12600
rect 11420 12540 11440 12600
rect 11500 12540 11510 12600
rect 11270 12530 11510 12540
rect 12110 13550 12190 13560
rect 12110 13490 12120 13550
rect 12180 13490 12190 13550
rect 11060 11330 11120 11340
rect 10870 11230 10880 11270
rect 10920 11230 10930 11270
rect 10870 11170 10930 11230
rect 10870 11130 10880 11170
rect 10920 11130 10930 11170
rect 10870 11070 10930 11130
rect 10870 11030 10880 11070
rect 10920 11030 10930 11070
rect 10870 10970 10930 11030
rect 10870 10930 10880 10970
rect 10920 10930 10930 10970
rect 10870 10910 10930 10930
rect 11250 11270 11310 11290
rect 11250 11230 11260 11270
rect 11300 11230 11310 11270
rect 11250 11170 11310 11230
rect 11250 11130 11260 11170
rect 11300 11130 11310 11170
rect 11250 11070 11310 11130
rect 11250 11030 11260 11070
rect 11300 11030 11310 11070
rect 11250 10970 11310 11030
rect 11250 10930 11260 10970
rect 11300 10930 11310 10970
rect 11250 10860 11310 10930
rect 9680 10840 9760 10860
rect 9680 10800 9700 10840
rect 9740 10800 9760 10840
rect 9680 10750 9760 10800
rect 9680 10690 9690 10750
rect 9750 10690 9760 10750
rect 9680 10680 9760 10690
rect 10200 10840 10280 10860
rect 10200 10800 10220 10840
rect 10260 10800 10280 10840
rect 10200 10750 10280 10800
rect 10200 10690 10210 10750
rect 10270 10690 10280 10750
rect 10200 10680 10280 10690
rect 10720 10840 10800 10860
rect 10720 10800 10740 10840
rect 10780 10800 10800 10840
rect 10720 10750 10800 10800
rect 10720 10690 10730 10750
rect 10790 10690 10800 10750
rect 10720 10680 10800 10690
rect 11240 10840 11320 10860
rect 11240 10800 11260 10840
rect 11300 10800 11320 10840
rect 11240 10750 11320 10800
rect 11240 10690 11250 10750
rect 11310 10690 11320 10750
rect 11240 10680 11320 10690
rect 9090 10520 9200 10540
rect 3800 10510 3880 10520
rect -640 10450 -560 10460
rect -640 10390 -630 10450
rect -570 10390 -560 10450
rect -640 10380 -560 10390
rect -420 10450 -340 10460
rect -420 10390 -410 10450
rect -350 10390 -340 10450
rect -420 10380 -340 10390
rect -120 10450 -40 10460
rect -120 10390 -110 10450
rect -50 10390 -40 10450
rect -120 10380 -40 10390
rect 100 10450 180 10460
rect 100 10390 110 10450
rect 170 10390 180 10450
rect 100 10380 180 10390
rect 260 10450 340 10460
rect 260 10390 270 10450
rect 330 10390 340 10450
rect 260 10380 340 10390
rect 480 10450 560 10460
rect 480 10390 490 10450
rect 550 10390 560 10450
rect 480 10380 560 10390
rect 780 10450 860 10460
rect 780 10390 790 10450
rect 850 10390 860 10450
rect 780 10380 860 10390
rect 1000 10450 1080 10460
rect 1000 10390 1010 10450
rect 1070 10390 1080 10450
rect 1000 10380 1080 10390
rect 1300 10450 1380 10460
rect 1300 10390 1310 10450
rect 1370 10390 1380 10450
rect 1300 10380 1380 10390
rect 1740 10450 1820 10460
rect 1740 10390 1750 10450
rect 1810 10390 1820 10450
rect 1740 10380 1820 10390
rect 2070 10450 2150 10460
rect 2070 10390 2080 10450
rect 2140 10390 2150 10450
rect 2070 10380 2150 10390
rect 2500 10450 2580 10460
rect 2500 10390 2510 10450
rect 2570 10390 2580 10450
rect 2500 10380 2580 10390
rect 2890 10450 2970 10460
rect 2890 10390 2900 10450
rect 2960 10390 2970 10450
rect 2890 10380 2970 10390
rect 3280 10450 3360 10460
rect 3280 10390 3290 10450
rect 3350 10390 3360 10450
rect 3280 10380 3360 10390
rect 3800 10450 3810 10510
rect 3870 10450 3880 10510
rect -230 10340 -150 10350
rect -230 10280 -220 10340
rect -160 10280 -150 10340
rect -230 10270 -150 10280
rect 1490 10340 1570 10350
rect 1490 10280 1500 10340
rect 1560 10280 1570 10340
rect 3570 10340 3650 10350
rect 1490 10270 1570 10280
rect 2340 10320 2420 10330
rect 2340 10260 2350 10320
rect 2410 10260 2420 10320
rect 3570 10280 3580 10340
rect 3640 10280 3650 10340
rect 3570 10270 3650 10280
rect 2340 10250 2420 10260
rect 1140 9990 1220 10000
rect -760 9960 -680 9970
rect -760 9900 -750 9960
rect -690 9900 -680 9960
rect 1140 9930 1150 9990
rect 1210 9930 1220 9990
rect 2360 9990 2400 10250
rect 2360 9970 2440 9990
rect 1140 9920 1220 9930
rect -760 9890 -680 9900
rect -640 9270 -560 9280
rect -640 9210 -630 9270
rect -570 9210 -560 9270
rect -640 9200 -560 9210
rect 100 9270 180 9280
rect 100 9210 110 9270
rect 170 9210 180 9270
rect 100 9200 180 9210
rect 260 9270 340 9280
rect 260 9210 270 9270
rect 330 9210 340 9270
rect 260 9200 340 9210
rect 1000 9270 1080 9280
rect 1000 9210 1010 9270
rect 1070 9210 1080 9270
rect 1000 9200 1080 9210
rect -190 9160 -110 9170
rect -190 9100 -180 9160
rect -120 9100 -110 9160
rect -190 9090 -110 9100
rect 1180 8600 1220 9920
rect 2230 9950 2310 9960
rect 2230 9890 2240 9950
rect 2300 9890 2310 9950
rect 2360 9930 2380 9970
rect 2420 9930 2440 9970
rect 2360 9910 2440 9930
rect 3800 9920 3880 10450
rect 9090 10450 9110 10520
rect 9180 10450 9200 10520
rect 9090 10430 9200 10450
rect 4510 10340 4590 10350
rect 4510 10280 4520 10340
rect 4580 10280 4590 10340
rect 4110 10000 4190 10010
rect 4110 9940 4120 10000
rect 4180 9940 4190 10000
rect 4110 9930 4190 9940
rect 4400 10000 4480 10010
rect 4400 9940 4410 10000
rect 4470 9940 4480 10000
rect 2230 9880 2310 9890
rect 1360 9380 1440 9390
rect 1360 9320 1370 9380
rect 1430 9320 1440 9380
rect 1250 9270 1330 9280
rect 1250 9210 1260 9270
rect 1320 9210 1330 9270
rect 1250 9200 1330 9210
rect 1360 9170 1400 9320
rect 1440 9270 1600 9280
rect 1440 9210 1450 9270
rect 1510 9210 1530 9270
rect 1590 9210 1600 9270
rect 1440 9200 1600 9210
rect 1730 9270 1810 9280
rect 1730 9210 1740 9270
rect 1800 9210 1810 9270
rect 1730 9200 1810 9210
rect 2060 9270 2140 9280
rect 2060 9210 2070 9270
rect 2130 9210 2140 9270
rect 2060 9200 2140 9210
rect 1340 9160 1420 9170
rect 1340 9100 1350 9160
rect 1410 9100 1420 9160
rect 1340 9090 1420 9100
rect 2270 8600 2310 9880
rect 3800 9860 3810 9920
rect 3870 9860 3880 9920
rect 3800 9850 3880 9860
rect 2500 9270 2580 9280
rect 2500 9210 2510 9270
rect 2570 9210 2580 9270
rect 2500 9200 2580 9210
rect 2890 9270 2970 9280
rect 2890 9210 2900 9270
rect 2960 9210 2970 9270
rect 2890 9200 2970 9210
rect 3100 9270 3180 9280
rect 3100 9210 3110 9270
rect 3170 9210 3180 9270
rect 3100 9200 3180 9210
rect 3280 9270 3360 9280
rect 3280 9210 3290 9270
rect 3350 9210 3360 9270
rect 3280 9200 3360 9210
rect 3960 9270 4040 9280
rect 3960 9210 3970 9270
rect 4030 9210 4040 9270
rect 3960 9200 4040 9210
rect 1160 8590 1240 8600
rect -1780 8520 -1770 8580
rect -1710 8520 -1700 8580
rect -1780 8510 -1700 8520
rect -760 8580 -680 8590
rect -760 8520 -750 8580
rect -690 8520 -680 8580
rect 1160 8530 1170 8590
rect 1230 8530 1240 8590
rect 1160 8520 1240 8530
rect 2190 8590 2310 8600
rect 2190 8530 2200 8590
rect 2260 8530 2310 8590
rect 2190 8520 2310 8530
rect 2340 9150 2420 9160
rect 2340 9090 2350 9150
rect 2410 9090 2420 9150
rect 2760 9100 2770 9160
rect 2830 9100 2840 9160
rect 2930 9100 2940 9160
rect 3000 9100 3010 9160
rect 2340 9080 2420 9090
rect 2340 8590 2380 9080
rect 2340 8570 2420 8590
rect 2340 8530 2360 8570
rect 2400 8530 2420 8570
rect -760 8510 -680 8520
rect 2340 8510 2420 8530
rect 2780 8100 2820 9100
rect 2930 9090 3010 9100
rect 3120 8210 3160 9200
rect 3570 9160 3650 9170
rect 3570 9100 3580 9160
rect 3640 9100 3650 9160
rect 3570 9090 3650 9100
rect 4290 9160 4370 9170
rect 4290 9100 4300 9160
rect 4360 9100 4370 9160
rect 4290 9010 4370 9100
rect 4400 9120 4480 9940
rect 4510 9230 4590 10280
rect 5650 10000 5730 10010
rect 5650 9940 5660 10000
rect 5720 9940 5730 10000
rect 5650 9880 5730 9940
rect 5650 9840 5670 9880
rect 5710 9840 5730 9880
rect 5650 9760 5730 9840
rect 5650 9720 5670 9760
rect 5710 9720 5730 9760
rect 5650 9660 5730 9720
rect 5650 9620 5670 9660
rect 5710 9620 5730 9660
rect 5650 9560 5730 9620
rect 5650 9520 5670 9560
rect 5710 9520 5730 9560
rect 5650 9460 5730 9520
rect 5650 9420 5670 9460
rect 5710 9420 5730 9460
rect 5650 9400 5730 9420
rect 5870 10000 5950 10010
rect 5870 9940 5880 10000
rect 5940 9940 5950 10000
rect 5870 9760 5950 9940
rect 6310 10000 6390 10010
rect 6310 9940 6320 10000
rect 6380 9940 6390 10000
rect 5870 9720 5890 9760
rect 5930 9720 5950 9760
rect 5870 9660 5950 9720
rect 5870 9620 5890 9660
rect 5930 9620 5950 9660
rect 5870 9560 5950 9620
rect 5870 9520 5890 9560
rect 5930 9520 5950 9560
rect 5870 9460 5950 9520
rect 5870 9420 5890 9460
rect 5930 9420 5950 9460
rect 5870 9400 5950 9420
rect 6090 9760 6170 9780
rect 6090 9720 6110 9760
rect 6150 9720 6170 9760
rect 6090 9660 6170 9720
rect 6090 9620 6110 9660
rect 6150 9620 6170 9660
rect 6090 9560 6170 9620
rect 6090 9520 6110 9560
rect 6150 9520 6170 9560
rect 6090 9460 6170 9520
rect 6090 9420 6110 9460
rect 6150 9420 6170 9460
rect 4510 9170 4520 9230
rect 4580 9170 4590 9230
rect 4510 9160 4590 9170
rect 5030 9350 5110 9360
rect 5030 9290 5040 9350
rect 5100 9290 5110 9350
rect 4400 9060 4410 9120
rect 4470 9060 4480 9120
rect 4400 9050 4480 9060
rect 4290 8950 4300 9010
rect 4360 8950 4370 9010
rect 4290 8940 4370 8950
rect 4760 9010 5000 9020
rect 4760 8950 4770 9010
rect 4830 8950 4850 9010
rect 4910 8950 4930 9010
rect 4990 8950 5000 9010
rect 4290 8900 4370 8910
rect 4290 8840 4300 8900
rect 4360 8840 4370 8900
rect 4110 8540 4190 8550
rect 4110 8480 4120 8540
rect 4180 8480 4190 8540
rect 4110 8470 4190 8480
rect 4290 8540 4370 8840
rect 4290 8480 4300 8540
rect 4360 8480 4370 8540
rect 4290 8470 4370 8480
rect 3010 8200 3160 8210
rect 3010 8140 3020 8200
rect 3080 8140 3160 8200
rect 3010 8130 3160 8140
rect 3640 8200 3720 8210
rect 3640 8140 3650 8200
rect 3710 8140 3720 8200
rect 3640 8130 3720 8140
rect 4210 8200 4290 8210
rect 4210 8140 4220 8200
rect 4280 8140 4290 8200
rect -640 8090 -560 8100
rect -640 8030 -630 8090
rect -570 8030 -560 8090
rect -640 8020 -560 8030
rect -420 8090 -340 8100
rect -420 8030 -410 8090
rect -350 8030 -340 8090
rect -420 8020 -340 8030
rect -120 8090 -40 8100
rect -120 8030 -110 8090
rect -50 8030 -40 8090
rect -120 8020 -40 8030
rect 110 8090 190 8100
rect 110 8030 120 8090
rect 180 8030 190 8090
rect 110 8020 190 8030
rect 260 8090 340 8100
rect 260 8030 270 8090
rect 330 8030 340 8090
rect 260 8020 340 8030
rect 480 8090 560 8100
rect 480 8030 490 8090
rect 550 8030 560 8090
rect 480 8020 560 8030
rect 780 8090 860 8100
rect 780 8030 790 8090
rect 850 8030 860 8090
rect 780 8020 860 8030
rect 1000 8090 1080 8100
rect 1000 8030 1010 8090
rect 1070 8030 1080 8090
rect 1000 8020 1080 8030
rect 1400 8090 1480 8100
rect 1400 8030 1410 8090
rect 1470 8030 1480 8090
rect 1400 8020 1480 8030
rect 1730 8090 1810 8100
rect 1730 8030 1740 8090
rect 1800 8030 1810 8090
rect 1730 8020 1810 8030
rect 2060 8090 2140 8100
rect 2060 8030 2070 8090
rect 2130 8030 2140 8090
rect 2060 8020 2140 8030
rect 2500 8090 2580 8100
rect 2500 8030 2510 8090
rect 2570 8030 2580 8090
rect 2500 8020 2580 8030
rect 2760 8090 2840 8100
rect 2760 8030 2770 8090
rect 2830 8030 2840 8090
rect 2760 8020 2840 8030
rect 3280 8090 3360 8100
rect 3280 8030 3290 8090
rect 3350 8030 3360 8090
rect 3280 8020 3360 8030
rect 3960 8090 4040 8100
rect 3960 8030 3970 8090
rect 4030 8030 4040 8090
rect 3960 8020 4040 8030
rect 4210 8020 4290 8140
rect 4210 7960 4220 8020
rect 4280 7960 4290 8020
rect 4210 7950 4290 7960
rect 650 7250 730 7260
rect 650 7190 660 7250
rect 720 7190 730 7250
rect 650 7170 730 7190
rect 650 7110 660 7170
rect 720 7110 730 7170
rect 650 7090 730 7110
rect -2640 7080 -2560 7090
rect -2640 7020 -2630 7080
rect -2570 7020 -2560 7080
rect -2870 6630 -2790 6640
rect -2870 6570 -2860 6630
rect -2800 6570 -2790 6630
rect -2980 5300 -2900 5310
rect -2980 5240 -2970 5300
rect -2910 5240 -2900 5300
rect -2980 2180 -2900 5240
rect -2980 2120 -2970 2180
rect -2910 2120 -2900 2180
rect -2980 2110 -2900 2120
rect -2870 4810 -2790 6570
rect -2870 4750 -2860 4810
rect -2800 4750 -2790 4810
rect -2870 -440 -2790 4750
rect -2750 5190 -2670 5200
rect -2750 5130 -2740 5190
rect -2680 5130 -2670 5190
rect -2750 3870 -2670 5130
rect -2750 3810 -2740 3870
rect -2680 3810 -2670 3870
rect -2750 -386 -2670 3810
rect -2640 3640 -2560 7020
rect -1250 7080 -1170 7090
rect -1250 7020 -1240 7080
rect -1180 7020 -1170 7080
rect -1250 7010 -1170 7020
rect -1030 7080 -950 7090
rect -1030 7020 -1020 7080
rect -960 7020 -950 7080
rect -1030 7010 -950 7020
rect -810 7080 -730 7090
rect -810 7020 -800 7080
rect -740 7020 -730 7080
rect -810 7010 -730 7020
rect -590 7080 -510 7090
rect -590 7020 -580 7080
rect -520 7020 -510 7080
rect -590 7010 -510 7020
rect -370 7080 -290 7090
rect -370 7020 -360 7080
rect -300 7020 -290 7080
rect -370 7010 -290 7020
rect -150 7080 -70 7090
rect -150 7020 -140 7080
rect -80 7020 -70 7080
rect 650 7030 660 7090
rect 720 7030 730 7090
rect 650 7020 730 7030
rect 870 7250 950 7260
rect 870 7190 880 7250
rect 940 7190 950 7250
rect 870 7170 950 7190
rect 870 7110 880 7170
rect 940 7110 950 7170
rect 870 7090 950 7110
rect 870 7030 880 7090
rect 940 7030 950 7090
rect 870 7020 950 7030
rect 1090 7250 1170 7260
rect 1090 7190 1100 7250
rect 1160 7190 1170 7250
rect 1090 7170 1170 7190
rect 1090 7110 1100 7170
rect 1160 7110 1170 7170
rect 1090 7090 1170 7110
rect 1090 7030 1100 7090
rect 1160 7030 1170 7090
rect 1090 7020 1170 7030
rect 1310 7250 1390 7260
rect 1310 7190 1320 7250
rect 1380 7190 1390 7250
rect 1310 7170 1390 7190
rect 1310 7110 1320 7170
rect 1380 7110 1390 7170
rect 1310 7090 1390 7110
rect 1310 7030 1320 7090
rect 1380 7030 1390 7090
rect 1310 7020 1390 7030
rect 1530 7250 1610 7260
rect 1530 7190 1540 7250
rect 1600 7190 1610 7250
rect 1530 7170 1610 7190
rect 1530 7110 1540 7170
rect 1600 7110 1610 7170
rect 1530 7090 1610 7110
rect 1530 7030 1540 7090
rect 1600 7030 1610 7090
rect 1530 7020 1610 7030
rect 1750 7250 1830 7260
rect 1750 7190 1760 7250
rect 1820 7190 1830 7250
rect 1750 7170 1830 7190
rect 1750 7110 1760 7170
rect 1820 7110 1830 7170
rect 1750 7090 1830 7110
rect 1750 7030 1760 7090
rect 1820 7030 1830 7090
rect 1750 7020 1830 7030
rect 4760 7250 5000 8950
rect 4760 7190 4770 7250
rect 4830 7190 4850 7250
rect 4910 7190 4930 7250
rect 4990 7190 5000 7250
rect 4760 7170 5000 7190
rect 4760 7110 4770 7170
rect 4830 7110 4850 7170
rect 4910 7110 4930 7170
rect 4990 7110 5000 7170
rect 4760 7090 5000 7110
rect 4760 7030 4770 7090
rect 4830 7030 4850 7090
rect 4910 7030 4930 7090
rect 4990 7030 5000 7090
rect 4760 7020 5000 7030
rect -150 7010 -70 7020
rect -1360 6970 -1280 6980
rect -1360 6910 -1350 6970
rect -1290 6910 -1280 6970
rect -1360 6900 -1280 6910
rect -1350 6860 -1290 6900
rect -1430 6840 -1290 6860
rect -1430 6800 -1420 6840
rect -1380 6800 -1340 6840
rect -1300 6800 -1290 6840
rect -1430 6740 -1290 6800
rect -1430 6700 -1420 6740
rect -1380 6700 -1340 6740
rect -1300 6700 -1290 6740
rect -1430 6680 -1290 6700
rect -1240 6840 -1180 7010
rect -1140 6970 -1060 6980
rect -1140 6910 -1130 6970
rect -1070 6910 -1060 6970
rect -1140 6900 -1060 6910
rect -1240 6800 -1230 6840
rect -1190 6800 -1180 6840
rect -1240 6740 -1180 6800
rect -1240 6700 -1230 6740
rect -1190 6700 -1180 6740
rect -1240 6680 -1180 6700
rect -1130 6840 -1070 6900
rect -1130 6800 -1120 6840
rect -1080 6800 -1070 6840
rect -1130 6740 -1070 6800
rect -1130 6700 -1120 6740
rect -1080 6700 -1070 6740
rect -1130 6680 -1070 6700
rect -1020 6840 -960 7010
rect -920 6970 -840 6980
rect -920 6910 -910 6970
rect -850 6910 -840 6970
rect -920 6900 -840 6910
rect -1020 6800 -1010 6840
rect -970 6800 -960 6840
rect -1020 6740 -960 6800
rect -1020 6700 -1010 6740
rect -970 6700 -960 6740
rect -1020 6680 -960 6700
rect -910 6840 -850 6900
rect -910 6800 -900 6840
rect -860 6800 -850 6840
rect -910 6740 -850 6800
rect -910 6700 -900 6740
rect -860 6700 -850 6740
rect -910 6680 -850 6700
rect -800 6840 -740 7010
rect -700 6970 -620 6980
rect -700 6910 -690 6970
rect -630 6910 -620 6970
rect -700 6900 -620 6910
rect -800 6800 -790 6840
rect -750 6800 -740 6840
rect -800 6740 -740 6800
rect -800 6700 -790 6740
rect -750 6700 -740 6740
rect -800 6680 -740 6700
rect -690 6840 -630 6900
rect -690 6800 -680 6840
rect -640 6800 -630 6840
rect -690 6740 -630 6800
rect -690 6700 -680 6740
rect -640 6700 -630 6740
rect -690 6680 -630 6700
rect -580 6840 -520 7010
rect -480 6970 -400 6980
rect -480 6910 -470 6970
rect -410 6910 -400 6970
rect -480 6900 -400 6910
rect -580 6800 -570 6840
rect -530 6800 -520 6840
rect -580 6740 -520 6800
rect -580 6700 -570 6740
rect -530 6700 -520 6740
rect -580 6680 -520 6700
rect -470 6840 -410 6900
rect -470 6800 -460 6840
rect -420 6800 -410 6840
rect -470 6740 -410 6800
rect -470 6700 -460 6740
rect -420 6700 -410 6740
rect -470 6680 -410 6700
rect -360 6840 -300 7010
rect -260 6970 -180 6980
rect -260 6910 -250 6970
rect -190 6910 -180 6970
rect -260 6900 -180 6910
rect -360 6800 -350 6840
rect -310 6800 -300 6840
rect -360 6740 -300 6800
rect -360 6700 -350 6740
rect -310 6700 -300 6740
rect -360 6680 -300 6700
rect -250 6840 -190 6900
rect -250 6800 -240 6840
rect -200 6800 -190 6840
rect -250 6740 -190 6800
rect -250 6700 -240 6740
rect -200 6700 -190 6740
rect -250 6680 -190 6700
rect -140 6840 -80 7010
rect -40 6970 40 6980
rect -40 6910 -30 6970
rect 30 6910 40 6970
rect -40 6900 40 6910
rect 540 6970 620 6980
rect 540 6910 550 6970
rect 610 6910 620 6970
rect 540 6900 620 6910
rect -140 6800 -130 6840
rect -90 6800 -80 6840
rect -140 6740 -80 6800
rect -140 6700 -130 6740
rect -90 6700 -80 6740
rect -140 6680 -80 6700
rect -30 6860 30 6900
rect 550 6860 610 6900
rect -30 6840 110 6860
rect -30 6800 -20 6840
rect 20 6800 60 6840
rect 100 6800 110 6840
rect -30 6740 110 6800
rect -30 6700 -20 6740
rect 20 6700 60 6740
rect 100 6700 110 6740
rect -30 6680 110 6700
rect 470 6840 610 6860
rect 470 6800 480 6840
rect 520 6800 560 6840
rect 600 6800 610 6840
rect 470 6740 610 6800
rect 470 6700 480 6740
rect 520 6700 560 6740
rect 600 6700 610 6740
rect 470 6680 610 6700
rect 660 6840 720 7020
rect 760 6970 840 6980
rect 760 6910 770 6970
rect 830 6910 840 6970
rect 760 6900 840 6910
rect 660 6800 670 6840
rect 710 6800 720 6840
rect 660 6740 720 6800
rect 660 6700 670 6740
rect 710 6700 720 6740
rect 660 6680 720 6700
rect 770 6840 830 6900
rect 770 6800 780 6840
rect 820 6800 830 6840
rect 770 6740 830 6800
rect 770 6700 780 6740
rect 820 6700 830 6740
rect 770 6680 830 6700
rect 880 6840 940 7020
rect 980 6970 1060 6980
rect 980 6910 990 6970
rect 1050 6910 1060 6970
rect 980 6900 1060 6910
rect 880 6800 890 6840
rect 930 6800 940 6840
rect 880 6740 940 6800
rect 880 6700 890 6740
rect 930 6700 940 6740
rect 880 6680 940 6700
rect 990 6840 1050 6900
rect 990 6800 1000 6840
rect 1040 6800 1050 6840
rect 990 6740 1050 6800
rect 990 6700 1000 6740
rect 1040 6700 1050 6740
rect 990 6680 1050 6700
rect 1100 6840 1160 7020
rect 1200 6970 1280 6980
rect 1200 6910 1210 6970
rect 1270 6910 1280 6970
rect 1200 6900 1280 6910
rect 1100 6800 1110 6840
rect 1150 6800 1160 6840
rect 1100 6740 1160 6800
rect 1100 6700 1110 6740
rect 1150 6700 1160 6740
rect 1100 6680 1160 6700
rect 1210 6840 1270 6900
rect 1210 6800 1220 6840
rect 1260 6800 1270 6840
rect 1210 6740 1270 6800
rect 1210 6700 1220 6740
rect 1260 6700 1270 6740
rect 1210 6680 1270 6700
rect 1320 6840 1380 7020
rect 1420 6970 1500 6980
rect 1420 6910 1430 6970
rect 1490 6910 1500 6970
rect 1420 6900 1500 6910
rect 1320 6800 1330 6840
rect 1370 6800 1380 6840
rect 1320 6740 1380 6800
rect 1320 6700 1330 6740
rect 1370 6700 1380 6740
rect 1320 6680 1380 6700
rect 1430 6840 1490 6900
rect 1430 6800 1440 6840
rect 1480 6800 1490 6840
rect 1430 6740 1490 6800
rect 1430 6700 1440 6740
rect 1480 6700 1490 6740
rect 1430 6680 1490 6700
rect 1540 6840 1600 7020
rect 1640 6970 1720 6980
rect 1640 6910 1650 6970
rect 1710 6910 1720 6970
rect 1640 6900 1720 6910
rect 1540 6800 1550 6840
rect 1590 6800 1600 6840
rect 1540 6740 1600 6800
rect 1540 6700 1550 6740
rect 1590 6700 1600 6740
rect 1540 6680 1600 6700
rect 1650 6840 1710 6900
rect 1650 6800 1660 6840
rect 1700 6800 1710 6840
rect 1650 6740 1710 6800
rect 1650 6700 1660 6740
rect 1700 6700 1710 6740
rect 1650 6680 1710 6700
rect 1760 6840 1820 7020
rect 1860 6970 1940 6980
rect 1860 6910 1870 6970
rect 1930 6910 1940 6970
rect 1860 6900 1940 6910
rect 1760 6800 1770 6840
rect 1810 6800 1820 6840
rect 1760 6740 1820 6800
rect 1760 6700 1770 6740
rect 1810 6700 1820 6740
rect 1760 6680 1820 6700
rect 1870 6860 1930 6900
rect 1870 6840 2010 6860
rect 1870 6800 1880 6840
rect 1920 6800 1960 6840
rect 2000 6800 2010 6840
rect 1870 6740 2010 6800
rect 1870 6700 1880 6740
rect 1920 6700 1960 6740
rect 2000 6700 2010 6740
rect 1870 6680 2010 6700
rect -1184 6632 -1126 6640
rect -1184 6580 -1182 6632
rect -1130 6580 -1126 6632
rect -1184 6570 -1126 6580
rect -1074 6632 -1016 6640
rect -1074 6580 -1072 6632
rect -1020 6580 -1016 6632
rect -1074 6570 -1016 6580
rect -964 6632 -906 6640
rect -964 6580 -962 6632
rect -910 6580 -906 6632
rect -964 6570 -906 6580
rect -854 6632 -796 6640
rect -854 6580 -852 6632
rect -800 6580 -796 6632
rect -854 6570 -796 6580
rect -744 6632 -686 6640
rect -744 6580 -742 6632
rect -690 6580 -686 6632
rect -744 6570 -686 6580
rect -634 6632 -576 6640
rect -634 6580 -632 6632
rect -580 6580 -576 6632
rect -634 6570 -576 6580
rect -524 6632 -466 6640
rect -524 6580 -522 6632
rect -470 6580 -466 6632
rect -524 6570 -466 6580
rect -414 6632 -356 6640
rect -414 6580 -412 6632
rect -360 6580 -356 6632
rect -414 6570 -356 6580
rect -304 6632 -246 6640
rect -304 6580 -302 6632
rect -250 6580 -246 6632
rect -304 6570 -246 6580
rect -194 6632 -136 6640
rect -194 6580 -192 6632
rect -140 6580 -136 6632
rect -194 6570 -136 6580
rect 716 6632 774 6640
rect 716 6580 718 6632
rect 770 6580 774 6632
rect 716 6570 774 6580
rect 826 6632 884 6640
rect 826 6580 828 6632
rect 880 6580 884 6632
rect 826 6570 884 6580
rect 936 6632 994 6640
rect 936 6580 938 6632
rect 990 6580 994 6632
rect 936 6570 994 6580
rect 1046 6632 1104 6640
rect 1046 6580 1048 6632
rect 1100 6580 1104 6632
rect 1046 6570 1104 6580
rect 1156 6632 1214 6640
rect 1156 6580 1158 6632
rect 1210 6580 1214 6632
rect 1156 6570 1214 6580
rect 1266 6632 1324 6640
rect 1266 6580 1268 6632
rect 1320 6580 1324 6632
rect 1266 6570 1324 6580
rect 1376 6632 1434 6640
rect 1376 6580 1378 6632
rect 1430 6580 1434 6632
rect 1376 6570 1434 6580
rect 1486 6632 1544 6640
rect 1486 6580 1488 6632
rect 1540 6580 1544 6632
rect 1486 6570 1544 6580
rect 1596 6632 1654 6640
rect 1596 6580 1598 6632
rect 1650 6580 1654 6632
rect 1596 6570 1654 6580
rect 1706 6632 1764 6640
rect 1706 6580 1708 6632
rect 1760 6580 1764 6632
rect 1706 6570 1764 6580
rect -1370 6530 -1290 6540
rect -1370 6470 -1360 6530
rect -1300 6470 -1290 6530
rect -1370 6450 -1290 6470
rect -1370 6390 -1360 6450
rect -1300 6390 -1290 6450
rect -1370 6370 -1290 6390
rect -1370 6310 -1360 6370
rect -1300 6310 -1290 6370
rect -1370 6300 -1290 6310
rect -1010 6530 -930 6540
rect -1010 6470 -1000 6530
rect -940 6470 -930 6530
rect -1010 6450 -930 6470
rect -1010 6390 -1000 6450
rect -940 6390 -930 6450
rect -1010 6370 -930 6390
rect -1010 6310 -1000 6370
rect -940 6310 -930 6370
rect -1010 6300 -930 6310
rect -650 6530 -570 6540
rect -650 6470 -640 6530
rect -580 6470 -570 6530
rect -650 6450 -570 6470
rect -650 6390 -640 6450
rect -580 6390 -570 6450
rect -650 6370 -570 6390
rect -650 6310 -640 6370
rect -580 6310 -570 6370
rect -650 6300 -570 6310
rect -290 6530 -210 6540
rect -290 6470 -280 6530
rect -220 6470 -210 6530
rect -290 6450 -210 6470
rect -290 6390 -280 6450
rect -220 6390 -210 6450
rect -290 6370 -210 6390
rect -290 6310 -280 6370
rect -220 6310 -210 6370
rect -290 6300 -210 6310
rect 70 6530 150 6540
rect 70 6470 80 6530
rect 140 6470 150 6530
rect 70 6450 150 6470
rect 70 6390 80 6450
rect 140 6390 150 6450
rect 70 6370 150 6390
rect 70 6310 80 6370
rect 140 6310 150 6370
rect 70 6300 150 6310
rect 430 6530 510 6540
rect 430 6470 440 6530
rect 500 6470 510 6530
rect 430 6450 510 6470
rect 430 6390 440 6450
rect 500 6390 510 6450
rect 430 6370 510 6390
rect 430 6310 440 6370
rect 500 6310 510 6370
rect 430 6300 510 6310
rect 790 6530 870 6540
rect 790 6470 800 6530
rect 860 6470 870 6530
rect 790 6450 870 6470
rect 790 6390 800 6450
rect 860 6390 870 6450
rect 790 6370 870 6390
rect 790 6310 800 6370
rect 860 6310 870 6370
rect 790 6300 870 6310
rect 1150 6530 1230 6540
rect 1150 6470 1160 6530
rect 1220 6470 1230 6530
rect 1150 6450 1230 6470
rect 1150 6390 1160 6450
rect 1220 6390 1230 6450
rect 1150 6370 1230 6390
rect 1150 6310 1160 6370
rect 1220 6310 1230 6370
rect 1150 6300 1230 6310
rect 1510 6530 1590 6540
rect 1510 6470 1520 6530
rect 1580 6470 1590 6530
rect 1510 6450 1590 6470
rect 1510 6390 1520 6450
rect 1580 6390 1590 6450
rect 1510 6370 1590 6390
rect 1510 6310 1520 6370
rect 1580 6310 1590 6370
rect 1510 6300 1590 6310
rect 1870 6530 1950 6540
rect 1870 6470 1880 6530
rect 1940 6470 1950 6530
rect 1870 6450 1950 6470
rect 1870 6390 1880 6450
rect 1940 6390 1950 6450
rect 1870 6370 1950 6390
rect 1870 6310 1880 6370
rect 1940 6310 1950 6370
rect 1870 6300 1950 6310
rect 2500 6530 2580 6540
rect 2500 6470 2510 6530
rect 2570 6470 2580 6530
rect 2500 6450 2580 6470
rect 2500 6390 2510 6450
rect 2570 6390 2580 6450
rect 2500 6370 2580 6390
rect 2500 6310 2510 6370
rect 2570 6310 2580 6370
rect 2500 6300 2580 6310
rect 2940 6530 3020 6540
rect 2940 6470 2950 6530
rect 3010 6470 3020 6530
rect 2940 6450 3020 6470
rect 2940 6390 2950 6450
rect 3010 6390 3020 6450
rect 2940 6370 3020 6390
rect 2940 6310 2950 6370
rect 3010 6310 3020 6370
rect 2940 6300 3020 6310
rect -1360 6240 -1300 6260
rect -1360 6200 -1350 6240
rect -1310 6200 -1300 6240
rect -1360 6140 -1300 6200
rect -1360 6100 -1350 6140
rect -1310 6100 -1300 6140
rect -1360 6040 -1300 6100
rect -1360 6000 -1350 6040
rect -1310 6000 -1300 6040
rect -1360 5940 -1300 6000
rect -1360 5900 -1350 5940
rect -1310 5900 -1300 5940
rect -1360 5840 -1300 5900
rect -1360 5800 -1350 5840
rect -1310 5800 -1300 5840
rect -1360 5740 -1300 5800
rect -1360 5700 -1350 5740
rect -1310 5700 -1300 5740
rect -1360 5680 -1300 5700
rect -1180 6240 -1120 6260
rect -1180 6200 -1170 6240
rect -1130 6200 -1120 6240
rect -1180 6140 -1120 6200
rect -1180 6100 -1170 6140
rect -1130 6100 -1120 6140
rect -1180 6040 -1120 6100
rect -1180 6000 -1170 6040
rect -1130 6000 -1120 6040
rect -1180 5940 -1120 6000
rect -1180 5900 -1170 5940
rect -1130 5900 -1120 5940
rect -1180 5840 -1120 5900
rect -1180 5800 -1170 5840
rect -1130 5800 -1120 5840
rect -1180 5740 -1120 5800
rect -1180 5700 -1170 5740
rect -1130 5700 -1120 5740
rect -1180 5200 -1120 5700
rect -1000 6240 -940 6260
rect -1000 6200 -990 6240
rect -950 6200 -940 6240
rect -1000 6140 -940 6200
rect -1000 6100 -990 6140
rect -950 6100 -940 6140
rect -1000 6040 -940 6100
rect -1000 6000 -990 6040
rect -950 6000 -940 6040
rect -1000 5940 -940 6000
rect -1000 5900 -990 5940
rect -950 5900 -940 5940
rect -1000 5840 -940 5900
rect -1000 5800 -990 5840
rect -950 5800 -940 5840
rect -1000 5740 -940 5800
rect -1000 5700 -990 5740
rect -950 5700 -940 5740
rect -1000 5680 -940 5700
rect -820 6240 -760 6260
rect -820 6200 -810 6240
rect -770 6200 -760 6240
rect -820 6140 -760 6200
rect -820 6100 -810 6140
rect -770 6100 -760 6140
rect -820 6040 -760 6100
rect -820 6000 -810 6040
rect -770 6000 -760 6040
rect -820 5940 -760 6000
rect -820 5900 -810 5940
rect -770 5900 -760 5940
rect -820 5840 -760 5900
rect -820 5800 -810 5840
rect -770 5800 -760 5840
rect -820 5740 -760 5800
rect -820 5700 -810 5740
rect -770 5700 -760 5740
rect -820 5680 -760 5700
rect -640 6240 -580 6260
rect -640 6200 -630 6240
rect -590 6200 -580 6240
rect -640 6140 -580 6200
rect -640 6100 -630 6140
rect -590 6100 -580 6140
rect -640 6040 -580 6100
rect -640 6000 -630 6040
rect -590 6000 -580 6040
rect -640 5940 -580 6000
rect -640 5900 -630 5940
rect -590 5900 -580 5940
rect -640 5840 -580 5900
rect -640 5800 -630 5840
rect -590 5800 -580 5840
rect -640 5740 -580 5800
rect -640 5700 -630 5740
rect -590 5700 -580 5740
rect -640 5680 -580 5700
rect -460 6240 -400 6260
rect -460 6200 -450 6240
rect -410 6200 -400 6240
rect -460 6140 -400 6200
rect -460 6100 -450 6140
rect -410 6100 -400 6140
rect -460 6040 -400 6100
rect -460 6000 -450 6040
rect -410 6000 -400 6040
rect -460 5940 -400 6000
rect -460 5900 -450 5940
rect -410 5900 -400 5940
rect -460 5840 -400 5900
rect -460 5800 -450 5840
rect -410 5800 -400 5840
rect -460 5740 -400 5800
rect -460 5700 -450 5740
rect -410 5700 -400 5740
rect -460 5680 -400 5700
rect -280 6240 -220 6260
rect -280 6200 -270 6240
rect -230 6200 -220 6240
rect -280 6140 -220 6200
rect -280 6100 -270 6140
rect -230 6100 -220 6140
rect -280 6040 -220 6100
rect -280 6000 -270 6040
rect -230 6000 -220 6040
rect -280 5940 -220 6000
rect -280 5900 -270 5940
rect -230 5900 -220 5940
rect -280 5840 -220 5900
rect -280 5800 -270 5840
rect -230 5800 -220 5840
rect -280 5740 -220 5800
rect -280 5700 -270 5740
rect -230 5700 -220 5740
rect -280 5680 -220 5700
rect -100 6240 -40 6260
rect -100 6200 -90 6240
rect -50 6200 -40 6240
rect -100 6140 -40 6200
rect -100 6100 -90 6140
rect -50 6100 -40 6140
rect -100 6040 -40 6100
rect -100 6000 -90 6040
rect -50 6000 -40 6040
rect -100 5940 -40 6000
rect -100 5900 -90 5940
rect -50 5900 -40 5940
rect -100 5840 -40 5900
rect -100 5800 -90 5840
rect -50 5800 -40 5840
rect -100 5740 -40 5800
rect -100 5700 -90 5740
rect -50 5700 -40 5740
rect -100 5680 -40 5700
rect 80 6240 140 6260
rect 80 6200 90 6240
rect 130 6200 140 6240
rect 80 6140 140 6200
rect 80 6100 90 6140
rect 130 6100 140 6140
rect 80 6040 140 6100
rect 80 6000 90 6040
rect 130 6000 140 6040
rect 80 5940 140 6000
rect 80 5900 90 5940
rect 130 5900 140 5940
rect 80 5840 140 5900
rect 80 5800 90 5840
rect 130 5800 140 5840
rect 80 5740 140 5800
rect 80 5700 90 5740
rect 130 5700 140 5740
rect 80 5680 140 5700
rect 260 6240 320 6260
rect 260 6200 270 6240
rect 310 6200 320 6240
rect 260 6140 320 6200
rect 260 6100 270 6140
rect 310 6100 320 6140
rect 260 6040 320 6100
rect 260 6000 270 6040
rect 310 6000 320 6040
rect 260 5940 320 6000
rect 260 5900 270 5940
rect 310 5900 320 5940
rect 260 5840 320 5900
rect 260 5800 270 5840
rect 310 5800 320 5840
rect 260 5740 320 5800
rect 260 5700 270 5740
rect 310 5700 320 5740
rect -1090 5630 -1020 5640
rect -1030 5570 -1020 5630
rect -1090 5560 -1020 5570
rect -920 5630 -840 5640
rect -920 5570 -910 5630
rect -850 5570 -840 5630
rect -920 5560 -840 5570
rect -810 5310 -770 5680
rect -740 5630 -660 5640
rect -740 5570 -730 5630
rect -670 5570 -660 5630
rect -740 5560 -660 5570
rect -560 5630 -480 5640
rect -560 5570 -550 5630
rect -490 5570 -480 5630
rect -560 5560 -480 5570
rect -450 5420 -410 5680
rect -380 5630 -300 5640
rect -380 5570 -370 5630
rect -310 5570 -300 5630
rect -380 5560 -300 5570
rect -200 5630 -120 5640
rect -200 5570 -190 5630
rect -130 5570 -120 5630
rect -200 5560 -120 5570
rect -90 5530 -50 5680
rect -20 5630 60 5640
rect -20 5570 -10 5630
rect 50 5570 60 5630
rect -20 5560 60 5570
rect 160 5630 230 5640
rect 160 5570 170 5630
rect 160 5560 230 5570
rect -110 5520 -30 5530
rect -110 5460 -100 5520
rect -40 5460 -30 5520
rect -110 5450 -30 5460
rect -470 5410 -390 5420
rect -470 5350 -460 5410
rect -400 5350 -390 5410
rect -470 5340 -390 5350
rect -830 5300 -750 5310
rect -830 5240 -820 5300
rect -760 5240 -750 5300
rect -830 5230 -750 5240
rect 260 5200 320 5700
rect 440 6240 500 6260
rect 440 6200 450 6240
rect 490 6200 500 6240
rect 440 6140 500 6200
rect 440 6100 450 6140
rect 490 6100 500 6140
rect 440 6040 500 6100
rect 440 6000 450 6040
rect 490 6000 500 6040
rect 440 5940 500 6000
rect 440 5900 450 5940
rect 490 5900 500 5940
rect 440 5840 500 5900
rect 440 5800 450 5840
rect 490 5800 500 5840
rect 440 5740 500 5800
rect 440 5700 450 5740
rect 490 5700 500 5740
rect 440 5680 500 5700
rect 620 6240 680 6260
rect 620 6200 630 6240
rect 670 6200 680 6240
rect 620 6140 680 6200
rect 620 6100 630 6140
rect 670 6100 680 6140
rect 620 6040 680 6100
rect 620 6000 630 6040
rect 670 6000 680 6040
rect 620 5940 680 6000
rect 620 5900 630 5940
rect 670 5900 680 5940
rect 620 5840 680 5900
rect 620 5800 630 5840
rect 670 5800 680 5840
rect 620 5740 680 5800
rect 620 5700 630 5740
rect 670 5700 680 5740
rect 620 5680 680 5700
rect 800 6240 860 6260
rect 800 6200 810 6240
rect 850 6200 860 6240
rect 800 6140 860 6200
rect 800 6100 810 6140
rect 850 6100 860 6140
rect 800 6040 860 6100
rect 800 6000 810 6040
rect 850 6000 860 6040
rect 800 5940 860 6000
rect 800 5900 810 5940
rect 850 5900 860 5940
rect 800 5840 860 5900
rect 800 5800 810 5840
rect 850 5800 860 5840
rect 800 5740 860 5800
rect 800 5700 810 5740
rect 850 5700 860 5740
rect 800 5680 860 5700
rect 980 6240 1040 6260
rect 980 6200 990 6240
rect 1030 6200 1040 6240
rect 980 6140 1040 6200
rect 980 6100 990 6140
rect 1030 6100 1040 6140
rect 980 6040 1040 6100
rect 980 6000 990 6040
rect 1030 6000 1040 6040
rect 980 5940 1040 6000
rect 980 5900 990 5940
rect 1030 5900 1040 5940
rect 980 5840 1040 5900
rect 980 5800 990 5840
rect 1030 5800 1040 5840
rect 980 5740 1040 5800
rect 980 5700 990 5740
rect 1030 5700 1040 5740
rect 980 5680 1040 5700
rect 1160 6240 1220 6260
rect 1160 6200 1170 6240
rect 1210 6200 1220 6240
rect 1160 6140 1220 6200
rect 1160 6100 1170 6140
rect 1210 6100 1220 6140
rect 1160 6040 1220 6100
rect 1160 6000 1170 6040
rect 1210 6000 1220 6040
rect 1160 5940 1220 6000
rect 1160 5900 1170 5940
rect 1210 5900 1220 5940
rect 1160 5840 1220 5900
rect 1160 5800 1170 5840
rect 1210 5800 1220 5840
rect 1160 5740 1220 5800
rect 1160 5700 1170 5740
rect 1210 5700 1220 5740
rect 1160 5680 1220 5700
rect 1340 6240 1400 6260
rect 1340 6200 1350 6240
rect 1390 6200 1400 6240
rect 1340 6140 1400 6200
rect 1340 6100 1350 6140
rect 1390 6100 1400 6140
rect 1340 6040 1400 6100
rect 1340 6000 1350 6040
rect 1390 6000 1400 6040
rect 1340 5940 1400 6000
rect 1340 5900 1350 5940
rect 1390 5900 1400 5940
rect 1340 5840 1400 5900
rect 1340 5800 1350 5840
rect 1390 5800 1400 5840
rect 1340 5740 1400 5800
rect 1340 5700 1350 5740
rect 1390 5700 1400 5740
rect 1340 5680 1400 5700
rect 1520 6240 1580 6260
rect 1520 6200 1530 6240
rect 1570 6200 1580 6240
rect 1520 6140 1580 6200
rect 1520 6100 1530 6140
rect 1570 6100 1580 6140
rect 1520 6040 1580 6100
rect 1520 6000 1530 6040
rect 1570 6000 1580 6040
rect 1520 5940 1580 6000
rect 1520 5900 1530 5940
rect 1570 5900 1580 5940
rect 1520 5840 1580 5900
rect 1520 5800 1530 5840
rect 1570 5800 1580 5840
rect 1520 5740 1580 5800
rect 1520 5700 1530 5740
rect 1570 5700 1580 5740
rect 1520 5680 1580 5700
rect 1700 6240 1760 6260
rect 1700 6200 1710 6240
rect 1750 6200 1760 6240
rect 1700 6140 1760 6200
rect 1700 6100 1710 6140
rect 1750 6100 1760 6140
rect 1700 6040 1760 6100
rect 1700 6000 1710 6040
rect 1750 6000 1760 6040
rect 1700 5940 1760 6000
rect 1700 5900 1710 5940
rect 1750 5900 1760 5940
rect 1700 5840 1760 5900
rect 1700 5800 1710 5840
rect 1750 5800 1760 5840
rect 1700 5740 1760 5800
rect 1700 5700 1710 5740
rect 1750 5700 1760 5740
rect 350 5630 600 5640
rect 410 5570 440 5630
rect 500 5570 530 5630
rect 590 5570 600 5630
rect 350 5560 600 5570
rect -1190 5190 -1110 5200
rect -1190 5130 -1180 5190
rect -1120 5130 -1110 5190
rect -1190 5120 -1110 5130
rect 250 5190 330 5200
rect 250 5130 260 5190
rect 320 5130 330 5190
rect 250 5120 330 5130
rect -2470 5080 -2390 5090
rect -2470 5020 -2460 5080
rect -2400 5020 -2390 5080
rect -2470 5000 -2390 5020
rect -2470 4940 -2460 5000
rect -2400 4940 -2390 5000
rect -2470 4920 -2390 4940
rect -2470 4860 -2460 4920
rect -2400 4860 -2390 4920
rect -2470 4850 -2390 4860
rect -2230 5080 -2150 5090
rect -2230 5020 -2220 5080
rect -2160 5020 -2150 5080
rect -2230 5000 -2150 5020
rect -2230 4940 -2220 5000
rect -2160 4940 -2150 5000
rect -2230 4920 -2150 4940
rect -2230 4860 -2220 4920
rect -2160 4860 -2150 4920
rect -2230 4850 -2150 4860
rect -1990 5080 -1910 5090
rect -1990 5020 -1980 5080
rect -1920 5020 -1910 5080
rect -1990 5000 -1910 5020
rect -1990 4940 -1980 5000
rect -1920 4940 -1910 5000
rect -1990 4920 -1910 4940
rect -1990 4860 -1980 4920
rect -1920 4860 -1910 4920
rect -1990 4850 -1910 4860
rect -1750 5080 -1670 5090
rect -1750 5020 -1740 5080
rect -1680 5020 -1670 5080
rect -1750 5000 -1670 5020
rect -1750 4940 -1740 5000
rect -1680 4940 -1670 5000
rect -1750 4920 -1670 4940
rect -1750 4860 -1740 4920
rect -1680 4860 -1670 4920
rect -1750 4850 -1670 4860
rect -1510 5080 -1430 5090
rect -1510 5020 -1500 5080
rect -1440 5020 -1430 5080
rect -1510 5000 -1430 5020
rect -1510 4940 -1500 5000
rect -1440 4940 -1430 5000
rect -1510 4920 -1430 4940
rect -1510 4860 -1500 4920
rect -1440 4860 -1430 4920
rect -1510 4850 -1430 4860
rect -1270 5080 -1190 5090
rect -1270 5020 -1260 5080
rect -1200 5020 -1190 5080
rect -1270 5000 -1190 5020
rect -1270 4940 -1260 5000
rect -1200 4940 -1190 5000
rect -1270 4920 -1190 4940
rect -1270 4860 -1260 4920
rect -1200 4860 -1190 4920
rect -1270 4850 -1190 4860
rect -1030 5080 -950 5090
rect -1030 5020 -1020 5080
rect -960 5020 -950 5080
rect -1030 5000 -950 5020
rect -1030 4940 -1020 5000
rect -960 4940 -950 5000
rect -1030 4920 -950 4940
rect -1030 4860 -1020 4920
rect -960 4860 -950 4920
rect -1030 4850 -950 4860
rect -790 5080 -710 5090
rect -790 5020 -780 5080
rect -720 5020 -710 5080
rect -790 5000 -710 5020
rect -790 4940 -780 5000
rect -720 4940 -710 5000
rect -790 4920 -710 4940
rect -790 4860 -780 4920
rect -720 4860 -710 4920
rect -790 4850 -710 4860
rect -550 5080 -470 5090
rect -550 5020 -540 5080
rect -480 5020 -470 5080
rect -550 5000 -470 5020
rect -550 4940 -540 5000
rect -480 4940 -470 5000
rect -550 4920 -470 4940
rect -550 4860 -540 4920
rect -480 4860 -470 4920
rect -550 4850 -470 4860
rect -310 5080 -230 5090
rect -310 5020 -300 5080
rect -240 5020 -230 5080
rect -310 5000 -230 5020
rect -310 4940 -300 5000
rect -240 4940 -230 5000
rect -310 4920 -230 4940
rect -310 4860 -300 4920
rect -240 4860 -230 4920
rect -310 4850 -230 4860
rect -70 5080 10 5090
rect -70 5020 -60 5080
rect 0 5020 10 5080
rect -70 5000 10 5020
rect -70 4940 -60 5000
rect 0 4940 10 5000
rect -70 4920 10 4940
rect -70 4860 -60 4920
rect 0 4860 10 4920
rect -70 4850 10 4860
rect -2460 4800 -2400 4850
rect -2460 4760 -2450 4800
rect -2410 4760 -2400 4800
rect -2460 4680 -2400 4760
rect -2350 4810 -2270 4820
rect -2350 4750 -2340 4810
rect -2280 4750 -2270 4810
rect -2350 4740 -2270 4750
rect -2460 4640 -2450 4680
rect -2410 4640 -2400 4680
rect -2460 4580 -2400 4640
rect -2460 4540 -2450 4580
rect -2410 4540 -2400 4580
rect -2460 4520 -2400 4540
rect -2340 4680 -2280 4740
rect -2340 4640 -2330 4680
rect -2290 4640 -2280 4680
rect -2340 4580 -2280 4640
rect -2340 4540 -2330 4580
rect -2290 4540 -2280 4580
rect -2340 4520 -2280 4540
rect -2220 4680 -2160 4850
rect -2220 4640 -2210 4680
rect -2170 4640 -2160 4680
rect -2220 4580 -2160 4640
rect -2220 4540 -2210 4580
rect -2170 4540 -2160 4580
rect -2220 4520 -2160 4540
rect -2100 4680 -2040 4700
rect -2100 4640 -2090 4680
rect -2050 4640 -2040 4680
rect -2100 4580 -2040 4640
rect -2100 4540 -2090 4580
rect -2050 4540 -2040 4580
rect -2100 4480 -2040 4540
rect -1980 4680 -1920 4850
rect -1980 4640 -1970 4680
rect -1930 4640 -1920 4680
rect -1980 4580 -1920 4640
rect -1980 4540 -1970 4580
rect -1930 4540 -1920 4580
rect -1980 4520 -1920 4540
rect -1860 4680 -1800 4700
rect -1860 4640 -1850 4680
rect -1810 4640 -1800 4680
rect -1860 4580 -1800 4640
rect -1860 4540 -1850 4580
rect -1810 4540 -1800 4580
rect -2110 4470 -2030 4480
rect -2280 4450 -2220 4470
rect -2280 4410 -2270 4450
rect -2230 4410 -2220 4450
rect -2280 4360 -2220 4410
rect -2110 4410 -2100 4470
rect -2040 4410 -2030 4470
rect -2110 4400 -2030 4410
rect -1860 4360 -1800 4540
rect -1740 4680 -1680 4850
rect -1630 4810 -1550 4820
rect -1630 4750 -1620 4810
rect -1560 4750 -1550 4810
rect -1630 4740 -1550 4750
rect -1740 4640 -1730 4680
rect -1690 4640 -1680 4680
rect -1740 4580 -1680 4640
rect -1740 4540 -1730 4580
rect -1690 4540 -1680 4580
rect -1740 4520 -1680 4540
rect -1620 4680 -1560 4740
rect -1620 4640 -1610 4680
rect -1570 4640 -1560 4680
rect -1620 4580 -1560 4640
rect -1620 4540 -1610 4580
rect -1570 4540 -1560 4580
rect -1620 4520 -1560 4540
rect -1500 4680 -1440 4850
rect -1500 4640 -1490 4680
rect -1450 4640 -1440 4680
rect -1500 4580 -1440 4640
rect -1500 4540 -1490 4580
rect -1450 4540 -1440 4580
rect -1500 4520 -1440 4540
rect -1380 4680 -1320 4700
rect -1380 4640 -1370 4680
rect -1330 4640 -1320 4680
rect -1380 4580 -1320 4640
rect -1380 4540 -1370 4580
rect -1330 4540 -1320 4580
rect -1380 4480 -1320 4540
rect -1260 4680 -1200 4850
rect -1260 4640 -1250 4680
rect -1210 4640 -1200 4680
rect -1260 4580 -1200 4640
rect -1260 4540 -1250 4580
rect -1210 4540 -1200 4580
rect -1260 4520 -1200 4540
rect -1140 4680 -1080 4700
rect -1140 4640 -1130 4680
rect -1090 4640 -1080 4680
rect -1140 4580 -1080 4640
rect -1140 4540 -1130 4580
rect -1090 4540 -1080 4580
rect -1620 4460 -1560 4480
rect -1620 4420 -1610 4460
rect -1570 4420 -1560 4460
rect -1620 4360 -1560 4420
rect -1390 4470 -1310 4480
rect -1390 4410 -1380 4470
rect -1320 4410 -1310 4470
rect -2640 3580 -2630 3640
rect -2570 3580 -2560 3640
rect -2640 1900 -2560 3580
rect -2370 4350 -2210 4360
rect -2370 4290 -2360 4350
rect -2300 4290 -2280 4350
rect -2220 4290 -2210 4350
rect -2370 4280 -2210 4290
rect -1870 4350 -1790 4360
rect -1870 4290 -1860 4350
rect -1800 4290 -1790 4350
rect -1870 4280 -1790 4290
rect -1630 4350 -1550 4360
rect -1630 4290 -1620 4350
rect -1560 4290 -1550 4350
rect -2370 2010 -2290 4280
rect -1630 4080 -1550 4290
rect -1630 4020 -1620 4080
rect -1560 4020 -1550 4080
rect -1630 4010 -1550 4020
rect -1620 3740 -1560 4010
rect -1390 3970 -1310 4410
rect -1140 4360 -1080 4540
rect -1020 4680 -960 4850
rect -910 4810 -830 4820
rect -910 4750 -900 4810
rect -840 4750 -830 4810
rect -910 4740 -830 4750
rect -1020 4640 -1010 4680
rect -970 4640 -960 4680
rect -1020 4580 -960 4640
rect -1020 4540 -1010 4580
rect -970 4540 -960 4580
rect -1020 4520 -960 4540
rect -900 4680 -840 4740
rect -900 4640 -890 4680
rect -850 4640 -840 4680
rect -900 4580 -840 4640
rect -900 4540 -890 4580
rect -850 4540 -840 4580
rect -900 4520 -840 4540
rect -780 4680 -720 4850
rect -780 4640 -770 4680
rect -730 4640 -720 4680
rect -780 4580 -720 4640
rect -780 4540 -770 4580
rect -730 4540 -720 4580
rect -780 4520 -720 4540
rect -660 4680 -600 4700
rect -660 4640 -650 4680
rect -610 4640 -600 4680
rect -660 4580 -600 4640
rect -660 4540 -650 4580
rect -610 4540 -600 4580
rect -660 4480 -600 4540
rect -540 4680 -480 4850
rect -540 4640 -530 4680
rect -490 4640 -480 4680
rect -540 4580 -480 4640
rect -540 4540 -530 4580
rect -490 4540 -480 4580
rect -540 4520 -480 4540
rect -420 4680 -360 4700
rect -420 4640 -410 4680
rect -370 4640 -360 4680
rect -420 4580 -360 4640
rect -420 4540 -410 4580
rect -370 4540 -360 4580
rect -900 4460 -840 4480
rect -900 4420 -890 4460
rect -850 4420 -840 4460
rect -900 4360 -840 4420
rect -670 4470 -590 4480
rect -670 4410 -660 4470
rect -600 4410 -590 4470
rect -670 4400 -590 4410
rect -420 4360 -360 4540
rect -300 4680 -240 4850
rect -190 4810 -110 4820
rect -190 4750 -180 4810
rect -120 4750 -110 4810
rect -190 4740 -110 4750
rect -60 4800 0 4850
rect -60 4760 -50 4800
rect -10 4760 0 4800
rect -300 4640 -290 4680
rect -250 4640 -240 4680
rect -300 4580 -240 4640
rect -300 4540 -290 4580
rect -250 4540 -240 4580
rect -300 4520 -240 4540
rect -180 4680 -120 4740
rect -180 4640 -170 4680
rect -130 4640 -120 4680
rect -180 4580 -120 4640
rect -180 4540 -170 4580
rect -130 4540 -120 4580
rect -180 4520 -120 4540
rect -60 4680 0 4760
rect 70 4810 150 4820
rect 70 4750 80 4810
rect 140 4750 150 4810
rect 70 4740 150 4750
rect 430 4810 510 5560
rect 630 5530 670 5680
rect 700 5630 780 5640
rect 700 5570 710 5630
rect 770 5570 780 5630
rect 700 5560 780 5570
rect 880 5630 960 5640
rect 880 5570 890 5630
rect 950 5570 960 5630
rect 880 5560 960 5570
rect 610 5520 690 5530
rect 610 5460 620 5520
rect 680 5460 690 5520
rect 610 5450 690 5460
rect 990 5420 1030 5680
rect 1060 5630 1140 5640
rect 1060 5570 1070 5630
rect 1130 5570 1140 5630
rect 1060 5560 1140 5570
rect 1240 5630 1320 5640
rect 1240 5570 1250 5630
rect 1310 5570 1320 5630
rect 1240 5560 1320 5570
rect 970 5410 1050 5420
rect 970 5350 980 5410
rect 1040 5350 1050 5410
rect 970 5340 1050 5350
rect 1350 5310 1390 5680
rect 1420 5630 1500 5640
rect 1420 5570 1430 5630
rect 1490 5570 1500 5630
rect 1420 5560 1500 5570
rect 1600 5630 1670 5640
rect 1600 5570 1610 5630
rect 1600 5560 1670 5570
rect 1330 5300 1410 5310
rect 1330 5240 1340 5300
rect 1400 5240 1410 5300
rect 1330 5230 1410 5240
rect 1700 5200 1760 5700
rect 1880 6240 1940 6260
rect 1880 6200 1890 6240
rect 1930 6200 1940 6240
rect 1880 6140 1940 6200
rect 2510 6180 2570 6300
rect 2950 6180 3010 6300
rect 1880 6100 1890 6140
rect 1930 6100 1940 6140
rect 2250 6170 2330 6180
rect 2250 6110 2260 6170
rect 2320 6110 2330 6170
rect 2250 6100 2330 6110
rect 2500 6160 2580 6180
rect 2500 6120 2520 6160
rect 2560 6120 2580 6160
rect 2500 6100 2580 6120
rect 2720 6170 2800 6180
rect 2720 6110 2730 6170
rect 2790 6110 2800 6170
rect 2720 6100 2800 6110
rect 2940 6160 3020 6180
rect 2940 6120 2960 6160
rect 3000 6120 3020 6160
rect 2940 6100 3020 6120
rect 1880 6040 1940 6100
rect 1880 6000 1890 6040
rect 1930 6000 1940 6040
rect 1880 5940 1940 6000
rect 1880 5900 1890 5940
rect 1930 5900 1940 5940
rect 1880 5840 1940 5900
rect 1880 5800 1890 5840
rect 1930 5800 1940 5840
rect 1880 5740 1940 5800
rect 1880 5700 1890 5740
rect 1930 5700 1940 5740
rect 1880 5680 1940 5700
rect 2270 5420 2310 6100
rect 2510 6040 2570 6100
rect 2510 6000 2520 6040
rect 2560 6000 2570 6040
rect 2510 5940 2570 6000
rect 2510 5900 2520 5940
rect 2560 5900 2570 5940
rect 2510 5880 2570 5900
rect 2620 6040 2680 6060
rect 2620 6000 2630 6040
rect 2670 6000 2680 6040
rect 2620 5940 2680 6000
rect 2620 5900 2630 5940
rect 2670 5900 2680 5940
rect 2620 5840 2680 5900
rect 2730 6040 2790 6100
rect 2730 6000 2740 6040
rect 2780 6000 2790 6040
rect 2730 5940 2790 6000
rect 2730 5900 2740 5940
rect 2780 5900 2790 5940
rect 2730 5880 2790 5900
rect 2840 6040 2900 6060
rect 2840 6000 2850 6040
rect 2890 6000 2900 6040
rect 2840 5940 2900 6000
rect 2840 5900 2850 5940
rect 2890 5900 2900 5940
rect 2840 5840 2900 5900
rect 2950 6040 3010 6100
rect 2950 6000 2960 6040
rect 3000 6000 3010 6040
rect 2950 5940 3010 6000
rect 2950 5900 2960 5940
rect 3000 5900 3010 5940
rect 2950 5880 3010 5900
rect 2600 5830 2680 5840
rect 2600 5770 2610 5830
rect 2670 5770 2680 5830
rect 2600 5760 2680 5770
rect 2720 5820 2800 5840
rect 2720 5780 2740 5820
rect 2780 5780 2800 5820
rect 2250 5410 2330 5420
rect 2250 5350 2260 5410
rect 2320 5350 2330 5410
rect 2250 5340 2330 5350
rect 2720 5300 2800 5780
rect 2840 5830 2920 5840
rect 2840 5770 2850 5830
rect 2910 5770 2920 5830
rect 2840 5760 2920 5770
rect 2720 5240 2730 5300
rect 2790 5240 2800 5300
rect 2720 5230 2800 5240
rect 1690 5190 1770 5200
rect 1690 5130 1700 5190
rect 1760 5130 1770 5190
rect 1690 5120 1770 5130
rect 570 5080 650 5090
rect 570 5020 580 5080
rect 640 5020 650 5080
rect 570 5000 650 5020
rect 570 4940 580 5000
rect 640 4940 650 5000
rect 570 4920 650 4940
rect 570 4860 580 4920
rect 640 4860 650 4920
rect 570 4850 650 4860
rect 810 5080 890 5090
rect 810 5020 820 5080
rect 880 5020 890 5080
rect 810 5000 890 5020
rect 810 4940 820 5000
rect 880 4940 890 5000
rect 810 4920 890 4940
rect 810 4860 820 4920
rect 880 4860 890 4920
rect 810 4850 890 4860
rect 1050 5080 1130 5090
rect 1050 5020 1060 5080
rect 1120 5020 1130 5080
rect 1050 5000 1130 5020
rect 1050 4940 1060 5000
rect 1120 4940 1130 5000
rect 1050 4920 1130 4940
rect 1050 4860 1060 4920
rect 1120 4860 1130 4920
rect 1050 4850 1130 4860
rect 1290 5080 1370 5090
rect 1290 5020 1300 5080
rect 1360 5020 1370 5080
rect 1290 5000 1370 5020
rect 1290 4940 1300 5000
rect 1360 4940 1370 5000
rect 1290 4920 1370 4940
rect 1290 4860 1300 4920
rect 1360 4860 1370 4920
rect 1290 4850 1370 4860
rect 1530 5080 1610 5090
rect 1530 5020 1540 5080
rect 1600 5020 1610 5080
rect 1530 5000 1610 5020
rect 1530 4940 1540 5000
rect 1600 4940 1610 5000
rect 1530 4920 1610 4940
rect 1530 4860 1540 4920
rect 1600 4860 1610 4920
rect 1530 4850 1610 4860
rect 1770 5080 1850 5090
rect 1770 5020 1780 5080
rect 1840 5020 1850 5080
rect 1770 5000 1850 5020
rect 1770 4940 1780 5000
rect 1840 4940 1850 5000
rect 1770 4920 1850 4940
rect 1770 4860 1780 4920
rect 1840 4860 1850 4920
rect 1770 4850 1850 4860
rect 2010 5080 2090 5090
rect 2010 5020 2020 5080
rect 2080 5020 2090 5080
rect 2010 5000 2090 5020
rect 2010 4940 2020 5000
rect 2080 4940 2090 5000
rect 2010 4920 2090 4940
rect 2010 4860 2020 4920
rect 2080 4860 2090 4920
rect 2010 4850 2090 4860
rect 2250 5080 2330 5090
rect 2250 5020 2260 5080
rect 2320 5020 2330 5080
rect 2250 5000 2330 5020
rect 2250 4940 2260 5000
rect 2320 4940 2330 5000
rect 2250 4920 2330 4940
rect 2250 4860 2260 4920
rect 2320 4860 2330 4920
rect 2250 4850 2330 4860
rect 2490 5080 2570 5090
rect 2490 5020 2500 5080
rect 2560 5020 2570 5080
rect 2490 5000 2570 5020
rect 2490 4940 2500 5000
rect 2560 4940 2570 5000
rect 2490 4920 2570 4940
rect 2490 4860 2500 4920
rect 2560 4860 2570 4920
rect 2490 4850 2570 4860
rect 2730 5080 2810 5090
rect 2730 5020 2740 5080
rect 2800 5020 2810 5080
rect 2730 5000 2810 5020
rect 2730 4940 2740 5000
rect 2800 4940 2810 5000
rect 2730 4920 2810 4940
rect 2730 4860 2740 4920
rect 2800 4860 2810 4920
rect 2730 4850 2810 4860
rect 430 4750 440 4810
rect 500 4750 510 4810
rect 430 4740 510 4750
rect 580 4800 640 4850
rect 580 4760 590 4800
rect 630 4760 640 4800
rect -60 4640 -50 4680
rect -10 4640 0 4680
rect -60 4580 0 4640
rect -60 4540 -50 4580
rect -10 4540 0 4580
rect -60 4520 0 4540
rect -240 4460 -180 4480
rect -240 4420 -230 4460
rect -190 4420 -180 4460
rect -240 4360 -180 4420
rect -1150 4350 -1070 4360
rect -1150 4290 -1140 4350
rect -1080 4290 -1070 4350
rect -1150 4280 -1070 4290
rect -910 4350 -830 4360
rect -910 4290 -900 4350
rect -840 4290 -830 4350
rect -910 4280 -830 4290
rect -430 4350 -350 4360
rect -430 4290 -420 4350
rect -360 4290 -350 4350
rect -430 4280 -350 4290
rect -250 4350 -170 4360
rect -250 4290 -240 4350
rect -180 4290 -170 4350
rect -250 4280 -170 4290
rect -1150 4080 -1070 4090
rect -1150 4020 -1140 4080
rect -1080 4020 -1070 4080
rect -1150 4010 -1070 4020
rect -670 4080 -590 4090
rect -670 4020 -660 4080
rect -600 4020 -590 4080
rect -670 4010 -590 4020
rect -1390 3910 -1380 3970
rect -1320 3910 -1310 3970
rect -1390 3900 -1310 3910
rect -1458 3860 -1400 3870
rect -1458 3808 -1454 3860
rect -1402 3808 -1400 3860
rect -1458 3800 -1400 3808
rect -1370 3760 -1330 3900
rect -1300 3860 -1242 3870
rect -1300 3808 -1296 3860
rect -1244 3808 -1242 3860
rect -1300 3800 -1242 3808
rect -1130 3760 -1090 4010
rect -910 3970 -830 3980
rect -910 3910 -900 3970
rect -840 3910 -830 3970
rect -910 3900 -830 3910
rect -976 3860 -918 3870
rect -976 3808 -972 3860
rect -920 3808 -918 3860
rect -976 3800 -918 3808
rect -890 3760 -850 3900
rect -822 3860 -764 3870
rect -822 3808 -818 3860
rect -766 3808 -764 3860
rect -822 3800 -764 3808
rect -650 3760 -610 4010
rect -430 3970 -350 3980
rect -430 3910 -420 3970
rect -360 3910 -350 3970
rect -430 3900 -350 3910
rect -498 3860 -440 3870
rect -498 3808 -494 3860
rect -442 3808 -440 3860
rect -498 3800 -440 3808
rect -410 3760 -370 3900
rect -190 3820 -110 3830
rect -190 3760 -180 3820
rect -120 3760 -110 3820
rect -1620 3700 -1610 3740
rect -1570 3700 -1560 3740
rect -1620 3680 -1560 3700
rect -1500 3740 -1440 3760
rect -1500 3700 -1490 3740
rect -1450 3700 -1440 3740
rect -1500 3680 -1440 3700
rect -1380 3740 -1320 3760
rect -1380 3700 -1370 3740
rect -1330 3700 -1320 3740
rect -1380 3680 -1320 3700
rect -1260 3740 -1200 3760
rect -1260 3700 -1250 3740
rect -1210 3700 -1200 3740
rect -1260 3680 -1200 3700
rect -1140 3740 -1080 3760
rect -1140 3700 -1130 3740
rect -1090 3700 -1080 3740
rect -1140 3680 -1080 3700
rect -1020 3740 -960 3760
rect -1020 3700 -1010 3740
rect -970 3700 -960 3740
rect -1020 3680 -960 3700
rect -900 3740 -840 3760
rect -900 3700 -890 3740
rect -850 3700 -840 3740
rect -900 3680 -840 3700
rect -780 3740 -720 3760
rect -780 3700 -770 3740
rect -730 3700 -720 3740
rect -780 3680 -720 3700
rect -660 3740 -600 3760
rect -660 3700 -650 3740
rect -610 3700 -600 3740
rect -660 3680 -600 3700
rect -540 3740 -480 3760
rect -540 3700 -530 3740
rect -490 3700 -480 3740
rect -540 3680 -480 3700
rect -420 3740 -360 3760
rect -420 3700 -410 3740
rect -370 3700 -360 3740
rect -420 3680 -360 3700
rect -190 3740 -110 3760
rect -190 3680 -180 3740
rect -120 3680 -110 3740
rect -1559 3632 -1501 3640
rect -1559 3580 -1557 3632
rect -1505 3580 -1501 3632
rect -1559 3570 -1501 3580
rect -1470 3540 -1440 3680
rect -1260 3540 -1230 3680
rect -1199 3632 -1141 3640
rect -1199 3580 -1197 3632
rect -1145 3580 -1141 3632
rect -1199 3570 -1141 3580
rect -1079 3632 -1021 3640
rect -1079 3580 -1077 3632
rect -1025 3580 -1021 3632
rect -1079 3570 -1021 3580
rect -990 3540 -960 3680
rect -780 3540 -750 3680
rect -719 3632 -661 3640
rect -719 3580 -717 3632
rect -665 3580 -661 3632
rect -719 3570 -661 3580
rect -599 3632 -541 3640
rect -599 3580 -597 3632
rect -545 3580 -541 3632
rect -599 3570 -541 3580
rect -510 3540 -480 3680
rect -190 3660 -110 3680
rect -190 3600 -180 3660
rect -120 3600 -110 3660
rect -190 3590 -110 3600
rect -2250 3530 -2170 3540
rect -2250 3470 -2240 3530
rect -2180 3470 -2170 3530
rect -2250 3460 -2170 3470
rect -1500 3530 -1420 3540
rect -1500 3470 -1490 3530
rect -1430 3470 -1420 3530
rect -1500 3460 -1420 3470
rect -1280 3530 -1200 3540
rect -1280 3470 -1270 3530
rect -1210 3470 -1200 3530
rect -1280 3460 -1200 3470
rect -1020 3530 -940 3540
rect -1020 3470 -1010 3530
rect -950 3470 -940 3530
rect -1020 3460 -940 3470
rect -800 3530 -720 3540
rect -800 3470 -790 3530
rect -730 3470 -720 3530
rect -800 3460 -720 3470
rect -540 3530 -460 3540
rect -540 3470 -530 3530
rect -470 3470 -460 3530
rect -540 3460 -460 3470
rect -2230 3230 -2190 3460
rect -2070 3420 -1990 3430
rect -2070 3360 -2060 3420
rect -2000 3360 -1990 3420
rect -2070 3340 -1990 3360
rect -2070 3280 -2060 3340
rect -2000 3280 -1990 3340
rect -2070 3260 -1990 3280
rect -2250 3210 -2170 3230
rect -2250 3170 -2230 3210
rect -2190 3170 -2170 3210
rect -2070 3200 -2060 3260
rect -2000 3200 -1990 3260
rect -2070 3190 -1990 3200
rect -1830 3420 -1750 3430
rect -1830 3360 -1820 3420
rect -1760 3360 -1750 3420
rect -1830 3340 -1750 3360
rect -1830 3280 -1820 3340
rect -1760 3280 -1750 3340
rect -1830 3260 -1750 3280
rect -1830 3200 -1820 3260
rect -1760 3200 -1750 3260
rect -1830 3190 -1750 3200
rect -1590 3420 -1510 3430
rect -1590 3360 -1580 3420
rect -1520 3360 -1510 3420
rect -1590 3340 -1510 3360
rect -1590 3280 -1580 3340
rect -1520 3280 -1510 3340
rect -1590 3260 -1510 3280
rect -1590 3200 -1580 3260
rect -1520 3200 -1510 3260
rect -1590 3190 -1510 3200
rect -1350 3420 -1270 3430
rect -1350 3360 -1340 3420
rect -1280 3360 -1270 3420
rect -1350 3340 -1270 3360
rect -1350 3280 -1340 3340
rect -1280 3280 -1270 3340
rect -1350 3260 -1270 3280
rect -1350 3200 -1340 3260
rect -1280 3200 -1270 3260
rect -1350 3190 -1270 3200
rect -710 3420 -630 3430
rect -710 3360 -700 3420
rect -640 3360 -630 3420
rect -710 3340 -630 3360
rect -710 3280 -700 3340
rect -640 3280 -630 3340
rect -710 3260 -630 3280
rect -710 3200 -700 3260
rect -640 3200 -630 3260
rect -710 3190 -630 3200
rect -470 3420 -390 3430
rect -470 3360 -460 3420
rect -400 3360 -390 3420
rect -470 3340 -390 3360
rect -470 3280 -460 3340
rect -400 3280 -390 3340
rect -470 3260 -390 3280
rect -470 3200 -460 3260
rect -400 3200 -390 3260
rect -470 3190 -390 3200
rect -230 3420 -150 3430
rect -230 3360 -220 3420
rect -160 3360 -150 3420
rect -230 3340 -150 3360
rect -230 3280 -220 3340
rect -160 3280 -150 3340
rect -230 3260 -150 3280
rect -230 3200 -220 3260
rect -160 3200 -150 3260
rect -230 3190 -150 3200
rect 80 3220 140 4740
rect -2250 3150 -2170 3170
rect 80 3180 90 3220
rect 130 3180 140 3220
rect 80 3160 140 3180
rect 170 3820 410 3830
rect 170 3760 180 3820
rect 240 3760 260 3820
rect 320 3760 340 3820
rect 400 3760 410 3820
rect 170 3740 410 3760
rect 170 3680 180 3740
rect 240 3680 260 3740
rect 320 3680 340 3740
rect 400 3680 410 3740
rect 170 3660 410 3680
rect 170 3600 180 3660
rect 240 3600 260 3660
rect 320 3600 340 3660
rect 400 3600 410 3660
rect -1090 2620 -1010 2630
rect -1090 2560 -1080 2620
rect -1020 2560 -1010 2620
rect -1090 2540 -1010 2560
rect -1090 2480 -1080 2540
rect -1020 2480 -1010 2540
rect -1090 2460 -1010 2480
rect -1090 2400 -1080 2460
rect -1020 2400 -1010 2460
rect -1090 2390 -1010 2400
rect 170 2620 410 3600
rect 440 3220 500 4740
rect 580 4680 640 4760
rect 690 4810 770 4820
rect 690 4750 700 4810
rect 760 4750 770 4810
rect 690 4740 770 4750
rect 580 4640 590 4680
rect 630 4640 640 4680
rect 580 4580 640 4640
rect 580 4540 590 4580
rect 630 4540 640 4580
rect 580 4520 640 4540
rect 700 4680 760 4740
rect 700 4640 710 4680
rect 750 4640 760 4680
rect 700 4580 760 4640
rect 700 4540 710 4580
rect 750 4540 760 4580
rect 700 4520 760 4540
rect 820 4680 880 4850
rect 820 4640 830 4680
rect 870 4640 880 4680
rect 820 4580 880 4640
rect 820 4540 830 4580
rect 870 4540 880 4580
rect 820 4520 880 4540
rect 940 4680 1000 4700
rect 940 4640 950 4680
rect 990 4640 1000 4680
rect 940 4580 1000 4640
rect 940 4540 950 4580
rect 990 4540 1000 4580
rect 760 4460 820 4480
rect 760 4420 770 4460
rect 810 4420 820 4460
rect 760 4360 820 4420
rect 940 4360 1000 4540
rect 1060 4680 1120 4850
rect 1060 4640 1070 4680
rect 1110 4640 1120 4680
rect 1060 4580 1120 4640
rect 1060 4540 1070 4580
rect 1110 4540 1120 4580
rect 1060 4520 1120 4540
rect 1180 4680 1240 4700
rect 1180 4640 1190 4680
rect 1230 4640 1240 4680
rect 1180 4580 1240 4640
rect 1180 4540 1190 4580
rect 1230 4540 1240 4580
rect 1180 4480 1240 4540
rect 1300 4680 1360 4850
rect 1410 4810 1490 4820
rect 1410 4750 1420 4810
rect 1480 4750 1490 4810
rect 1410 4740 1490 4750
rect 1300 4640 1310 4680
rect 1350 4640 1360 4680
rect 1300 4580 1360 4640
rect 1300 4540 1310 4580
rect 1350 4540 1360 4580
rect 1300 4520 1360 4540
rect 1420 4680 1480 4740
rect 1420 4640 1430 4680
rect 1470 4640 1480 4680
rect 1420 4580 1480 4640
rect 1420 4540 1430 4580
rect 1470 4540 1480 4580
rect 1420 4520 1480 4540
rect 1540 4680 1600 4850
rect 1540 4640 1550 4680
rect 1590 4640 1600 4680
rect 1540 4580 1600 4640
rect 1540 4540 1550 4580
rect 1590 4540 1600 4580
rect 1540 4520 1600 4540
rect 1660 4680 1720 4700
rect 1660 4640 1670 4680
rect 1710 4640 1720 4680
rect 1660 4580 1720 4640
rect 1660 4540 1670 4580
rect 1710 4540 1720 4580
rect 1170 4470 1250 4480
rect 1170 4410 1180 4470
rect 1240 4410 1250 4470
rect 1170 4400 1250 4410
rect 1420 4460 1480 4480
rect 1420 4420 1430 4460
rect 1470 4420 1480 4460
rect 1420 4360 1480 4420
rect 1660 4360 1720 4540
rect 1780 4680 1840 4850
rect 1780 4640 1790 4680
rect 1830 4640 1840 4680
rect 1780 4580 1840 4640
rect 1780 4540 1790 4580
rect 1830 4540 1840 4580
rect 1780 4520 1840 4540
rect 1900 4680 1960 4700
rect 1900 4640 1910 4680
rect 1950 4640 1960 4680
rect 1900 4580 1960 4640
rect 1900 4540 1910 4580
rect 1950 4540 1960 4580
rect 1900 4480 1960 4540
rect 2020 4680 2080 4850
rect 2130 4810 2210 4820
rect 2130 4750 2140 4810
rect 2200 4750 2210 4810
rect 2130 4740 2210 4750
rect 2020 4640 2030 4680
rect 2070 4640 2080 4680
rect 2020 4580 2080 4640
rect 2020 4540 2030 4580
rect 2070 4540 2080 4580
rect 2020 4520 2080 4540
rect 2140 4680 2200 4740
rect 2140 4640 2150 4680
rect 2190 4640 2200 4680
rect 2140 4580 2200 4640
rect 2140 4540 2150 4580
rect 2190 4540 2200 4580
rect 2140 4520 2200 4540
rect 2260 4680 2320 4850
rect 2260 4640 2270 4680
rect 2310 4640 2320 4680
rect 2260 4580 2320 4640
rect 2260 4540 2270 4580
rect 2310 4540 2320 4580
rect 2260 4520 2320 4540
rect 2380 4680 2440 4700
rect 2380 4640 2390 4680
rect 2430 4640 2440 4680
rect 2380 4580 2440 4640
rect 2380 4540 2390 4580
rect 2430 4540 2440 4580
rect 1890 4470 1970 4480
rect 1890 4410 1900 4470
rect 1960 4410 1970 4470
rect 750 4350 830 4360
rect 750 4290 760 4350
rect 820 4290 830 4350
rect 750 4270 830 4290
rect 750 4210 760 4270
rect 820 4210 830 4270
rect 750 4190 830 4210
rect 750 4130 760 4190
rect 820 4130 830 4190
rect 750 4120 830 4130
rect 930 4350 1010 4360
rect 930 4290 940 4350
rect 1000 4290 1010 4350
rect 930 4270 1010 4290
rect 930 4210 940 4270
rect 1000 4210 1010 4270
rect 930 4190 1010 4210
rect 930 4130 940 4190
rect 1000 4130 1010 4190
rect 930 4120 1010 4130
rect 1170 4350 1250 4360
rect 1170 4290 1180 4350
rect 1240 4290 1250 4350
rect 1170 4270 1250 4290
rect 1170 4210 1180 4270
rect 1240 4210 1250 4270
rect 1170 4190 1250 4210
rect 1170 4130 1180 4190
rect 1240 4130 1250 4190
rect 1170 4120 1250 4130
rect 1410 4350 1490 4360
rect 1410 4290 1420 4350
rect 1480 4290 1490 4350
rect 1410 4270 1490 4290
rect 1410 4210 1420 4270
rect 1480 4210 1490 4270
rect 1410 4190 1490 4210
rect 1410 4130 1420 4190
rect 1480 4130 1490 4190
rect 1410 4120 1490 4130
rect 1650 4350 1730 4360
rect 1650 4290 1660 4350
rect 1720 4290 1730 4350
rect 1650 4270 1730 4290
rect 1650 4210 1660 4270
rect 1720 4210 1730 4270
rect 1650 4190 1730 4210
rect 1650 4130 1660 4190
rect 1720 4130 1730 4190
rect 1650 4120 1730 4130
rect 1170 4080 1250 4090
rect 1170 4020 1180 4080
rect 1240 4020 1250 4080
rect 1170 4010 1250 4020
rect 1650 4080 1730 4090
rect 1650 4020 1660 4080
rect 1720 4020 1730 4080
rect 1650 4010 1730 4020
rect 930 3970 1010 3980
rect 930 3910 940 3970
rect 1000 3910 1010 3970
rect 930 3900 1010 3910
rect 690 3820 770 3830
rect 690 3760 700 3820
rect 760 3760 770 3820
rect 950 3760 990 3900
rect 1020 3860 1078 3870
rect 1020 3808 1022 3860
rect 1074 3808 1078 3860
rect 1020 3800 1078 3808
rect 1190 3760 1230 4010
rect 1410 3970 1490 3980
rect 1410 3910 1420 3970
rect 1480 3910 1490 3970
rect 1410 3900 1490 3910
rect 1344 3860 1402 3870
rect 1344 3808 1346 3860
rect 1398 3808 1402 3860
rect 1344 3800 1402 3808
rect 1430 3760 1470 3900
rect 1498 3860 1556 3870
rect 1498 3808 1500 3860
rect 1552 3808 1556 3860
rect 1498 3800 1556 3808
rect 1670 3760 1710 4010
rect 1890 3970 1970 4410
rect 2140 4460 2200 4480
rect 2140 4420 2150 4460
rect 2190 4420 2200 4460
rect 2140 4360 2200 4420
rect 2380 4360 2440 4540
rect 2500 4680 2560 4850
rect 2500 4640 2510 4680
rect 2550 4640 2560 4680
rect 2500 4580 2560 4640
rect 2500 4540 2510 4580
rect 2550 4540 2560 4580
rect 2500 4520 2560 4540
rect 2620 4680 2680 4700
rect 2620 4640 2630 4680
rect 2670 4640 2680 4680
rect 2620 4580 2680 4640
rect 2620 4540 2630 4580
rect 2670 4540 2680 4580
rect 2620 4480 2680 4540
rect 2740 4680 2800 4850
rect 2850 4810 2930 5760
rect 3160 5520 3240 5530
rect 3160 5460 3170 5520
rect 3230 5460 3240 5520
rect 3160 5450 3240 5460
rect 2970 5080 3050 5090
rect 2970 5020 2980 5080
rect 3040 5020 3050 5080
rect 2970 5000 3050 5020
rect 2970 4940 2980 5000
rect 3040 4940 3050 5000
rect 2970 4920 3050 4940
rect 2970 4860 2980 4920
rect 3040 4860 3050 4920
rect 2970 4850 3050 4860
rect 2850 4750 2860 4810
rect 2920 4750 2930 4810
rect 2850 4740 2930 4750
rect 2980 4800 3040 4850
rect 2980 4760 2990 4800
rect 3030 4760 3040 4800
rect 2740 4640 2750 4680
rect 2790 4640 2800 4680
rect 2740 4580 2800 4640
rect 2740 4540 2750 4580
rect 2790 4540 2800 4580
rect 2740 4520 2800 4540
rect 2860 4680 2920 4740
rect 2860 4640 2870 4680
rect 2910 4640 2920 4680
rect 2860 4580 2920 4640
rect 2860 4540 2870 4580
rect 2910 4540 2920 4580
rect 2860 4520 2920 4540
rect 2980 4680 3040 4760
rect 2980 4640 2990 4680
rect 3030 4640 3040 4680
rect 2980 4580 3040 4640
rect 2980 4540 2990 4580
rect 3030 4540 3040 4580
rect 2980 4520 3040 4540
rect 2610 4470 2690 4480
rect 2610 4410 2620 4470
rect 2680 4410 2690 4470
rect 2610 4400 2690 4410
rect 2800 4450 2860 4470
rect 2800 4410 2810 4450
rect 2850 4410 2860 4450
rect 2800 4360 2860 4410
rect 2130 4350 2210 4360
rect 2130 4290 2140 4350
rect 2200 4290 2210 4350
rect 2130 4270 2210 4290
rect 2130 4210 2140 4270
rect 2200 4210 2210 4270
rect 2130 4190 2210 4210
rect 2130 4130 2140 4190
rect 2200 4130 2210 4190
rect 2130 4080 2210 4130
rect 2370 4350 2450 4360
rect 2370 4290 2380 4350
rect 2440 4290 2450 4350
rect 2370 4270 2450 4290
rect 2370 4210 2380 4270
rect 2440 4210 2450 4270
rect 2370 4190 2450 4210
rect 2370 4130 2380 4190
rect 2440 4130 2450 4190
rect 2370 4120 2450 4130
rect 2790 4350 2870 4360
rect 2790 4290 2800 4350
rect 2860 4290 2870 4350
rect 2790 4270 2870 4290
rect 2790 4210 2800 4270
rect 2860 4210 2870 4270
rect 2790 4190 2870 4210
rect 2790 4130 2800 4190
rect 2860 4130 2870 4190
rect 2790 4120 2870 4130
rect 2130 4020 2140 4080
rect 2200 4020 2210 4080
rect 2130 4010 2210 4020
rect 1890 3910 1900 3970
rect 1960 3910 1970 3970
rect 1890 3900 1970 3910
rect 1822 3860 1880 3870
rect 1822 3808 1824 3860
rect 1876 3808 1880 3860
rect 1822 3800 1880 3808
rect 1910 3760 1950 3900
rect 1980 3860 2038 3870
rect 1980 3808 1982 3860
rect 2034 3808 2038 3860
rect 1980 3800 2038 3808
rect 690 3740 770 3760
rect 690 3680 700 3740
rect 760 3680 770 3740
rect 940 3740 1000 3760
rect 940 3700 950 3740
rect 990 3700 1000 3740
rect 940 3680 1000 3700
rect 1060 3740 1120 3760
rect 1060 3700 1070 3740
rect 1110 3700 1120 3740
rect 1060 3680 1120 3700
rect 1180 3740 1240 3760
rect 1180 3700 1190 3740
rect 1230 3700 1240 3740
rect 1180 3680 1240 3700
rect 1300 3740 1360 3760
rect 1300 3700 1310 3740
rect 1350 3700 1360 3740
rect 1300 3680 1360 3700
rect 1420 3740 1480 3760
rect 1420 3700 1430 3740
rect 1470 3700 1480 3740
rect 1420 3680 1480 3700
rect 1540 3740 1600 3760
rect 1540 3700 1550 3740
rect 1590 3700 1600 3740
rect 1540 3680 1600 3700
rect 1660 3740 1720 3760
rect 1660 3700 1670 3740
rect 1710 3700 1720 3740
rect 1660 3680 1720 3700
rect 1780 3740 1840 3760
rect 1780 3700 1790 3740
rect 1830 3700 1840 3740
rect 1780 3680 1840 3700
rect 1900 3740 1960 3760
rect 1900 3700 1910 3740
rect 1950 3700 1960 3740
rect 1900 3680 1960 3700
rect 2020 3740 2080 3760
rect 2020 3700 2030 3740
rect 2070 3700 2080 3740
rect 2020 3680 2080 3700
rect 2140 3740 2200 4010
rect 2140 3700 2150 3740
rect 2190 3700 2200 3740
rect 2140 3680 2200 3700
rect 690 3660 770 3680
rect 690 3600 700 3660
rect 760 3600 770 3660
rect 690 3590 770 3600
rect 1060 3540 1090 3680
rect 1121 3632 1179 3640
rect 1121 3580 1125 3632
rect 1177 3580 1179 3632
rect 1121 3570 1179 3580
rect 1241 3632 1299 3640
rect 1241 3580 1245 3632
rect 1297 3580 1299 3632
rect 1241 3570 1299 3580
rect 1330 3540 1360 3680
rect 1540 3540 1570 3680
rect 1601 3632 1659 3640
rect 1601 3580 1605 3632
rect 1657 3580 1659 3632
rect 1601 3570 1659 3580
rect 1721 3632 1779 3640
rect 1721 3580 1725 3632
rect 1777 3580 1779 3632
rect 1721 3570 1779 3580
rect 1810 3540 1840 3680
rect 2020 3540 2050 3680
rect 3180 3650 3220 5450
rect 3250 5410 3330 5420
rect 3250 5350 3260 5410
rect 3320 5350 3330 5410
rect 3250 5340 3330 5350
rect 3270 3880 3310 5340
rect 5030 5140 5110 9290
rect 6090 9350 6170 9420
rect 6310 9760 6390 9940
rect 6750 10000 6830 10010
rect 6750 9940 6760 10000
rect 6820 9940 6830 10000
rect 6310 9720 6330 9760
rect 6370 9720 6390 9760
rect 6310 9660 6390 9720
rect 6310 9620 6330 9660
rect 6370 9620 6390 9660
rect 6310 9560 6390 9620
rect 6310 9520 6330 9560
rect 6370 9520 6390 9560
rect 6310 9460 6390 9520
rect 6310 9420 6330 9460
rect 6370 9420 6390 9460
rect 6310 9400 6390 9420
rect 6530 9760 6610 9780
rect 6530 9720 6550 9760
rect 6590 9720 6610 9760
rect 6530 9660 6610 9720
rect 6530 9620 6550 9660
rect 6590 9620 6610 9660
rect 6530 9560 6610 9620
rect 6530 9520 6550 9560
rect 6590 9520 6610 9560
rect 6530 9460 6610 9520
rect 6530 9420 6550 9460
rect 6590 9420 6610 9460
rect 6090 9290 6100 9350
rect 6160 9290 6170 9350
rect 6090 9280 6170 9290
rect 6310 9340 6390 9360
rect 6310 9300 6330 9340
rect 6370 9300 6390 9340
rect 5250 9230 5330 9240
rect 5250 9170 5260 9230
rect 5320 9170 5330 9230
rect 5250 7890 5330 9170
rect 6310 9230 6390 9300
rect 6530 9350 6610 9420
rect 6750 9760 6830 9940
rect 7070 10000 7150 10010
rect 7070 9940 7080 10000
rect 7140 9940 7150 10000
rect 7070 9780 7150 9940
rect 7390 10000 7470 10010
rect 7390 9940 7400 10000
rect 7460 9940 7470 10000
rect 6750 9720 6770 9760
rect 6810 9720 6830 9760
rect 6750 9660 6830 9720
rect 6750 9620 6770 9660
rect 6810 9620 6830 9660
rect 6750 9560 6830 9620
rect 6750 9520 6770 9560
rect 6810 9520 6830 9560
rect 6750 9460 6830 9520
rect 6750 9420 6770 9460
rect 6810 9420 6830 9460
rect 6750 9400 6830 9420
rect 6970 9760 7250 9780
rect 6970 9720 6990 9760
rect 7030 9720 7090 9760
rect 7130 9720 7190 9760
rect 7230 9720 7250 9760
rect 6970 9660 7250 9720
rect 6970 9620 6990 9660
rect 7030 9620 7090 9660
rect 7130 9620 7190 9660
rect 7230 9620 7250 9660
rect 6970 9560 7250 9620
rect 6970 9520 6990 9560
rect 7030 9520 7090 9560
rect 7130 9520 7190 9560
rect 7230 9520 7250 9560
rect 6970 9460 7250 9520
rect 6970 9420 6990 9460
rect 7030 9420 7090 9460
rect 7130 9420 7190 9460
rect 7230 9420 7250 9460
rect 6970 9400 7250 9420
rect 7390 9760 7470 9940
rect 7830 10000 7910 10010
rect 7830 9940 7840 10000
rect 7900 9940 7910 10000
rect 7390 9720 7410 9760
rect 7450 9720 7470 9760
rect 7390 9660 7470 9720
rect 7390 9620 7410 9660
rect 7450 9620 7470 9660
rect 7390 9560 7470 9620
rect 7390 9520 7410 9560
rect 7450 9520 7470 9560
rect 7390 9460 7470 9520
rect 7390 9420 7410 9460
rect 7450 9420 7470 9460
rect 7390 9400 7470 9420
rect 7610 9760 7690 9780
rect 7610 9720 7630 9760
rect 7670 9720 7690 9760
rect 7610 9660 7690 9720
rect 7610 9620 7630 9660
rect 7670 9620 7690 9660
rect 7610 9560 7690 9620
rect 7610 9520 7630 9560
rect 7670 9520 7690 9560
rect 7610 9460 7690 9520
rect 7610 9420 7630 9460
rect 7670 9420 7690 9460
rect 6530 9290 6540 9350
rect 6600 9290 6610 9350
rect 6530 9280 6610 9290
rect 6970 9350 7050 9360
rect 6970 9290 6980 9350
rect 7040 9290 7050 9350
rect 7610 9350 7690 9420
rect 7830 9760 7910 9940
rect 8270 10000 8350 10010
rect 8270 9940 8280 10000
rect 8340 9940 8350 10000
rect 7830 9720 7850 9760
rect 7890 9720 7910 9760
rect 7830 9660 7910 9720
rect 7830 9620 7850 9660
rect 7890 9620 7910 9660
rect 7830 9560 7910 9620
rect 7830 9520 7850 9560
rect 7890 9520 7910 9560
rect 7830 9460 7910 9520
rect 7830 9420 7850 9460
rect 7890 9420 7910 9460
rect 7830 9400 7910 9420
rect 8050 9760 8130 9780
rect 8050 9720 8070 9760
rect 8110 9720 8130 9760
rect 8050 9660 8130 9720
rect 8050 9620 8070 9660
rect 8110 9620 8130 9660
rect 8050 9560 8130 9620
rect 8050 9520 8070 9560
rect 8110 9520 8130 9560
rect 8050 9460 8130 9520
rect 8050 9420 8070 9460
rect 8110 9420 8130 9460
rect 6310 9170 6320 9230
rect 6380 9170 6390 9230
rect 6310 9160 6390 9170
rect 5890 9010 5970 9020
rect 5890 8950 5900 9010
rect 5960 8950 5970 9010
rect 5890 8770 5970 8950
rect 5890 8730 5910 8770
rect 5950 8730 5970 8770
rect 5890 8710 5970 8730
rect 5450 8660 5530 8680
rect 5450 8620 5470 8660
rect 5510 8620 5530 8660
rect 5450 8560 5530 8620
rect 5450 8520 5470 8560
rect 5510 8520 5530 8560
rect 5450 8460 5530 8520
rect 5450 8420 5470 8460
rect 5510 8420 5530 8460
rect 5450 8360 5530 8420
rect 5450 8320 5470 8360
rect 5510 8320 5530 8360
rect 5450 8240 5530 8320
rect 5450 8200 5470 8240
rect 5510 8200 5530 8240
rect 5450 8160 5530 8200
rect 5450 8100 5460 8160
rect 5520 8100 5530 8160
rect 5450 8090 5530 8100
rect 5670 8660 5750 8680
rect 5670 8620 5690 8660
rect 5730 8620 5750 8660
rect 5670 8560 5750 8620
rect 5670 8520 5690 8560
rect 5730 8520 5750 8560
rect 5670 8460 5750 8520
rect 5670 8420 5690 8460
rect 5730 8420 5750 8460
rect 5670 8360 5750 8420
rect 5670 8320 5690 8360
rect 5730 8320 5750 8360
rect 5670 8160 5750 8320
rect 5890 8660 5970 8680
rect 5890 8620 5910 8660
rect 5950 8620 5970 8660
rect 5890 8560 5970 8620
rect 5890 8520 5910 8560
rect 5950 8520 5970 8560
rect 5890 8460 5970 8520
rect 5890 8420 5910 8460
rect 5950 8420 5970 8460
rect 5890 8360 5970 8420
rect 5890 8320 5910 8360
rect 5950 8320 5970 8360
rect 5890 8300 5970 8320
rect 6110 8660 6190 8680
rect 6110 8620 6130 8660
rect 6170 8620 6190 8660
rect 6110 8560 6190 8620
rect 6110 8520 6130 8560
rect 6170 8520 6190 8560
rect 6110 8460 6190 8520
rect 6110 8420 6130 8460
rect 6170 8420 6190 8460
rect 6110 8360 6190 8420
rect 6110 8320 6130 8360
rect 6170 8320 6190 8360
rect 5670 8100 5680 8160
rect 5740 8100 5750 8160
rect 5670 8090 5750 8100
rect 6110 8160 6190 8320
rect 6330 8660 6610 8680
rect 6330 8620 6350 8660
rect 6390 8620 6450 8660
rect 6490 8620 6550 8660
rect 6590 8620 6610 8660
rect 6330 8560 6610 8620
rect 6330 8520 6350 8560
rect 6390 8520 6450 8560
rect 6490 8520 6550 8560
rect 6590 8520 6610 8560
rect 6330 8460 6610 8520
rect 6330 8420 6350 8460
rect 6390 8420 6450 8460
rect 6490 8420 6550 8460
rect 6590 8420 6610 8460
rect 6330 8360 6610 8420
rect 6330 8320 6350 8360
rect 6390 8320 6450 8360
rect 6490 8320 6550 8360
rect 6590 8320 6610 8360
rect 6330 8300 6610 8320
rect 6750 8660 6830 8680
rect 6750 8620 6770 8660
rect 6810 8620 6830 8660
rect 6750 8560 6830 8620
rect 6750 8520 6770 8560
rect 6810 8520 6830 8560
rect 6750 8460 6830 8520
rect 6750 8420 6770 8460
rect 6810 8420 6830 8460
rect 6750 8360 6830 8420
rect 6750 8320 6770 8360
rect 6810 8320 6830 8360
rect 6110 8100 6120 8160
rect 6180 8100 6190 8160
rect 6110 8090 6190 8100
rect 6430 8160 6510 8300
rect 6430 8100 6440 8160
rect 6500 8100 6510 8160
rect 6430 8090 6510 8100
rect 6750 8160 6830 8320
rect 6970 8660 7050 9290
rect 7480 9320 7560 9330
rect 7480 9260 7490 9320
rect 7550 9260 7560 9320
rect 7610 9290 7620 9350
rect 7680 9290 7690 9350
rect 7610 9280 7690 9290
rect 8050 9350 8130 9420
rect 8270 9760 8350 9940
rect 8270 9720 8290 9760
rect 8330 9720 8350 9760
rect 8270 9660 8350 9720
rect 8270 9620 8290 9660
rect 8330 9620 8350 9660
rect 8270 9560 8350 9620
rect 8270 9520 8290 9560
rect 8330 9520 8350 9560
rect 8270 9460 8350 9520
rect 8270 9420 8290 9460
rect 8330 9420 8350 9460
rect 8270 9400 8350 9420
rect 8490 10000 8570 10010
rect 8490 9940 8500 10000
rect 8560 9940 8570 10000
rect 8490 9880 8570 9940
rect 8490 9840 8510 9880
rect 8550 9840 8570 9880
rect 8490 9760 8570 9840
rect 8490 9720 8510 9760
rect 8550 9720 8570 9760
rect 8490 9660 8570 9720
rect 8490 9620 8510 9660
rect 8550 9620 8570 9660
rect 8490 9560 8570 9620
rect 8490 9520 8510 9560
rect 8550 9520 8570 9560
rect 8490 9460 8570 9520
rect 8490 9420 8510 9460
rect 8550 9420 8570 9460
rect 8490 9400 8570 9420
rect 8050 9290 8060 9350
rect 8120 9290 8130 9350
rect 8850 9340 8960 9360
rect 7480 9120 7560 9260
rect 7480 9060 7490 9120
rect 7550 9060 7560 9120
rect 7480 9050 7560 9060
rect 8050 9070 8130 9290
rect 8180 9320 8260 9330
rect 8180 9260 8190 9320
rect 8250 9260 8260 9320
rect 8180 9250 8260 9260
rect 8850 9270 8870 9340
rect 8940 9270 8960 9340
rect 8850 9250 8960 9270
rect 8050 9010 8060 9070
rect 8120 9010 8130 9070
rect 7920 8820 8000 8830
rect 7920 8760 7930 8820
rect 7990 8760 8000 8820
rect 7920 8750 8000 8760
rect 6970 8620 6990 8660
rect 7030 8620 7050 8660
rect 6970 8560 7050 8620
rect 6970 8520 6990 8560
rect 7030 8520 7050 8560
rect 6970 8460 7050 8520
rect 6970 8420 6990 8460
rect 7030 8420 7050 8460
rect 6970 8360 7050 8420
rect 6970 8320 6990 8360
rect 7030 8320 7050 8360
rect 6970 8300 7050 8320
rect 7190 8660 7270 8680
rect 7190 8620 7210 8660
rect 7250 8620 7270 8660
rect 7190 8560 7270 8620
rect 7190 8520 7210 8560
rect 7250 8520 7270 8560
rect 7190 8460 7270 8520
rect 7190 8420 7210 8460
rect 7250 8420 7270 8460
rect 7190 8360 7270 8420
rect 7190 8320 7210 8360
rect 7250 8320 7270 8360
rect 6750 8100 6760 8160
rect 6820 8100 6830 8160
rect 6750 8090 6830 8100
rect 7190 8160 7270 8320
rect 7410 8660 7690 8680
rect 7410 8620 7430 8660
rect 7470 8620 7530 8660
rect 7570 8620 7630 8660
rect 7670 8620 7690 8660
rect 7410 8560 7690 8620
rect 7410 8520 7430 8560
rect 7470 8520 7530 8560
rect 7570 8520 7630 8560
rect 7670 8520 7690 8560
rect 7410 8460 7690 8520
rect 7410 8420 7430 8460
rect 7470 8420 7530 8460
rect 7570 8420 7630 8460
rect 7670 8420 7690 8460
rect 7410 8360 7690 8420
rect 7410 8320 7430 8360
rect 7470 8320 7530 8360
rect 7570 8320 7630 8360
rect 7670 8320 7690 8360
rect 7410 8300 7690 8320
rect 7830 8660 7910 8680
rect 7830 8620 7850 8660
rect 7890 8620 7910 8660
rect 7830 8560 7910 8620
rect 7830 8520 7850 8560
rect 7890 8520 7910 8560
rect 7830 8460 7910 8520
rect 7830 8420 7850 8460
rect 7890 8420 7910 8460
rect 7830 8360 7910 8420
rect 7830 8320 7850 8360
rect 7890 8320 7910 8360
rect 7190 8100 7200 8160
rect 7260 8100 7270 8160
rect 7190 8090 7270 8100
rect 7510 8160 7590 8300
rect 7510 8100 7520 8160
rect 7580 8100 7590 8160
rect 7510 8090 7590 8100
rect 7830 8160 7910 8320
rect 8050 8660 8130 9010
rect 12110 9070 12190 13490
rect 12110 9010 12120 9070
rect 12180 9010 12190 9070
rect 8180 8820 8260 8830
rect 8180 8760 8190 8820
rect 8250 8760 8260 8820
rect 8180 8750 8260 8760
rect 8850 8810 8960 8830
rect 8850 8740 8870 8810
rect 8940 8740 8960 8810
rect 8850 8720 8960 8740
rect 8050 8620 8070 8660
rect 8110 8620 8130 8660
rect 8050 8560 8130 8620
rect 8050 8520 8070 8560
rect 8110 8520 8130 8560
rect 8050 8460 8130 8520
rect 8050 8420 8070 8460
rect 8110 8420 8130 8460
rect 8050 8360 8130 8420
rect 8050 8320 8070 8360
rect 8110 8320 8130 8360
rect 8050 8300 8130 8320
rect 8270 8660 8350 8680
rect 8270 8620 8290 8660
rect 8330 8620 8350 8660
rect 8270 8560 8350 8620
rect 8270 8520 8290 8560
rect 8330 8520 8350 8560
rect 8270 8460 8350 8520
rect 8270 8420 8290 8460
rect 8330 8420 8350 8460
rect 8270 8360 8350 8420
rect 8270 8320 8290 8360
rect 8330 8320 8350 8360
rect 7830 8100 7840 8160
rect 7900 8100 7910 8160
rect 7830 8090 7910 8100
rect 8270 8160 8350 8320
rect 8270 8100 8280 8160
rect 8340 8100 8350 8160
rect 8270 8090 8350 8100
rect 8490 8660 8570 8680
rect 8490 8620 8510 8660
rect 8550 8620 8570 8660
rect 8490 8560 8570 8620
rect 8490 8520 8510 8560
rect 8550 8520 8570 8560
rect 8490 8460 8570 8520
rect 8490 8420 8510 8460
rect 8550 8420 8570 8460
rect 8490 8360 8570 8420
rect 8490 8320 8510 8360
rect 8550 8320 8570 8360
rect 8490 8240 8570 8320
rect 8490 8200 8510 8240
rect 8550 8200 8570 8240
rect 8490 8160 8570 8200
rect 8490 8100 8500 8160
rect 8560 8100 8570 8160
rect 8490 8090 8570 8100
rect 9200 8020 9310 8040
rect 9200 7950 9220 8020
rect 9290 7950 9310 8020
rect 9200 7930 9310 7950
rect 5250 7830 5260 7890
rect 5320 7830 5330 7890
rect 5250 7820 5330 7830
rect 12000 7890 12080 7900
rect 12000 7830 12010 7890
rect 12070 7830 12080 7890
rect 5030 5080 5040 5140
rect 5100 5080 5110 5140
rect 5030 5070 5110 5080
rect 5140 7780 5220 7790
rect 5140 7720 5150 7780
rect 5210 7720 5220 7780
rect 5140 7700 5220 7720
rect 5140 7640 5150 7700
rect 5210 7640 5220 7700
rect 5140 7620 5220 7640
rect 5140 7560 5150 7620
rect 5210 7560 5220 7620
rect 5140 4980 5220 7560
rect 9320 7260 9420 7280
rect 9320 7200 9340 7260
rect 9400 7200 9420 7260
rect 9320 7180 9420 7200
rect 9120 6740 9200 6750
rect 9120 6680 9130 6740
rect 9190 6680 9200 6740
rect 9120 6670 9200 6680
rect 5140 4920 5150 4980
rect 5210 4920 5220 4980
rect 5140 4910 5220 4920
rect 5250 6350 5330 6360
rect 5250 6290 5260 6350
rect 5320 6290 5330 6350
rect 3480 4810 3560 4820
rect 3480 4750 3490 4810
rect 3550 4750 3560 4810
rect 3250 3870 3330 3880
rect 3250 3810 3260 3870
rect 3320 3810 3330 3870
rect 3250 3800 3330 3810
rect 3160 3640 3240 3650
rect 2081 3632 2139 3640
rect 2081 3580 2085 3632
rect 2137 3580 2139 3632
rect 2081 3570 2139 3580
rect 3160 3580 3170 3640
rect 3230 3580 3240 3640
rect 3160 3570 3240 3580
rect 1040 3530 1120 3540
rect 1040 3470 1050 3530
rect 1110 3470 1120 3530
rect 1040 3460 1120 3470
rect 1300 3530 1380 3540
rect 1300 3470 1310 3530
rect 1370 3470 1380 3530
rect 1300 3460 1380 3470
rect 1520 3530 1600 3540
rect 1520 3470 1530 3530
rect 1590 3470 1600 3530
rect 1520 3460 1600 3470
rect 1780 3530 1860 3540
rect 1780 3470 1790 3530
rect 1850 3470 1860 3530
rect 1780 3460 1860 3470
rect 2000 3530 2080 3540
rect 2000 3470 2010 3530
rect 2070 3470 2080 3530
rect 2000 3460 2080 3470
rect 2750 3530 2830 3540
rect 2750 3470 2760 3530
rect 2820 3470 2830 3530
rect 2750 3460 2830 3470
rect 440 3180 450 3220
rect 490 3180 500 3220
rect 730 3420 810 3430
rect 730 3360 740 3420
rect 800 3360 810 3420
rect 730 3340 810 3360
rect 730 3280 740 3340
rect 800 3280 810 3340
rect 730 3260 810 3280
rect 730 3200 740 3260
rect 800 3200 810 3260
rect 730 3190 810 3200
rect 970 3420 1050 3430
rect 970 3360 980 3420
rect 1040 3360 1050 3420
rect 970 3340 1050 3360
rect 970 3280 980 3340
rect 1040 3280 1050 3340
rect 970 3260 1050 3280
rect 970 3200 980 3260
rect 1040 3200 1050 3260
rect 970 3190 1050 3200
rect 1210 3420 1290 3430
rect 1210 3360 1220 3420
rect 1280 3360 1290 3420
rect 1210 3340 1290 3360
rect 1210 3280 1220 3340
rect 1280 3280 1290 3340
rect 1210 3260 1290 3280
rect 1210 3200 1220 3260
rect 1280 3200 1290 3260
rect 1210 3190 1290 3200
rect 1850 3420 1930 3430
rect 1850 3360 1860 3420
rect 1920 3360 1930 3420
rect 1850 3340 1930 3360
rect 1850 3280 1860 3340
rect 1920 3280 1930 3340
rect 1850 3260 1930 3280
rect 1850 3200 1860 3260
rect 1920 3200 1930 3260
rect 1850 3190 1930 3200
rect 2090 3420 2170 3430
rect 2090 3360 2100 3420
rect 2160 3360 2170 3420
rect 2090 3340 2170 3360
rect 2090 3280 2100 3340
rect 2160 3280 2170 3340
rect 2090 3260 2170 3280
rect 2090 3200 2100 3260
rect 2160 3200 2170 3260
rect 2090 3190 2170 3200
rect 2330 3420 2410 3430
rect 2330 3360 2340 3420
rect 2400 3360 2410 3420
rect 2330 3340 2410 3360
rect 2330 3280 2340 3340
rect 2400 3280 2410 3340
rect 2330 3260 2410 3280
rect 2330 3200 2340 3260
rect 2400 3200 2410 3260
rect 2330 3190 2410 3200
rect 2570 3420 2650 3430
rect 2570 3360 2580 3420
rect 2640 3360 2650 3420
rect 2570 3340 2650 3360
rect 2570 3280 2580 3340
rect 2640 3280 2650 3340
rect 2570 3260 2650 3280
rect 2570 3200 2580 3260
rect 2640 3200 2650 3260
rect 2570 3190 2650 3200
rect 440 3160 500 3180
rect 2760 3130 2820 3460
rect 2760 3090 2770 3130
rect 2810 3090 2820 3130
rect 2760 3030 2820 3090
rect 2760 2990 2770 3030
rect 2810 2990 2820 3030
rect 2760 2930 2820 2990
rect 2760 2890 2770 2930
rect 2810 2890 2820 2930
rect 2760 2830 2820 2890
rect 2760 2790 2770 2830
rect 2810 2790 2820 2830
rect 2760 2730 2820 2790
rect 2760 2690 2770 2730
rect 2810 2690 2820 2730
rect 2760 2670 2820 2690
rect 170 2560 180 2620
rect 240 2560 260 2620
rect 320 2560 340 2620
rect 400 2560 410 2620
rect 170 2540 410 2560
rect 170 2480 180 2540
rect 240 2480 260 2540
rect 320 2480 340 2540
rect 400 2480 410 2540
rect 170 2460 410 2480
rect 170 2400 180 2460
rect 240 2400 260 2460
rect 320 2400 340 2460
rect 400 2400 410 2460
rect 170 2390 410 2400
rect 1590 2620 1670 2630
rect 1590 2560 1600 2620
rect 1660 2560 1670 2620
rect 1590 2540 1670 2560
rect 1590 2480 1600 2540
rect 1660 2480 1670 2540
rect 1590 2460 1670 2480
rect 1590 2400 1600 2460
rect 1660 2400 1670 2460
rect 1590 2390 1670 2400
rect -1830 2350 -1750 2360
rect -1830 2290 -1820 2350
rect -1760 2290 -1750 2350
rect -1830 2280 -1750 2290
rect -1670 2350 -1590 2360
rect -1670 2290 -1660 2350
rect -1600 2290 -1590 2350
rect -1670 2280 -1590 2290
rect -1510 2350 -1430 2360
rect -1510 2290 -1500 2350
rect -1440 2290 -1430 2350
rect -1510 2280 -1430 2290
rect -1350 2350 -1270 2360
rect -1350 2290 -1340 2350
rect -1280 2290 -1270 2350
rect -1350 2280 -1270 2290
rect -1190 2350 -1110 2360
rect -1190 2290 -1180 2350
rect -1120 2290 -1110 2350
rect -1190 2280 -1110 2290
rect -1030 2350 -950 2360
rect -1030 2290 -1020 2350
rect -960 2290 -950 2350
rect -1030 2280 -950 2290
rect -870 2350 -790 2360
rect -870 2290 -860 2350
rect -800 2290 -790 2350
rect -870 2280 -790 2290
rect -710 2350 -630 2360
rect -710 2290 -700 2350
rect -640 2290 -630 2350
rect -710 2280 -630 2290
rect -550 2350 -470 2360
rect -550 2290 -540 2350
rect -480 2290 -470 2350
rect -550 2280 -470 2290
rect -390 2350 -310 2360
rect -390 2290 -380 2350
rect -320 2290 -310 2350
rect -390 2280 -310 2290
rect -230 2350 -150 2360
rect -230 2290 -220 2350
rect -160 2290 -150 2350
rect -230 2280 -150 2290
rect -70 2350 10 2360
rect -70 2290 -60 2350
rect 0 2290 10 2350
rect -70 2280 10 2290
rect 90 2350 170 2360
rect 90 2290 100 2350
rect 160 2290 170 2350
rect 90 2280 170 2290
rect 250 2350 330 2360
rect 250 2290 260 2350
rect 320 2290 330 2350
rect 250 2280 330 2290
rect 410 2350 490 2360
rect 410 2290 420 2350
rect 480 2290 490 2350
rect 410 2280 490 2290
rect 570 2350 650 2360
rect 570 2290 580 2350
rect 640 2290 650 2350
rect 570 2280 650 2290
rect 730 2350 810 2360
rect 730 2290 740 2350
rect 800 2290 810 2350
rect 730 2280 810 2290
rect 890 2350 970 2360
rect 890 2290 900 2350
rect 960 2290 970 2350
rect 890 2280 970 2290
rect 1050 2350 1130 2360
rect 1050 2290 1060 2350
rect 1120 2290 1130 2350
rect 1050 2280 1130 2290
rect 1210 2350 1290 2360
rect 1210 2290 1220 2350
rect 1280 2290 1290 2350
rect 1210 2280 1290 2290
rect 1370 2350 1450 2360
rect 1370 2290 1380 2350
rect 1440 2290 1450 2350
rect 1370 2280 1450 2290
rect 1530 2350 1610 2360
rect 1530 2290 1540 2350
rect 1600 2290 1610 2350
rect 1530 2280 1610 2290
rect 1690 2350 1770 2360
rect 1690 2290 1700 2350
rect 1760 2290 1770 2350
rect 1690 2280 1770 2290
rect 1850 2350 1930 2360
rect 1850 2290 1860 2350
rect 1920 2290 1930 2350
rect 1850 2280 1930 2290
rect 2010 2350 2090 2360
rect 2010 2290 2020 2350
rect 2080 2290 2090 2350
rect 2010 2280 2090 2290
rect 2170 2350 2250 2360
rect 2170 2290 2180 2350
rect 2240 2290 2250 2350
rect 2170 2280 2250 2290
rect 2480 2220 2560 2230
rect -1910 2180 -1830 2190
rect -1910 2120 -1900 2180
rect -1840 2120 -1830 2180
rect -1910 2110 -1830 2120
rect 2480 2160 2490 2220
rect 2550 2160 2560 2220
rect 2480 2140 2560 2160
rect 2480 2080 2490 2140
rect 2550 2080 2560 2140
rect 2480 2070 2560 2080
rect -2370 1950 -2360 2010
rect -2300 1950 -2290 2010
rect -2370 1940 -2290 1950
rect -1960 2010 -1880 2020
rect -1960 1950 -1950 2010
rect -1890 1950 -1880 2010
rect -2640 1840 -2630 1900
rect -2570 1840 -2560 1900
rect -2640 1830 -2560 1840
rect -2320 1670 -2240 1680
rect -2320 1610 -2310 1670
rect -2250 1610 -2240 1670
rect -2320 0 -2240 1610
rect -2310 -10 -2240 0
rect -2310 -90 -2240 -80
rect -2740 -390 -2670 -386
rect -2740 -470 -2670 -460
rect -2860 -530 -2790 -510
rect -3040 -1390 -2960 -1360
rect -3040 -1430 -3020 -1390
rect -2980 -1430 -2960 -1390
rect -3040 -2530 -2960 -1430
rect -2860 -1788 -2790 -1778
rect -3040 -2590 -3030 -2530
rect -2970 -2590 -2960 -2530
rect -3040 -2610 -2960 -2590
rect -3040 -2670 -3030 -2610
rect -2970 -2670 -2960 -2610
rect -3040 -2690 -2960 -2670
rect -3040 -2750 -3030 -2690
rect -2970 -2750 -2960 -2690
rect -3040 -2760 -2960 -2750
rect -2870 -2800 -2790 -1858
rect -2500 -1998 -2430 -1988
rect -2500 -2530 -2420 -2068
rect -2500 -2590 -2490 -2530
rect -2430 -2590 -2420 -2530
rect -2500 -2610 -2420 -2590
rect -2500 -2670 -2490 -2610
rect -2430 -2670 -2420 -2610
rect -2500 -2690 -2420 -2670
rect -2500 -2750 -2490 -2690
rect -2430 -2750 -2420 -2690
rect -2500 -2760 -2420 -2750
rect -2070 -2148 -2000 -2138
rect -2070 -2220 -2000 -2218
rect -2070 -2530 -1990 -2220
rect -2070 -2590 -2060 -2530
rect -2000 -2590 -1990 -2530
rect -2070 -2610 -1990 -2590
rect -2070 -2670 -2060 -2610
rect -2000 -2670 -1990 -2610
rect -2070 -2690 -1990 -2670
rect -2070 -2750 -2060 -2690
rect -2000 -2750 -1990 -2690
rect -2070 -2760 -1990 -2750
rect -2870 -2860 -2860 -2800
rect -2800 -2860 -2790 -2800
rect -2870 -2870 -2790 -2860
rect -1960 -2870 -1880 1950
rect 2820 1900 2900 1910
rect 2820 1840 2830 1900
rect 2890 1840 2900 1900
rect -1850 1780 -1770 1790
rect -1850 1720 -1840 1780
rect -1780 1720 -1770 1780
rect -448 1720 -438 1790
rect -368 1720 -358 1790
rect 950 1720 960 1790
rect 1030 1720 1040 1790
rect -1850 -420 -1770 1720
rect 960 1670 1040 1720
rect 960 1610 970 1670
rect 1030 1610 1040 1670
rect 960 1600 1040 1610
rect 2350 1590 2430 1600
rect 2350 1530 2360 1590
rect 2420 1530 2430 1590
rect 2350 1520 2430 1530
rect 2700 1590 2780 1600
rect 2700 1530 2710 1590
rect 2770 1530 2780 1590
rect 2700 1520 2780 1530
rect -1850 -480 -1840 -420
rect -1780 -480 -1770 -420
rect -1850 -490 -1770 -480
rect -1420 1170 2000 1260
rect -1420 1136 -1330 1170
rect -1296 1136 -1230 1170
rect -1196 1136 -1130 1170
rect -1096 1136 -1030 1170
rect -996 1136 -930 1170
rect -896 1136 -830 1170
rect -796 1136 30 1170
rect 64 1136 130 1170
rect 164 1136 230 1170
rect 264 1136 330 1170
rect 364 1136 430 1170
rect 464 1136 530 1170
rect 564 1136 1390 1170
rect 1424 1136 1490 1170
rect 1524 1136 1590 1170
rect 1624 1136 1690 1170
rect 1724 1136 1790 1170
rect 1824 1136 1890 1170
rect 1924 1136 2000 1170
rect -1420 1070 2000 1136
rect -1420 1036 -1330 1070
rect -1296 1036 -1230 1070
rect -1196 1036 -1130 1070
rect -1096 1036 -1030 1070
rect -996 1036 -930 1070
rect -896 1036 -830 1070
rect -796 1036 30 1070
rect 64 1036 130 1070
rect 164 1036 230 1070
rect 264 1036 330 1070
rect 364 1036 430 1070
rect 464 1036 530 1070
rect 564 1036 1390 1070
rect 1424 1036 1490 1070
rect 1524 1036 1590 1070
rect 1624 1036 1690 1070
rect 1724 1036 1790 1070
rect 1824 1036 1890 1070
rect 1924 1036 2000 1070
rect -1420 970 2000 1036
rect -1420 936 -1330 970
rect -1296 936 -1230 970
rect -1196 936 -1130 970
rect -1096 936 -1030 970
rect -996 936 -930 970
rect -896 936 -830 970
rect -796 936 30 970
rect 64 936 130 970
rect 164 936 230 970
rect 264 936 330 970
rect 364 936 430 970
rect 464 936 530 970
rect 564 936 1390 970
rect 1424 936 1490 970
rect 1524 936 1590 970
rect 1624 936 1690 970
rect 1724 936 1790 970
rect 1824 936 1890 970
rect 1924 936 2000 970
rect -1420 870 2000 936
rect -1420 836 -1330 870
rect -1296 836 -1230 870
rect -1196 836 -1130 870
rect -1096 836 -1030 870
rect -996 836 -930 870
rect -896 836 -830 870
rect -796 836 30 870
rect 64 836 130 870
rect 164 836 230 870
rect 264 836 330 870
rect 364 836 430 870
rect 464 836 530 870
rect 564 836 1390 870
rect 1424 836 1490 870
rect 1524 836 1590 870
rect 1624 836 1690 870
rect 1724 836 1790 870
rect 1824 836 1890 870
rect 1924 836 2000 870
rect -1420 770 2000 836
rect -1420 736 -1330 770
rect -1296 736 -1230 770
rect -1196 736 -1130 770
rect -1096 736 -1030 770
rect -996 736 -930 770
rect -896 736 -830 770
rect -796 736 30 770
rect 64 736 130 770
rect 164 736 230 770
rect 264 736 330 770
rect 364 736 430 770
rect 464 736 530 770
rect 564 736 1390 770
rect 1424 736 1490 770
rect 1524 736 1590 770
rect 1624 736 1690 770
rect 1724 736 1790 770
rect 1824 736 1890 770
rect 1924 736 2000 770
rect -1420 670 2000 736
rect -1420 636 -1330 670
rect -1296 636 -1230 670
rect -1196 636 -1130 670
rect -1096 636 -1030 670
rect -996 636 -930 670
rect -896 636 -830 670
rect -796 636 30 670
rect 64 636 130 670
rect 164 636 230 670
rect 264 636 330 670
rect 364 636 430 670
rect 464 636 530 670
rect 564 636 1390 670
rect 1424 636 1490 670
rect 1524 636 1590 670
rect 1624 636 1690 670
rect 1724 636 1790 670
rect 1824 636 1890 670
rect 1924 636 2000 670
rect -1420 560 2000 636
rect -1420 -190 -720 560
rect -1420 -224 -1330 -190
rect -1296 -224 -1230 -190
rect -1196 -224 -1130 -190
rect -1096 -224 -1030 -190
rect -996 -224 -930 -190
rect -896 -224 -830 -190
rect -796 -224 -720 -190
rect -1420 -290 -720 -224
rect -1420 -324 -1330 -290
rect -1296 -324 -1230 -290
rect -1196 -324 -1130 -290
rect -1096 -324 -1030 -290
rect -996 -324 -930 -290
rect -896 -324 -830 -290
rect -796 -324 -720 -290
rect -1420 -390 -720 -324
rect -1420 -420 -1330 -390
rect -1420 -480 -1410 -420
rect -1350 -424 -1330 -420
rect -1296 -424 -1230 -390
rect -1196 -424 -1130 -390
rect -1096 -424 -1030 -390
rect -996 -424 -930 -390
rect -896 -424 -830 -390
rect -796 -424 -720 -390
rect -1350 -480 -720 -424
rect -1420 -490 -720 -480
rect -1420 -524 -1330 -490
rect -1296 -524 -1230 -490
rect -1196 -524 -1130 -490
rect -1096 -524 -1030 -490
rect -996 -524 -930 -490
rect -896 -524 -830 -490
rect -796 -524 -720 -490
rect -1420 -590 -720 -524
rect -1420 -624 -1330 -590
rect -1296 -624 -1230 -590
rect -1196 -624 -1130 -590
rect -1096 -624 -1030 -590
rect -996 -624 -930 -590
rect -896 -624 -830 -590
rect -796 -624 -720 -590
rect -1420 -690 -720 -624
rect -1420 -724 -1330 -690
rect -1296 -724 -1230 -690
rect -1196 -724 -1130 -690
rect -1096 -724 -1030 -690
rect -996 -724 -930 -690
rect -896 -724 -830 -690
rect -796 -724 -720 -690
rect -1420 -1460 -720 -724
rect -60 -190 640 -100
rect -60 -224 30 -190
rect 64 -224 130 -190
rect 164 -224 230 -190
rect 264 -224 330 -190
rect 364 -224 430 -190
rect 464 -224 530 -190
rect 564 -224 640 -190
rect -60 -290 640 -224
rect -60 -324 30 -290
rect 64 -324 130 -290
rect 164 -324 230 -290
rect 264 -324 330 -290
rect 364 -324 430 -290
rect 464 -324 530 -290
rect 564 -324 640 -290
rect -60 -390 640 -324
rect -60 -424 30 -390
rect 64 -424 130 -390
rect 164 -424 230 -390
rect 264 -420 330 -390
rect 320 -424 330 -420
rect 364 -424 430 -390
rect 464 -424 530 -390
rect 564 -424 640 -390
rect -60 -480 260 -424
rect 320 -480 640 -424
rect -60 -490 640 -480
rect -60 -524 30 -490
rect 64 -524 130 -490
rect 164 -524 230 -490
rect 264 -524 330 -490
rect 364 -524 430 -490
rect 464 -524 530 -490
rect 564 -524 640 -490
rect -60 -590 640 -524
rect -60 -624 30 -590
rect 64 -624 130 -590
rect 164 -624 230 -590
rect 264 -624 330 -590
rect 364 -624 430 -590
rect 464 -624 530 -590
rect 564 -624 640 -590
rect -60 -690 640 -624
rect -60 -724 30 -690
rect 64 -724 130 -690
rect 164 -724 230 -690
rect 264 -724 330 -690
rect 364 -724 430 -690
rect 464 -724 530 -690
rect 564 -724 640 -690
rect -60 -800 640 -724
rect 1300 -190 2000 560
rect 1300 -224 1390 -190
rect 1424 -224 1490 -190
rect 1524 -224 1590 -190
rect 1624 -224 1690 -190
rect 1724 -224 1790 -190
rect 1824 -224 1890 -190
rect 1924 -224 2000 -190
rect 1300 -290 2000 -224
rect 1300 -324 1390 -290
rect 1424 -324 1490 -290
rect 1524 -324 1590 -290
rect 1624 -324 1690 -290
rect 1724 -324 1790 -290
rect 1824 -324 1890 -290
rect 1924 -324 2000 -290
rect 1300 -390 2000 -324
rect 1300 -424 1390 -390
rect 1424 -424 1490 -390
rect 1524 -424 1590 -390
rect 1624 -424 1690 -390
rect 1724 -424 1790 -390
rect 1824 -424 1890 -390
rect 1924 -424 2000 -390
rect 2370 -410 2410 1520
rect 2720 0 2760 1520
rect 2700 -10 2770 0
rect 2700 -90 2770 -80
rect 1300 -490 2000 -424
rect 2350 -420 2430 -410
rect 2350 -480 2360 -420
rect 2420 -480 2430 -420
rect 2350 -490 2430 -480
rect 1300 -524 1390 -490
rect 1424 -524 1490 -490
rect 1524 -524 1590 -490
rect 1624 -524 1690 -490
rect 1724 -524 1790 -490
rect 1824 -524 1890 -490
rect 1924 -524 2000 -490
rect 1300 -590 2000 -524
rect 1300 -624 1390 -590
rect 1424 -624 1490 -590
rect 1524 -624 1590 -590
rect 1624 -624 1690 -590
rect 1724 -624 1790 -590
rect 1824 -624 1890 -590
rect 1924 -624 2000 -590
rect 1300 -690 2000 -624
rect 1300 -724 1390 -690
rect 1424 -724 1490 -690
rect 1524 -724 1590 -690
rect 1624 -724 1690 -690
rect 1724 -724 1790 -690
rect 1824 -724 1890 -690
rect 1924 -724 2000 -690
rect 1300 -1460 2000 -724
rect 2820 -850 2900 1840
rect 3180 1800 3220 3570
rect 3160 1790 3240 1800
rect 3160 1730 3170 1790
rect 3230 1730 3240 1790
rect 3160 1720 3240 1730
rect 3270 1600 3310 3800
rect 3250 1590 3330 1600
rect 3250 1530 3260 1590
rect 3320 1530 3330 1590
rect 3250 1520 3330 1530
rect 3480 -360 3560 4750
rect 3590 4350 3830 4360
rect 3590 4290 3600 4350
rect 3660 4290 3680 4350
rect 3740 4290 3760 4350
rect 3820 4290 3830 4350
rect 3590 4270 3830 4290
rect 3590 4210 3600 4270
rect 3660 4210 3680 4270
rect 3740 4210 3760 4270
rect 3820 4210 3830 4270
rect 3590 4190 3830 4210
rect 3590 4130 3600 4190
rect 3660 4130 3680 4190
rect 3740 4130 3760 4190
rect 3820 4130 3830 4190
rect 3590 1040 3830 4130
rect 5250 3600 5330 6290
rect 9330 6280 9410 7180
rect 5710 6030 5790 6050
rect 5710 5980 5730 6030
rect 5770 5980 5790 6030
rect 5710 5890 5790 5980
rect 5710 5840 5730 5890
rect 5770 5840 5790 5890
rect 5510 5760 5590 5780
rect 5510 5720 5530 5760
rect 5570 5720 5590 5760
rect 5510 5620 5590 5720
rect 5510 5560 5520 5620
rect 5580 5560 5590 5620
rect 5510 5550 5590 5560
rect 5710 5620 5790 5840
rect 6110 6030 6190 6050
rect 6110 5980 6130 6030
rect 6170 5980 6190 6030
rect 6110 5890 6190 5980
rect 6110 5840 6130 5890
rect 6170 5840 6190 5890
rect 5710 5560 5720 5620
rect 5780 5560 5790 5620
rect 5710 5550 5790 5560
rect 5950 5620 6030 5630
rect 5950 5560 5960 5620
rect 6020 5560 6030 5620
rect 5950 5550 6030 5560
rect 6110 5620 6190 5840
rect 6110 5560 6120 5620
rect 6180 5560 6190 5620
rect 6110 5550 6190 5560
rect 6510 6030 6590 6050
rect 6510 5980 6530 6030
rect 6570 5980 6590 6030
rect 6510 5890 6590 5980
rect 6510 5840 6530 5890
rect 6570 5840 6590 5890
rect 6510 5620 6590 5840
rect 6510 5560 6520 5620
rect 6580 5560 6590 5620
rect 6510 5550 6590 5560
rect 6910 6030 6990 6050
rect 6910 5980 6930 6030
rect 6970 5980 6990 6030
rect 6910 5890 6990 5980
rect 6910 5840 6930 5890
rect 6970 5840 6990 5890
rect 6910 5620 6990 5840
rect 7310 6030 7390 6050
rect 7310 5980 7330 6030
rect 7370 5980 7390 6030
rect 7310 5890 7390 5980
rect 7310 5840 7330 5890
rect 7370 5840 7390 5890
rect 6910 5560 6920 5620
rect 6980 5560 6990 5620
rect 6910 5550 6990 5560
rect 7090 5730 7170 5740
rect 7090 5670 7100 5730
rect 7160 5670 7170 5730
rect 7090 5510 7170 5670
rect 7310 5620 7390 5840
rect 7310 5560 7320 5620
rect 7380 5560 7390 5620
rect 7310 5550 7390 5560
rect 7510 5760 7590 5780
rect 7510 5720 7530 5760
rect 7570 5720 7590 5760
rect 7510 5620 7590 5720
rect 7510 5560 7520 5620
rect 7580 5560 7590 5620
rect 7510 5550 7590 5560
rect 8230 5620 8310 5630
rect 8230 5560 8240 5620
rect 8300 5560 8310 5620
rect 8230 5550 8310 5560
rect 7090 5450 7100 5510
rect 7160 5450 7170 5510
rect 7090 5440 7170 5450
rect 5560 5340 5640 5360
rect 5560 5300 5580 5340
rect 5620 5300 5640 5340
rect 5560 5280 5640 5300
rect 5690 5340 5770 5360
rect 5690 5300 5710 5340
rect 5750 5300 5770 5340
rect 5690 5280 5770 5300
rect 5820 5340 5900 5360
rect 5820 5300 5840 5340
rect 5880 5300 5900 5340
rect 5820 5220 5900 5300
rect 5950 5340 6030 5360
rect 5950 5300 5970 5340
rect 6010 5300 6030 5340
rect 5950 5280 6030 5300
rect 6080 5340 6160 5360
rect 6080 5300 6100 5340
rect 6140 5300 6160 5340
rect 6080 5240 6160 5300
rect 6210 5340 6290 5360
rect 6210 5300 6230 5340
rect 6270 5300 6290 5340
rect 6210 5280 6290 5300
rect 6340 5340 6420 5360
rect 6340 5300 6360 5340
rect 6400 5300 6420 5340
rect 6340 5280 6420 5300
rect 6700 5340 6780 5360
rect 6700 5300 6720 5340
rect 6760 5300 6780 5340
rect 6700 5280 6780 5300
rect 6830 5340 6910 5360
rect 6830 5300 6850 5340
rect 6890 5300 6910 5340
rect 6830 5280 6910 5300
rect 6960 5340 7040 5360
rect 6960 5300 6980 5340
rect 7020 5300 7040 5340
rect 6960 5280 7040 5300
rect 7090 5340 7170 5360
rect 7090 5300 7110 5340
rect 7150 5300 7170 5340
rect 7090 5280 7170 5300
rect 7220 5340 7300 5360
rect 7220 5300 7240 5340
rect 7280 5300 7300 5340
rect 7220 5280 7300 5300
rect 7350 5340 7430 5360
rect 7350 5300 7370 5340
rect 7410 5300 7430 5340
rect 7350 5280 7430 5300
rect 7480 5340 7560 5360
rect 7480 5300 7500 5340
rect 7540 5300 7560 5340
rect 7480 5280 7560 5300
rect 5820 5180 5840 5220
rect 5880 5180 5900 5220
rect 5820 5160 5900 5180
rect 5730 4890 5810 4900
rect 5730 4830 5740 4890
rect 5800 4830 5810 4890
rect 5730 4820 5810 4830
rect 5840 4780 5880 5160
rect 6100 5060 6140 5240
rect 6870 5230 6950 5240
rect 6870 5170 6880 5230
rect 6940 5170 6950 5230
rect 6170 5160 6250 5170
rect 6170 5100 6180 5160
rect 6240 5100 6250 5160
rect 6170 5090 6250 5100
rect 6870 5160 6950 5170
rect 6080 5000 6090 5060
rect 6150 5000 6160 5060
rect 6100 4780 6140 5000
rect 6190 4900 6230 5090
rect 6870 4980 6910 5160
rect 6830 4920 6840 4980
rect 6900 4920 6910 4980
rect 6980 4910 7020 5280
rect 7240 4920 7280 5280
rect 7310 5230 7390 5240
rect 7310 5170 7320 5230
rect 7380 5170 7390 5230
rect 7310 5160 7390 5170
rect 8850 5230 8930 5240
rect 8850 5170 8860 5230
rect 8920 5170 8930 5230
rect 8850 5160 8930 5170
rect 9330 5230 9410 6130
rect 9550 5330 9660 5350
rect 9550 5260 9570 5330
rect 9640 5260 9660 5330
rect 9550 5240 9660 5260
rect 9330 5170 9340 5230
rect 9400 5170 9410 5230
rect 9330 5160 9410 5170
rect 8010 5110 8090 5120
rect 8010 5050 8020 5110
rect 8080 5050 8090 5110
rect 8010 5040 8090 5050
rect 9720 5060 9800 5070
rect 9720 5000 9730 5060
rect 9790 5000 9800 5060
rect 9720 4990 9800 5000
rect 12000 4990 12080 7830
rect 12110 7780 12190 9010
rect 12110 7720 12120 7780
rect 12180 7720 12190 7780
rect 12110 7700 12190 7720
rect 12110 7640 12120 7700
rect 12180 7640 12190 7700
rect 12110 7620 12190 7640
rect 12110 7560 12120 7620
rect 12180 7560 12190 7620
rect 7240 4910 7320 4920
rect 6170 4890 6250 4900
rect 6170 4830 6180 4890
rect 6240 4830 6250 4890
rect 6170 4820 6250 4830
rect 6960 4890 7040 4910
rect 6960 4850 6980 4890
rect 7020 4850 7040 4890
rect 5560 4760 5640 4780
rect 5560 4720 5580 4760
rect 5620 4720 5640 4760
rect 5560 4660 5640 4720
rect 5560 4620 5580 4660
rect 5620 4620 5640 4660
rect 5560 4600 5640 4620
rect 5690 4760 5770 4780
rect 5690 4720 5710 4760
rect 5750 4720 5770 4760
rect 5690 4660 5770 4720
rect 5690 4620 5710 4660
rect 5750 4620 5770 4660
rect 5690 4600 5770 4620
rect 5820 4760 5900 4780
rect 5820 4720 5840 4760
rect 5880 4720 5900 4760
rect 5820 4660 5900 4720
rect 5820 4620 5840 4660
rect 5880 4620 5900 4660
rect 5820 4600 5900 4620
rect 5950 4760 6030 4780
rect 5950 4720 5970 4760
rect 6010 4720 6030 4760
rect 5950 4660 6030 4720
rect 5950 4620 5970 4660
rect 6010 4620 6030 4660
rect 5950 4600 6030 4620
rect 6080 4760 6160 4780
rect 6080 4720 6100 4760
rect 6140 4720 6160 4760
rect 6080 4660 6160 4720
rect 6080 4620 6100 4660
rect 6140 4620 6160 4660
rect 6080 4600 6160 4620
rect 6210 4760 6290 4780
rect 6210 4720 6230 4760
rect 6270 4720 6290 4760
rect 6210 4660 6290 4720
rect 6210 4620 6230 4660
rect 6270 4620 6290 4660
rect 6210 4600 6290 4620
rect 6340 4760 6420 4780
rect 6340 4720 6360 4760
rect 6400 4720 6420 4760
rect 6340 4660 6420 4720
rect 6340 4620 6360 4660
rect 6400 4620 6420 4660
rect 6340 4600 6420 4620
rect 6700 4760 6780 4780
rect 6700 4720 6720 4760
rect 6760 4720 6780 4760
rect 6700 4660 6780 4720
rect 6700 4620 6720 4660
rect 6760 4620 6780 4660
rect 6700 4600 6780 4620
rect 6830 4760 6910 4780
rect 6830 4720 6850 4760
rect 6890 4720 6910 4760
rect 6830 4660 6910 4720
rect 6830 4620 6850 4660
rect 6890 4620 6910 4660
rect 6830 4600 6910 4620
rect 6960 4760 7040 4850
rect 7240 4850 7250 4910
rect 7310 4850 7320 4910
rect 7240 4840 7320 4850
rect 8010 4890 8090 4900
rect 7240 4780 7280 4840
rect 8010 4830 8020 4890
rect 8080 4830 8090 4890
rect 8010 4820 8090 4830
rect 8850 4890 8930 4900
rect 8850 4830 8860 4890
rect 8920 4830 8930 4890
rect 8850 4820 8930 4830
rect 9330 4890 9410 4900
rect 9330 4830 9340 4890
rect 9400 4830 9410 4890
rect 6960 4720 6980 4760
rect 7020 4720 7040 4760
rect 6960 4660 7040 4720
rect 6960 4620 6980 4660
rect 7020 4620 7040 4660
rect 6960 4600 7040 4620
rect 7090 4760 7170 4780
rect 7090 4720 7110 4760
rect 7150 4720 7170 4760
rect 7090 4660 7170 4720
rect 7090 4620 7110 4660
rect 7150 4620 7170 4660
rect 7090 4600 7170 4620
rect 7220 4760 7300 4780
rect 7220 4720 7240 4760
rect 7280 4720 7300 4760
rect 7220 4660 7300 4720
rect 7220 4620 7240 4660
rect 7280 4620 7300 4660
rect 7220 4600 7300 4620
rect 7350 4760 7430 4780
rect 7350 4720 7370 4760
rect 7410 4720 7430 4760
rect 7350 4660 7430 4720
rect 7350 4620 7370 4660
rect 7410 4620 7430 4660
rect 7350 4600 7430 4620
rect 7480 4760 7560 4780
rect 7480 4720 7500 4760
rect 7540 4720 7560 4760
rect 7480 4660 7560 4720
rect 7480 4620 7500 4660
rect 7540 4620 7560 4660
rect 7480 4600 7560 4620
rect 6030 4510 6110 4520
rect 6030 4450 6040 4510
rect 6100 4450 6110 4510
rect 5630 4400 5710 4410
rect 5630 4340 5640 4400
rect 5700 4340 5710 4400
rect 5630 4230 5710 4340
rect 5630 4190 5650 4230
rect 5690 4190 5710 4230
rect 5630 4170 5710 4190
rect 5830 4400 5910 4410
rect 5830 4340 5840 4400
rect 5900 4340 5910 4400
rect 5630 4110 5710 4130
rect 5630 4070 5650 4110
rect 5690 4070 5710 4110
rect 5630 4010 5710 4070
rect 5630 3970 5650 4010
rect 5690 3970 5710 4010
rect 5630 3910 5710 3970
rect 5630 3870 5650 3910
rect 5690 3870 5710 3910
rect 5630 3810 5710 3870
rect 5630 3770 5650 3810
rect 5690 3770 5710 3810
rect 5630 3710 5710 3770
rect 5630 3670 5650 3710
rect 5690 3670 5710 3710
rect 5630 3650 5710 3670
rect 5830 4110 5910 4340
rect 5830 4070 5850 4110
rect 5890 4070 5910 4110
rect 5830 4010 5910 4070
rect 5830 3970 5850 4010
rect 5890 3970 5910 4010
rect 5830 3910 5910 3970
rect 5830 3870 5850 3910
rect 5890 3870 5910 3910
rect 5830 3810 5910 3870
rect 5830 3770 5850 3810
rect 5890 3770 5910 3810
rect 5830 3710 5910 3770
rect 5830 3670 5850 3710
rect 5890 3670 5910 3710
rect 5830 3650 5910 3670
rect 6030 4260 6110 4450
rect 6030 4200 6040 4260
rect 6100 4200 6110 4260
rect 6030 4110 6110 4200
rect 6030 4070 6050 4110
rect 6090 4070 6110 4110
rect 6030 4010 6110 4070
rect 6030 3970 6050 4010
rect 6090 3970 6110 4010
rect 6030 3910 6110 3970
rect 6030 3870 6050 3910
rect 6090 3870 6110 3910
rect 6030 3810 6110 3870
rect 6030 3770 6050 3810
rect 6090 3770 6110 3810
rect 6030 3710 6110 3770
rect 6030 3670 6050 3710
rect 6090 3670 6110 3710
rect 6030 3650 6110 3670
rect 6230 4400 6310 4410
rect 6230 4340 6240 4400
rect 6300 4340 6310 4400
rect 6230 4110 6310 4340
rect 6630 4400 6710 4410
rect 6630 4340 6640 4400
rect 6700 4340 6710 4400
rect 6230 4070 6250 4110
rect 6290 4070 6310 4110
rect 6230 4010 6310 4070
rect 6230 3970 6250 4010
rect 6290 3970 6310 4010
rect 6230 3910 6310 3970
rect 6230 3870 6250 3910
rect 6290 3870 6310 3910
rect 6230 3810 6310 3870
rect 6230 3770 6250 3810
rect 6290 3770 6310 3810
rect 6230 3710 6310 3770
rect 6230 3670 6250 3710
rect 6290 3670 6310 3710
rect 6230 3650 6310 3670
rect 6430 4110 6510 4130
rect 6430 4070 6450 4110
rect 6490 4070 6510 4110
rect 6430 4010 6510 4070
rect 6430 3970 6450 4010
rect 6490 3970 6510 4010
rect 6430 3910 6510 3970
rect 6430 3870 6450 3910
rect 6490 3870 6510 3910
rect 6430 3810 6510 3870
rect 6430 3770 6450 3810
rect 6490 3770 6510 3810
rect 6430 3710 6510 3770
rect 6430 3670 6450 3710
rect 6490 3670 6510 3710
rect 5250 3540 5260 3600
rect 5320 3540 5330 3600
rect 5250 3530 5330 3540
rect 6430 3600 6510 3670
rect 6630 4110 6710 4340
rect 7030 4400 7190 4410
rect 7030 4340 7040 4400
rect 7100 4340 7120 4400
rect 7180 4340 7190 4400
rect 7030 4330 7190 4340
rect 7430 4400 7510 4410
rect 7430 4340 7440 4400
rect 7500 4340 7510 4400
rect 6630 4070 6650 4110
rect 6690 4070 6710 4110
rect 6630 4010 6710 4070
rect 6630 3970 6650 4010
rect 6690 3970 6710 4010
rect 6630 3910 6710 3970
rect 6630 3870 6650 3910
rect 6690 3870 6710 3910
rect 6630 3810 6710 3870
rect 6630 3770 6650 3810
rect 6690 3770 6710 3810
rect 6630 3710 6710 3770
rect 6630 3670 6650 3710
rect 6690 3670 6710 3710
rect 6630 3650 6710 3670
rect 6830 4110 6910 4130
rect 6830 4070 6850 4110
rect 6890 4070 6910 4110
rect 6830 4010 6910 4070
rect 6830 3970 6850 4010
rect 6890 3970 6910 4010
rect 6830 3910 6910 3970
rect 6830 3870 6850 3910
rect 6890 3870 6910 3910
rect 6830 3810 6910 3870
rect 6830 3770 6850 3810
rect 6890 3770 6910 3810
rect 6830 3710 6910 3770
rect 6830 3670 6850 3710
rect 6890 3670 6910 3710
rect 6430 3540 6440 3600
rect 6500 3540 6510 3600
rect 6430 3530 6510 3540
rect 6830 3600 6910 3670
rect 7030 4110 7110 4330
rect 7030 4070 7050 4110
rect 7090 4070 7110 4110
rect 7030 4010 7110 4070
rect 7030 3970 7050 4010
rect 7090 3970 7110 4010
rect 7030 3910 7110 3970
rect 7030 3870 7050 3910
rect 7090 3870 7110 3910
rect 7030 3810 7110 3870
rect 7030 3770 7050 3810
rect 7090 3770 7110 3810
rect 7030 3710 7110 3770
rect 7030 3670 7050 3710
rect 7090 3670 7110 3710
rect 7030 3650 7110 3670
rect 7230 4260 7310 4270
rect 7230 4200 7240 4260
rect 7300 4200 7310 4260
rect 7230 4110 7310 4200
rect 7230 4070 7250 4110
rect 7290 4070 7310 4110
rect 7230 4010 7310 4070
rect 7230 3970 7250 4010
rect 7290 3970 7310 4010
rect 7230 3910 7310 3970
rect 7230 3870 7250 3910
rect 7290 3870 7310 3910
rect 7230 3810 7310 3870
rect 7230 3770 7250 3810
rect 7290 3770 7310 3810
rect 7230 3710 7310 3770
rect 7230 3670 7250 3710
rect 7290 3670 7310 3710
rect 7230 3650 7310 3670
rect 7430 4110 7510 4340
rect 7430 4070 7450 4110
rect 7490 4070 7510 4110
rect 7430 4010 7510 4070
rect 7430 3970 7450 4010
rect 7490 3970 7510 4010
rect 7430 3910 7510 3970
rect 7430 3870 7450 3910
rect 7490 3870 7510 3910
rect 7430 3810 7510 3870
rect 7430 3770 7450 3810
rect 7490 3770 7510 3810
rect 7430 3710 7510 3770
rect 7430 3670 7450 3710
rect 7490 3670 7510 3710
rect 7430 3650 7510 3670
rect 7630 4400 7710 4410
rect 7630 4340 7640 4400
rect 7700 4340 7710 4400
rect 7630 4230 7710 4340
rect 8230 4400 8310 4410
rect 8230 4340 8240 4400
rect 8300 4340 8310 4400
rect 8230 4330 8310 4340
rect 7630 4190 7650 4230
rect 7690 4190 7710 4230
rect 7630 4110 7710 4190
rect 7630 4070 7650 4110
rect 7690 4070 7710 4110
rect 7630 4010 7710 4070
rect 7630 3970 7650 4010
rect 7690 3970 7710 4010
rect 7630 3910 7710 3970
rect 7630 3870 7650 3910
rect 7690 3870 7710 3910
rect 7630 3810 7710 3870
rect 9330 3810 9410 4830
rect 9550 4820 9660 4840
rect 9550 4750 9570 4820
rect 9640 4750 9660 4820
rect 9550 4730 9660 4750
rect 7630 3770 7650 3810
rect 7690 3770 7710 3810
rect 7630 3710 7710 3770
rect 7630 3670 7650 3710
rect 7690 3670 7710 3710
rect 7630 3650 7710 3670
rect 6830 3540 6840 3600
rect 6900 3540 6910 3600
rect 6830 3530 6910 3540
rect 9120 3210 9200 3220
rect 9120 3150 9130 3210
rect 9190 3150 9200 3210
rect 9120 3140 9200 3150
rect 4150 2970 4390 2990
rect 4150 2910 4190 2970
rect 4250 2910 4290 2970
rect 4350 2910 4390 2970
rect 4150 2890 4390 2910
rect 9330 2900 9410 3610
rect 3590 980 3600 1040
rect 3660 980 3680 1040
rect 3740 980 3760 1040
rect 3820 980 3830 1040
rect 3590 960 3830 980
rect 3980 2010 4060 2020
rect 3980 1950 3990 2010
rect 4050 1950 4060 2010
rect 3480 -420 3490 -360
rect 3550 -420 3560 -360
rect 3480 -640 3560 -420
rect 3860 340 3940 350
rect 3860 280 3870 340
rect 3930 280 3940 340
rect 3480 -652 3550 -640
rect 3480 -732 3550 -722
rect 2820 -860 2890 -850
rect 2820 -940 2890 -930
rect -1420 -1550 2000 -1460
rect -1420 -1584 -1330 -1550
rect -1296 -1584 -1230 -1550
rect -1196 -1584 -1130 -1550
rect -1096 -1584 -1030 -1550
rect -996 -1584 -930 -1550
rect -896 -1584 -830 -1550
rect -796 -1584 30 -1550
rect 64 -1584 130 -1550
rect 164 -1584 230 -1550
rect 264 -1584 330 -1550
rect 364 -1584 430 -1550
rect 464 -1584 530 -1550
rect 564 -1584 1390 -1550
rect 1424 -1584 1490 -1550
rect 1524 -1584 1590 -1550
rect 1624 -1584 1690 -1550
rect 1724 -1584 1790 -1550
rect 1824 -1584 1890 -1550
rect 1924 -1584 2000 -1550
rect -1420 -1650 2000 -1584
rect -1420 -1684 -1330 -1650
rect -1296 -1684 -1230 -1650
rect -1196 -1684 -1130 -1650
rect -1096 -1684 -1030 -1650
rect -996 -1684 -930 -1650
rect -896 -1684 -830 -1650
rect -796 -1684 30 -1650
rect 64 -1684 130 -1650
rect 164 -1684 230 -1650
rect 264 -1684 330 -1650
rect 364 -1684 430 -1650
rect 464 -1684 530 -1650
rect 564 -1684 1390 -1650
rect 1424 -1684 1490 -1650
rect 1524 -1684 1590 -1650
rect 1624 -1684 1690 -1650
rect 1724 -1684 1790 -1650
rect 1824 -1684 1890 -1650
rect 1924 -1684 2000 -1650
rect -1420 -1750 2000 -1684
rect -1420 -1784 -1330 -1750
rect -1296 -1784 -1230 -1750
rect -1196 -1784 -1130 -1750
rect -1096 -1784 -1030 -1750
rect -996 -1784 -930 -1750
rect -896 -1784 -830 -1750
rect -796 -1784 30 -1750
rect 64 -1784 130 -1750
rect 164 -1784 230 -1750
rect 264 -1784 330 -1750
rect 364 -1784 430 -1750
rect 464 -1784 530 -1750
rect 564 -1784 1390 -1750
rect 1424 -1784 1490 -1750
rect 1524 -1784 1590 -1750
rect 1624 -1784 1690 -1750
rect 1724 -1784 1790 -1750
rect 1824 -1784 1890 -1750
rect 1924 -1784 2000 -1750
rect -1420 -1850 2000 -1784
rect -1420 -1884 -1330 -1850
rect -1296 -1884 -1230 -1850
rect -1196 -1884 -1130 -1850
rect -1096 -1884 -1030 -1850
rect -996 -1884 -930 -1850
rect -896 -1884 -830 -1850
rect -796 -1884 30 -1850
rect 64 -1884 130 -1850
rect 164 -1884 230 -1850
rect 264 -1884 330 -1850
rect 364 -1884 430 -1850
rect 464 -1884 530 -1850
rect 564 -1884 1390 -1850
rect 1424 -1884 1490 -1850
rect 1524 -1884 1590 -1850
rect 1624 -1884 1690 -1850
rect 1724 -1884 1790 -1850
rect 1824 -1884 1890 -1850
rect 1924 -1884 2000 -1850
rect -1420 -1950 2000 -1884
rect -1420 -1984 -1330 -1950
rect -1296 -1984 -1230 -1950
rect -1196 -1984 -1130 -1950
rect -1096 -1984 -1030 -1950
rect -996 -1984 -930 -1950
rect -896 -1984 -830 -1950
rect -796 -1984 30 -1950
rect 64 -1984 130 -1950
rect 164 -1984 230 -1950
rect 264 -1984 330 -1950
rect 364 -1984 430 -1950
rect 464 -1984 530 -1950
rect 564 -1984 1390 -1950
rect 1424 -1984 1490 -1950
rect 1524 -1984 1590 -1950
rect 1624 -1984 1690 -1950
rect 1724 -1984 1790 -1950
rect 1824 -1984 1890 -1950
rect 1924 -1984 2000 -1950
rect -1420 -2050 2000 -1984
rect 2990 -1450 3070 -1420
rect 2990 -1490 3010 -1450
rect 3050 -1490 3070 -1450
rect -1420 -2084 -1330 -2050
rect -1296 -2084 -1230 -2050
rect -1196 -2084 -1130 -2050
rect -1096 -2084 -1030 -2050
rect -996 -2084 -930 -2050
rect -896 -2084 -830 -2050
rect -796 -2084 30 -2050
rect 64 -2084 130 -2050
rect 164 -2084 230 -2050
rect 264 -2084 330 -2050
rect 364 -2084 430 -2050
rect 464 -2084 530 -2050
rect 564 -2084 1390 -2050
rect 1424 -2084 1490 -2050
rect 1524 -2084 1590 -2050
rect 1624 -2084 1690 -2050
rect 1724 -2084 1790 -2050
rect 1824 -2084 1890 -2050
rect 1924 -2084 2000 -2050
rect -1420 -2160 2000 -2084
rect 2820 -1998 2890 -1988
rect 2460 -2148 2530 -2138
rect 2460 -2520 2530 -2218
rect 2820 -2520 2890 -2068
rect 250 -2530 330 -2520
rect 250 -2590 260 -2530
rect 320 -2590 330 -2530
rect 250 -2610 330 -2590
rect 250 -2670 260 -2610
rect 320 -2670 330 -2610
rect 250 -2690 330 -2670
rect 250 -2750 260 -2690
rect 320 -2750 330 -2690
rect 250 -2760 330 -2750
rect 2450 -2530 2530 -2520
rect 2450 -2590 2460 -2530
rect 2520 -2590 2530 -2530
rect 2450 -2610 2530 -2590
rect 2450 -2670 2460 -2610
rect 2520 -2670 2530 -2610
rect 2450 -2690 2530 -2670
rect 2450 -2750 2460 -2690
rect 2520 -2750 2530 -2690
rect 2450 -2760 2530 -2750
rect 2810 -2530 2890 -2520
rect 2810 -2590 2820 -2530
rect 2880 -2590 2890 -2530
rect 2810 -2610 2890 -2590
rect 2810 -2670 2820 -2610
rect 2880 -2670 2890 -2610
rect 2810 -2690 2890 -2670
rect 2810 -2750 2820 -2690
rect 2880 -2750 2890 -2690
rect 2810 -2760 2890 -2750
rect 2990 -2530 3070 -1490
rect 3480 -1998 3550 -1988
rect 3860 -1990 3940 280
rect 3980 -1740 4060 1950
rect 4090 1040 4190 1060
rect 4090 980 4110 1040
rect 4170 980 4190 1040
rect 4090 960 4190 980
rect 4090 -360 4190 -340
rect 4090 -420 4110 -360
rect 4170 -420 4190 -360
rect 4090 -440 4190 -420
rect 4230 -1060 4310 2890
rect 9320 2880 9420 2900
rect 9320 2820 9340 2880
rect 9400 2820 9420 2880
rect 9320 2800 9420 2820
rect 4230 -1120 4240 -1060
rect 4300 -1120 4310 -1060
rect 4230 -1130 4310 -1120
rect 3970 -1760 4070 -1740
rect 3970 -1820 3990 -1760
rect 4050 -1820 4070 -1760
rect 3970 -1840 4070 -1820
rect 3480 -2080 3550 -2068
rect 3850 -2000 3940 -1990
rect 3850 -2070 3860 -2000
rect 3930 -2070 3940 -2000
rect 3850 -2080 3940 -2070
rect 2990 -2590 3000 -2530
rect 3060 -2590 3070 -2530
rect 2990 -2610 3070 -2590
rect 2990 -2670 3000 -2610
rect 3060 -2670 3070 -2610
rect 2990 -2690 3070 -2670
rect 2990 -2750 3000 -2690
rect 3060 -2750 3070 -2690
rect 2990 -2760 3070 -2750
rect 4300 -2460 4380 -2450
rect 4300 -2520 4310 -2460
rect 4370 -2520 4380 -2460
rect 4300 -2800 4380 -2520
rect 4300 -2860 4310 -2800
rect 4370 -2860 4380 -2800
rect 4300 -2870 4380 -2860
rect 2890 -2910 2970 -2900
rect 5340 -2910 5420 -2900
rect 2890 -2970 2900 -2910
rect 2960 -2970 2980 -2910
rect 2890 -2980 2980 -2970
rect 5330 -2970 5350 -2910
rect 5410 -2970 5420 -2910
rect 5330 -2980 5420 -2970
rect 12110 -2910 12190 7560
rect 12110 -2970 12120 -2910
rect 12180 -2970 12190 -2910
rect 12110 -2980 12190 -2970
<< via1 >>
rect 9420 14210 9480 14270
rect 8930 14100 8990 14160
rect 9010 14100 9070 14160
rect 9090 14100 9150 14160
rect 8930 14020 8990 14080
rect 9010 14020 9070 14080
rect 9090 14020 9150 14080
rect 8930 13940 8990 14000
rect 9010 13940 9070 14000
rect 9090 13940 9150 14000
rect -1340 13040 -1280 13050
rect -1340 13000 -1330 13040
rect -1330 13000 -1290 13040
rect -1290 13000 -1280 13040
rect -1340 12990 -1280 13000
rect -1120 13040 -1060 13050
rect -1120 13000 -1110 13040
rect -1110 13000 -1070 13040
rect -1070 13000 -1060 13040
rect -1120 12990 -1060 13000
rect -650 13040 -590 13050
rect -650 13000 -640 13040
rect -640 13000 -600 13040
rect -600 13000 -590 13040
rect -650 12990 -590 13000
rect -310 13040 -250 13050
rect -310 13000 -300 13040
rect -300 13000 -260 13040
rect -260 13000 -250 13040
rect -310 12990 -250 13000
rect -90 13040 -30 13050
rect -90 13000 -80 13040
rect -80 13000 -40 13040
rect -40 13000 -30 13040
rect -90 12990 -30 13000
rect 350 13040 410 13050
rect 350 13000 360 13040
rect 360 13000 400 13040
rect 400 13000 410 13040
rect 350 12990 410 13000
rect 1030 13040 1090 13050
rect 1030 13000 1040 13040
rect 1040 13000 1080 13040
rect 1080 13000 1090 13040
rect 1030 12990 1090 13000
rect 1250 13040 1310 13050
rect 1250 13000 1260 13040
rect 1260 13000 1300 13040
rect 1300 13000 1310 13040
rect 1250 12990 1310 13000
rect 1720 13040 1780 13050
rect 1720 13000 1730 13040
rect 1730 13000 1770 13040
rect 1770 13000 1780 13040
rect 1720 12990 1780 13000
rect 2180 13040 2240 13050
rect 2180 13000 2190 13040
rect 2190 13000 2230 13040
rect 2230 13000 2240 13040
rect 2180 12990 2240 13000
rect 2530 13040 2590 13050
rect 2530 13000 2540 13040
rect 2540 13000 2580 13040
rect 2580 13000 2590 13040
rect 2530 12990 2590 13000
rect 2780 13040 2840 13050
rect 2780 13000 2790 13040
rect 2790 13000 2830 13040
rect 2830 13000 2840 13040
rect 2780 12990 2840 13000
rect 3000 13040 3060 13050
rect 3000 13000 3010 13040
rect 3010 13000 3050 13040
rect 3050 13000 3060 13040
rect 3000 12990 3060 13000
rect 3330 13040 3390 13050
rect 3330 13000 3340 13040
rect 3340 13000 3380 13040
rect 3380 13000 3390 13040
rect 3330 12990 3390 13000
rect 3990 13040 4050 13050
rect 3990 13000 4000 13040
rect 4000 13000 4040 13040
rect 4040 13000 4050 13040
rect 3990 12990 4050 13000
rect 4210 13040 4270 13050
rect 4210 13000 4220 13040
rect 4220 13000 4260 13040
rect 4260 13000 4270 13040
rect 4210 12990 4270 13000
rect 4780 13040 4840 13050
rect 4780 13000 4790 13040
rect 4790 13000 4830 13040
rect 4830 13000 4840 13040
rect 4780 12990 4840 13000
rect 5040 13040 5100 13050
rect 5040 13000 5050 13040
rect 5050 13000 5090 13040
rect 5090 13000 5100 13040
rect 5040 12990 5100 13000
rect 5290 13040 5350 13050
rect 5290 13000 5300 13040
rect 5300 13000 5340 13040
rect 5340 13000 5350 13040
rect 5290 12990 5350 13000
rect 5510 13040 5570 13050
rect 5510 13000 5520 13040
rect 5520 13000 5560 13040
rect 5560 13000 5570 13040
rect 5510 12990 5570 13000
rect 6060 13040 6120 13050
rect 6060 13000 6070 13040
rect 6070 13000 6110 13040
rect 6110 13000 6120 13040
rect 6060 12990 6120 13000
rect 6340 13040 6400 13050
rect 6340 13000 6350 13040
rect 6350 13000 6390 13040
rect 6390 13000 6400 13040
rect 6340 12990 6400 13000
rect 6590 13040 6650 13050
rect 6590 13000 6600 13040
rect 6600 13000 6640 13040
rect 6640 13000 6650 13040
rect 6590 12990 6650 13000
rect 6810 13040 6870 13050
rect 6810 13000 6820 13040
rect 6820 13000 6860 13040
rect 6860 13000 6870 13040
rect 6810 12990 6870 13000
rect 7360 13040 7420 13050
rect 7360 13000 7370 13040
rect 7370 13000 7410 13040
rect 7410 13000 7420 13040
rect 7360 12990 7420 13000
rect 7640 13040 7700 13050
rect 7640 13000 7650 13040
rect 7650 13000 7690 13040
rect 7690 13000 7700 13040
rect 7640 12990 7700 13000
rect 7890 13040 7950 13050
rect 7890 13000 7900 13040
rect 7900 13000 7940 13040
rect 7940 13000 7950 13040
rect 7890 12990 7950 13000
rect 8110 13040 8170 13050
rect 8110 13000 8120 13040
rect 8120 13000 8160 13040
rect 8160 13000 8170 13040
rect 8110 12990 8170 13000
rect 8660 13040 8720 13050
rect 8660 13000 8670 13040
rect 8670 13000 8710 13040
rect 8710 13000 8720 13040
rect 8660 12990 8720 13000
rect -1770 12610 -1710 12670
rect -1560 12660 -1500 12670
rect -1560 12620 -1550 12660
rect -1550 12620 -1510 12660
rect -1510 12620 -1500 12660
rect -1560 12610 -1500 12620
rect 9940 14210 10000 14270
rect 10460 14210 10520 14270
rect 10950 14210 11010 14270
rect 11280 14100 11340 14160
rect 11360 14100 11420 14160
rect 11440 14100 11500 14160
rect 11280 14020 11340 14080
rect 11360 14020 11420 14080
rect 11440 14020 11500 14080
rect 11280 13940 11340 14000
rect 11360 13940 11420 14000
rect 11440 13940 11500 14000
rect 9370 13542 9422 13552
rect 9370 13508 9378 13542
rect 9378 13508 9412 13542
rect 9412 13508 9422 13542
rect 9370 13500 9422 13508
rect 9890 13542 9942 13552
rect 9890 13508 9898 13542
rect 9898 13508 9932 13542
rect 9932 13508 9942 13542
rect 9890 13500 9942 13508
rect 10410 13542 10462 13552
rect 10410 13508 10418 13542
rect 10418 13508 10452 13542
rect 10452 13508 10462 13542
rect 10410 13500 10462 13508
rect 10976 13542 11028 13552
rect 10976 13508 10986 13542
rect 10986 13508 11020 13542
rect 11020 13508 11028 13542
rect 10976 13500 11028 13508
rect 9420 13380 9480 13390
rect 9420 13340 9430 13380
rect 9430 13340 9470 13380
rect 9470 13340 9480 13380
rect 9420 13330 9480 13340
rect 9420 13280 9480 13290
rect 9420 13240 9430 13280
rect 9430 13240 9470 13280
rect 9470 13240 9480 13280
rect 9420 13230 9480 13240
rect 9630 13330 9690 13390
rect 9630 13230 9690 13290
rect 9384 13162 9436 13172
rect 9384 13128 9392 13162
rect 9392 13128 9426 13162
rect 9426 13128 9436 13162
rect 9384 13120 9436 13128
rect 9520 13110 9580 13170
rect 8930 12700 8990 12760
rect 9010 12700 9070 12760
rect 9090 12700 9150 12760
rect 8866 12662 8918 12672
rect 8866 12628 8874 12662
rect 8874 12628 8908 12662
rect 8908 12628 8918 12662
rect 8866 12620 8918 12628
rect 8930 12620 8990 12680
rect 9010 12620 9070 12680
rect 9090 12620 9150 12680
rect 8930 12540 8990 12600
rect 9010 12540 9070 12600
rect 9090 12540 9150 12600
rect 9350 12700 9410 12760
rect 9350 12620 9410 12680
rect 9350 12540 9410 12600
rect 9440 12700 9500 12760
rect 9440 12620 9500 12680
rect 9440 12540 9500 12600
rect -1180 12260 -1120 12270
rect -1180 12220 -1170 12260
rect -1170 12220 -1130 12260
rect -1130 12220 -1120 12260
rect -1180 12210 -1120 12220
rect -760 12260 -700 12270
rect -760 12220 -750 12260
rect -750 12220 -710 12260
rect -710 12220 -700 12260
rect -760 12210 -700 12220
rect -90 12260 -30 12270
rect -90 12220 -80 12260
rect -80 12220 -40 12260
rect -40 12220 -30 12260
rect -90 12210 -30 12220
rect 480 12260 540 12270
rect 480 12220 490 12260
rect 490 12220 530 12260
rect 530 12220 540 12260
rect 480 12210 540 12220
rect 1190 12260 1250 12270
rect 1190 12220 1200 12260
rect 1200 12220 1240 12260
rect 1240 12220 1250 12260
rect 1190 12210 1250 12220
rect 1620 12260 1680 12270
rect 1620 12220 1630 12260
rect 1630 12220 1670 12260
rect 1670 12220 1680 12260
rect 1620 12210 1680 12220
rect 2060 12260 2120 12270
rect 2060 12220 2070 12260
rect 2070 12220 2110 12260
rect 2110 12220 2120 12260
rect 2060 12210 2120 12220
rect 2310 12260 2370 12270
rect 2310 12220 2320 12260
rect 2320 12220 2360 12260
rect 2360 12220 2370 12260
rect 2310 12210 2370 12220
rect 2530 12260 2590 12270
rect 2530 12220 2540 12260
rect 2540 12220 2580 12260
rect 2580 12220 2590 12260
rect 2530 12210 2590 12220
rect 3000 12260 3060 12270
rect 3000 12220 3010 12260
rect 3010 12220 3050 12260
rect 3050 12220 3060 12260
rect 3000 12210 3060 12220
rect 3440 12260 3500 12270
rect 3440 12220 3450 12260
rect 3450 12220 3490 12260
rect 3490 12220 3500 12260
rect 3440 12210 3500 12220
rect 4060 12260 4120 12270
rect 4060 12220 4070 12260
rect 4070 12220 4110 12260
rect 4110 12220 4120 12260
rect 4060 12210 4120 12220
rect 4400 12260 4460 12270
rect 4400 12220 4410 12260
rect 4410 12220 4450 12260
rect 4450 12220 4460 12260
rect 4400 12210 4460 12220
rect 4760 12260 4820 12270
rect 4760 12220 4770 12260
rect 4770 12220 4810 12260
rect 4810 12220 4820 12260
rect 4760 12210 4820 12220
rect 5360 12260 5420 12270
rect 5360 12220 5370 12260
rect 5370 12220 5410 12260
rect 5410 12220 5420 12260
rect 5360 12210 5420 12220
rect 5700 12260 5760 12270
rect 5700 12220 5710 12260
rect 5710 12220 5750 12260
rect 5750 12220 5760 12260
rect 5700 12210 5760 12220
rect 6060 12260 6120 12270
rect 6060 12220 6070 12260
rect 6070 12220 6110 12260
rect 6110 12220 6120 12260
rect 6060 12210 6120 12220
rect 6660 12260 6720 12270
rect 6660 12220 6670 12260
rect 6670 12220 6710 12260
rect 6710 12220 6720 12260
rect 6660 12210 6720 12220
rect 7000 12260 7060 12270
rect 7000 12220 7010 12260
rect 7010 12220 7050 12260
rect 7050 12220 7060 12260
rect 7000 12210 7060 12220
rect 7360 12260 7420 12270
rect 7360 12220 7370 12260
rect 7370 12220 7410 12260
rect 7410 12220 7420 12260
rect 7360 12210 7420 12220
rect 7960 12260 8020 12270
rect 7960 12220 7970 12260
rect 7970 12220 8010 12260
rect 8010 12220 8020 12260
rect 7960 12210 8020 12220
rect 8300 12260 8360 12270
rect 8300 12220 8310 12260
rect 8310 12220 8350 12260
rect 8350 12220 8360 12260
rect 8300 12210 8360 12220
rect 8660 12260 8720 12270
rect 8660 12220 8670 12260
rect 8670 12220 8710 12260
rect 8710 12220 8720 12260
rect 8660 12210 8720 12220
rect 9384 12072 9436 12082
rect 9384 12038 9392 12072
rect 9392 12038 9426 12072
rect 9426 12038 9436 12072
rect 9384 12030 9436 12038
rect 9940 13380 10000 13390
rect 9940 13340 9950 13380
rect 9950 13340 9990 13380
rect 9990 13340 10000 13380
rect 9940 13330 10000 13340
rect 9940 13280 10000 13290
rect 9940 13240 9950 13280
rect 9950 13240 9990 13280
rect 9990 13240 10000 13280
rect 9940 13230 10000 13240
rect 10150 13330 10210 13390
rect 10150 13230 10210 13290
rect 9904 13162 9956 13172
rect 9904 13128 9912 13162
rect 9912 13128 9946 13162
rect 9946 13128 9956 13162
rect 9904 13120 9956 13128
rect 10040 13110 10100 13170
rect 9870 12700 9930 12760
rect 9870 12620 9930 12680
rect 9870 12540 9930 12600
rect 9960 12700 10020 12760
rect 9960 12620 10020 12680
rect 9960 12540 10020 12600
rect 9630 12030 9690 12090
rect 9420 11960 9480 11970
rect 9420 11920 9430 11960
rect 9430 11920 9470 11960
rect 9470 11920 9480 11960
rect 9420 11910 9480 11920
rect 9520 11910 9580 11970
rect 9904 12072 9956 12082
rect 9904 12038 9912 12072
rect 9912 12038 9946 12072
rect 9946 12038 9956 12072
rect 9904 12030 9956 12038
rect 10460 13380 10520 13390
rect 10460 13340 10470 13380
rect 10470 13340 10510 13380
rect 10510 13340 10520 13380
rect 10460 13330 10520 13340
rect 10460 13280 10520 13290
rect 10460 13240 10470 13280
rect 10470 13240 10510 13280
rect 10510 13240 10520 13280
rect 10460 13230 10520 13240
rect 10670 13330 10730 13390
rect 10670 13230 10730 13290
rect 10424 13162 10476 13172
rect 10424 13128 10432 13162
rect 10432 13128 10466 13162
rect 10466 13128 10476 13162
rect 10424 13120 10476 13128
rect 10560 13110 10620 13170
rect 10390 12700 10450 12760
rect 10390 12620 10450 12680
rect 10390 12540 10450 12600
rect 10480 12700 10540 12760
rect 10480 12620 10540 12680
rect 10480 12540 10540 12600
rect 10150 12030 10210 12090
rect 9420 11520 9480 11580
rect 9690 11520 9750 11580
rect 9500 11390 9560 11400
rect 9500 11350 9510 11390
rect 9510 11350 9550 11390
rect 9550 11350 9560 11390
rect 9500 11340 9560 11350
rect 9940 11960 10000 11970
rect 9940 11920 9950 11960
rect 9950 11920 9990 11960
rect 9990 11920 10000 11960
rect 9940 11910 10000 11920
rect 10040 11910 10100 11970
rect 10424 12072 10476 12082
rect 10424 12038 10432 12072
rect 10432 12038 10466 12072
rect 10466 12038 10476 12072
rect 10424 12030 10476 12038
rect 10670 12030 10730 12090
rect 9940 11520 10000 11580
rect 10210 11520 10270 11580
rect 10020 11390 10080 11400
rect 10020 11350 10030 11390
rect 10030 11350 10070 11390
rect 10070 11350 10080 11390
rect 10020 11340 10080 11350
rect 10460 11960 10520 11970
rect 10460 11920 10470 11960
rect 10470 11920 10510 11960
rect 10510 11920 10520 11960
rect 10460 11910 10520 11920
rect 10560 11910 10620 11970
rect 10460 11520 10520 11580
rect 10730 11520 10790 11580
rect 10540 11390 10600 11400
rect 10540 11350 10550 11390
rect 10550 11350 10590 11390
rect 10590 11350 10600 11390
rect 10540 11340 10600 11350
rect 10870 11340 10930 11400
rect 11280 12700 11340 12760
rect 11360 12700 11420 12760
rect 11440 12700 11500 12760
rect 11280 12620 11340 12680
rect 11360 12620 11420 12680
rect 11440 12620 11500 12680
rect 11280 12540 11340 12600
rect 11360 12540 11420 12600
rect 11440 12540 11500 12600
rect 12120 13490 12180 13550
rect 11060 11390 11120 11400
rect 11060 11350 11070 11390
rect 11070 11350 11110 11390
rect 11110 11350 11120 11390
rect 11060 11340 11120 11350
rect 9690 10690 9750 10750
rect 10210 10690 10270 10750
rect 10730 10690 10790 10750
rect 11250 10690 11310 10750
rect -630 10440 -570 10450
rect -630 10400 -620 10440
rect -620 10400 -580 10440
rect -580 10400 -570 10440
rect -630 10390 -570 10400
rect -410 10440 -350 10450
rect -410 10400 -400 10440
rect -400 10400 -360 10440
rect -360 10400 -350 10440
rect -410 10390 -350 10400
rect -110 10440 -50 10450
rect -110 10400 -100 10440
rect -100 10400 -60 10440
rect -60 10400 -50 10440
rect -110 10390 -50 10400
rect 110 10440 170 10450
rect 110 10400 120 10440
rect 120 10400 160 10440
rect 160 10400 170 10440
rect 110 10390 170 10400
rect 270 10440 330 10450
rect 270 10400 280 10440
rect 280 10400 320 10440
rect 320 10400 330 10440
rect 270 10390 330 10400
rect 490 10440 550 10450
rect 490 10400 500 10440
rect 500 10400 540 10440
rect 540 10400 550 10440
rect 490 10390 550 10400
rect 790 10440 850 10450
rect 790 10400 800 10440
rect 800 10400 840 10440
rect 840 10400 850 10440
rect 790 10390 850 10400
rect 1010 10440 1070 10450
rect 1010 10400 1020 10440
rect 1020 10400 1060 10440
rect 1060 10400 1070 10440
rect 1010 10390 1070 10400
rect 1310 10440 1370 10450
rect 1310 10400 1320 10440
rect 1320 10400 1360 10440
rect 1360 10400 1370 10440
rect 1310 10390 1370 10400
rect 1750 10440 1810 10450
rect 1750 10400 1760 10440
rect 1760 10400 1800 10440
rect 1800 10400 1810 10440
rect 1750 10390 1810 10400
rect 2080 10440 2140 10450
rect 2080 10400 2090 10440
rect 2090 10400 2130 10440
rect 2130 10400 2140 10440
rect 2080 10390 2140 10400
rect 2510 10440 2570 10450
rect 2510 10400 2520 10440
rect 2520 10400 2560 10440
rect 2560 10400 2570 10440
rect 2510 10390 2570 10400
rect 2900 10440 2960 10450
rect 2900 10400 2910 10440
rect 2910 10400 2950 10440
rect 2950 10400 2960 10440
rect 2900 10390 2960 10400
rect 3290 10440 3350 10450
rect 3290 10400 3300 10440
rect 3300 10400 3340 10440
rect 3340 10400 3350 10440
rect 3290 10390 3350 10400
rect 3810 10450 3870 10510
rect -220 10330 -160 10340
rect -220 10290 -210 10330
rect -210 10290 -170 10330
rect -170 10290 -160 10330
rect -220 10280 -160 10290
rect 1500 10330 1560 10340
rect 1500 10290 1510 10330
rect 1510 10290 1550 10330
rect 1550 10290 1560 10330
rect 1500 10280 1560 10290
rect 2350 10260 2410 10320
rect 3580 10330 3640 10340
rect 3580 10290 3590 10330
rect 3590 10290 3630 10330
rect 3630 10290 3640 10330
rect 3580 10280 3640 10290
rect -750 9950 -690 9960
rect -750 9910 -740 9950
rect -740 9910 -700 9950
rect -700 9910 -690 9950
rect -750 9900 -690 9910
rect 1150 9980 1210 9990
rect 1150 9940 1160 9980
rect 1160 9940 1200 9980
rect 1200 9940 1210 9980
rect 1150 9930 1210 9940
rect -630 9260 -570 9270
rect -630 9220 -620 9260
rect -620 9220 -580 9260
rect -580 9220 -570 9260
rect -630 9210 -570 9220
rect 110 9260 170 9270
rect 110 9220 120 9260
rect 120 9220 160 9260
rect 160 9220 170 9260
rect 110 9210 170 9220
rect 270 9260 330 9270
rect 270 9220 280 9260
rect 280 9220 320 9260
rect 320 9220 330 9260
rect 270 9210 330 9220
rect 1010 9260 1070 9270
rect 1010 9220 1020 9260
rect 1020 9220 1060 9260
rect 1060 9220 1070 9260
rect 1010 9210 1070 9220
rect -180 9150 -120 9160
rect -180 9110 -170 9150
rect -170 9110 -130 9150
rect -130 9110 -120 9150
rect -180 9100 -120 9110
rect 2240 9940 2300 9950
rect 2240 9900 2250 9940
rect 2250 9900 2290 9940
rect 2290 9900 2300 9940
rect 2240 9890 2300 9900
rect 9110 10450 9180 10520
rect 4520 10280 4580 10340
rect 4120 9990 4180 10000
rect 4120 9950 4130 9990
rect 4130 9950 4170 9990
rect 4170 9950 4180 9990
rect 4120 9940 4180 9950
rect 4410 9940 4470 10000
rect 1370 9370 1430 9380
rect 1370 9330 1380 9370
rect 1380 9330 1420 9370
rect 1420 9330 1430 9370
rect 1370 9320 1430 9330
rect 1260 9260 1320 9270
rect 1260 9220 1270 9260
rect 1270 9220 1310 9260
rect 1310 9220 1320 9260
rect 1260 9210 1320 9220
rect 1450 9260 1510 9270
rect 1450 9220 1460 9260
rect 1460 9220 1500 9260
rect 1500 9220 1510 9260
rect 1450 9210 1510 9220
rect 1530 9260 1590 9270
rect 1530 9220 1540 9260
rect 1540 9220 1580 9260
rect 1580 9220 1590 9260
rect 1530 9210 1590 9220
rect 1740 9260 1800 9270
rect 1740 9220 1750 9260
rect 1750 9220 1790 9260
rect 1790 9220 1800 9260
rect 1740 9210 1800 9220
rect 2070 9260 2130 9270
rect 2070 9220 2080 9260
rect 2080 9220 2120 9260
rect 2120 9220 2130 9260
rect 2070 9210 2130 9220
rect 1350 9100 1410 9160
rect 3810 9910 3870 9920
rect 3810 9870 3820 9910
rect 3820 9870 3860 9910
rect 3860 9870 3870 9910
rect 3810 9860 3870 9870
rect 2510 9260 2570 9270
rect 2510 9220 2520 9260
rect 2520 9220 2560 9260
rect 2560 9220 2570 9260
rect 2510 9210 2570 9220
rect 2900 9260 2960 9270
rect 2900 9220 2910 9260
rect 2910 9220 2950 9260
rect 2950 9220 2960 9260
rect 2900 9210 2960 9220
rect 3110 9210 3170 9270
rect 3290 9260 3350 9270
rect 3290 9220 3300 9260
rect 3300 9220 3340 9260
rect 3340 9220 3350 9260
rect 3290 9210 3350 9220
rect 3970 9260 4030 9270
rect 3970 9220 3980 9260
rect 3980 9220 4020 9260
rect 4020 9220 4030 9260
rect 3970 9210 4030 9220
rect -1770 8520 -1710 8580
rect -750 8570 -690 8580
rect -750 8530 -740 8570
rect -740 8530 -700 8570
rect -700 8530 -690 8570
rect -750 8520 -690 8530
rect 1170 8580 1230 8590
rect 1170 8540 1180 8580
rect 1180 8540 1220 8580
rect 1220 8540 1230 8580
rect 1170 8530 1230 8540
rect 2200 8580 2260 8590
rect 2200 8540 2210 8580
rect 2210 8540 2250 8580
rect 2250 8540 2260 8580
rect 2200 8530 2260 8540
rect 2350 9090 2410 9150
rect 2770 9100 2830 9160
rect 2940 9150 3000 9160
rect 2940 9110 2950 9150
rect 2950 9110 2990 9150
rect 2990 9110 3000 9150
rect 2940 9100 3000 9110
rect 3580 9150 3640 9160
rect 3580 9110 3590 9150
rect 3590 9110 3630 9150
rect 3630 9110 3640 9150
rect 3580 9100 3640 9110
rect 4300 9100 4360 9160
rect 5660 9940 5720 10000
rect 5880 9940 5940 10000
rect 6320 9940 6380 10000
rect 4520 9170 4580 9230
rect 5040 9290 5100 9350
rect 4410 9060 4470 9120
rect 4300 8950 4360 9010
rect 4770 8950 4830 9010
rect 4850 8950 4910 9010
rect 4930 8950 4990 9010
rect 4300 8840 4360 8900
rect 4120 8530 4180 8540
rect 4120 8490 4130 8530
rect 4130 8490 4170 8530
rect 4170 8490 4180 8530
rect 4120 8480 4180 8490
rect 4300 8480 4360 8540
rect 3020 8190 3080 8200
rect 3020 8150 3030 8190
rect 3030 8150 3070 8190
rect 3070 8150 3080 8190
rect 3020 8140 3080 8150
rect 3650 8190 3710 8200
rect 3650 8150 3660 8190
rect 3660 8150 3700 8190
rect 3700 8150 3710 8190
rect 3650 8140 3710 8150
rect 4220 8140 4280 8200
rect -630 8080 -570 8090
rect -630 8040 -620 8080
rect -620 8040 -580 8080
rect -580 8040 -570 8080
rect -630 8030 -570 8040
rect -410 8080 -350 8090
rect -410 8040 -400 8080
rect -400 8040 -360 8080
rect -360 8040 -350 8080
rect -410 8030 -350 8040
rect -110 8080 -50 8090
rect -110 8040 -100 8080
rect -100 8040 -60 8080
rect -60 8040 -50 8080
rect -110 8030 -50 8040
rect 120 8080 180 8090
rect 120 8040 130 8080
rect 130 8040 170 8080
rect 170 8040 180 8080
rect 120 8030 180 8040
rect 270 8080 330 8090
rect 270 8040 280 8080
rect 280 8040 320 8080
rect 320 8040 330 8080
rect 270 8030 330 8040
rect 490 8080 550 8090
rect 490 8040 500 8080
rect 500 8040 540 8080
rect 540 8040 550 8080
rect 490 8030 550 8040
rect 790 8080 850 8090
rect 790 8040 800 8080
rect 800 8040 840 8080
rect 840 8040 850 8080
rect 790 8030 850 8040
rect 1010 8080 1070 8090
rect 1010 8040 1020 8080
rect 1020 8040 1060 8080
rect 1060 8040 1070 8080
rect 1010 8030 1070 8040
rect 1410 8080 1470 8090
rect 1410 8040 1420 8080
rect 1420 8040 1460 8080
rect 1460 8040 1470 8080
rect 1410 8030 1470 8040
rect 1740 8080 1800 8090
rect 1740 8040 1750 8080
rect 1750 8040 1790 8080
rect 1790 8040 1800 8080
rect 1740 8030 1800 8040
rect 2070 8080 2130 8090
rect 2070 8040 2080 8080
rect 2080 8040 2120 8080
rect 2120 8040 2130 8080
rect 2070 8030 2130 8040
rect 2510 8080 2570 8090
rect 2510 8040 2520 8080
rect 2520 8040 2560 8080
rect 2560 8040 2570 8080
rect 2510 8030 2570 8040
rect 2770 8030 2830 8090
rect 3290 8080 3350 8090
rect 3290 8040 3300 8080
rect 3300 8040 3340 8080
rect 3340 8040 3350 8080
rect 3290 8030 3350 8040
rect 3970 8080 4030 8090
rect 3970 8040 3980 8080
rect 3980 8040 4020 8080
rect 4020 8040 4030 8080
rect 3970 8030 4030 8040
rect 4220 7960 4280 8020
rect 660 7190 720 7250
rect 660 7110 720 7170
rect -2630 7020 -2570 7080
rect -2860 6570 -2800 6630
rect -2970 5240 -2910 5300
rect -2970 2120 -2910 2180
rect -2860 4750 -2800 4810
rect -2740 5130 -2680 5190
rect -2740 3810 -2680 3870
rect -1240 7020 -1180 7080
rect -1020 7020 -960 7080
rect -800 7020 -740 7080
rect -580 7020 -520 7080
rect -360 7020 -300 7080
rect -140 7020 -80 7080
rect 660 7030 720 7090
rect 880 7190 940 7250
rect 880 7110 940 7170
rect 880 7030 940 7090
rect 1100 7190 1160 7250
rect 1100 7110 1160 7170
rect 1100 7030 1160 7090
rect 1320 7190 1380 7250
rect 1320 7110 1380 7170
rect 1320 7030 1380 7090
rect 1540 7190 1600 7250
rect 1540 7110 1600 7170
rect 1540 7030 1600 7090
rect 1760 7190 1820 7250
rect 1760 7110 1820 7170
rect 1760 7030 1820 7090
rect 4770 7190 4830 7250
rect 4850 7190 4910 7250
rect 4930 7190 4990 7250
rect 4770 7110 4830 7170
rect 4850 7110 4910 7170
rect 4930 7110 4990 7170
rect 4770 7030 4830 7090
rect 4850 7030 4910 7090
rect 4930 7030 4990 7090
rect -1350 6960 -1290 6970
rect -1350 6920 -1340 6960
rect -1340 6920 -1300 6960
rect -1300 6920 -1290 6960
rect -1350 6910 -1290 6920
rect -1130 6910 -1070 6970
rect -910 6910 -850 6970
rect -690 6910 -630 6970
rect -470 6910 -410 6970
rect -250 6910 -190 6970
rect -30 6960 30 6970
rect -30 6920 -20 6960
rect -20 6920 20 6960
rect 20 6920 30 6960
rect -30 6910 30 6920
rect 550 6960 610 6970
rect 550 6920 560 6960
rect 560 6920 600 6960
rect 600 6920 610 6960
rect 550 6910 610 6920
rect 770 6910 830 6970
rect 990 6910 1050 6970
rect 1210 6910 1270 6970
rect 1430 6910 1490 6970
rect 1650 6910 1710 6970
rect 1870 6960 1930 6970
rect 1870 6920 1880 6960
rect 1880 6920 1920 6960
rect 1920 6920 1930 6960
rect 1870 6910 1930 6920
rect -1182 6622 -1130 6632
rect -1182 6588 -1172 6622
rect -1172 6588 -1138 6622
rect -1138 6588 -1130 6622
rect -1182 6580 -1130 6588
rect -1072 6622 -1020 6632
rect -1072 6588 -1062 6622
rect -1062 6588 -1028 6622
rect -1028 6588 -1020 6622
rect -1072 6580 -1020 6588
rect -962 6622 -910 6632
rect -962 6588 -952 6622
rect -952 6588 -918 6622
rect -918 6588 -910 6622
rect -962 6580 -910 6588
rect -852 6622 -800 6632
rect -852 6588 -842 6622
rect -842 6588 -808 6622
rect -808 6588 -800 6622
rect -852 6580 -800 6588
rect -742 6622 -690 6632
rect -742 6588 -732 6622
rect -732 6588 -698 6622
rect -698 6588 -690 6622
rect -742 6580 -690 6588
rect -632 6622 -580 6632
rect -632 6588 -622 6622
rect -622 6588 -588 6622
rect -588 6588 -580 6622
rect -632 6580 -580 6588
rect -522 6622 -470 6632
rect -522 6588 -512 6622
rect -512 6588 -478 6622
rect -478 6588 -470 6622
rect -522 6580 -470 6588
rect -412 6622 -360 6632
rect -412 6588 -402 6622
rect -402 6588 -368 6622
rect -368 6588 -360 6622
rect -412 6580 -360 6588
rect -302 6622 -250 6632
rect -302 6588 -292 6622
rect -292 6588 -258 6622
rect -258 6588 -250 6622
rect -302 6580 -250 6588
rect -192 6622 -140 6632
rect -192 6588 -182 6622
rect -182 6588 -148 6622
rect -148 6588 -140 6622
rect -192 6580 -140 6588
rect 718 6622 770 6632
rect 718 6588 728 6622
rect 728 6588 762 6622
rect 762 6588 770 6622
rect 718 6580 770 6588
rect 828 6622 880 6632
rect 828 6588 838 6622
rect 838 6588 872 6622
rect 872 6588 880 6622
rect 828 6580 880 6588
rect 938 6622 990 6632
rect 938 6588 948 6622
rect 948 6588 982 6622
rect 982 6588 990 6622
rect 938 6580 990 6588
rect 1048 6622 1100 6632
rect 1048 6588 1058 6622
rect 1058 6588 1092 6622
rect 1092 6588 1100 6622
rect 1048 6580 1100 6588
rect 1158 6622 1210 6632
rect 1158 6588 1168 6622
rect 1168 6588 1202 6622
rect 1202 6588 1210 6622
rect 1158 6580 1210 6588
rect 1268 6622 1320 6632
rect 1268 6588 1278 6622
rect 1278 6588 1312 6622
rect 1312 6588 1320 6622
rect 1268 6580 1320 6588
rect 1378 6622 1430 6632
rect 1378 6588 1388 6622
rect 1388 6588 1422 6622
rect 1422 6588 1430 6622
rect 1378 6580 1430 6588
rect 1488 6622 1540 6632
rect 1488 6588 1498 6622
rect 1498 6588 1532 6622
rect 1532 6588 1540 6622
rect 1488 6580 1540 6588
rect 1598 6622 1650 6632
rect 1598 6588 1608 6622
rect 1608 6588 1642 6622
rect 1642 6588 1650 6622
rect 1598 6580 1650 6588
rect 1708 6622 1760 6632
rect 1708 6588 1718 6622
rect 1718 6588 1752 6622
rect 1752 6588 1760 6622
rect 1708 6580 1760 6588
rect -1360 6470 -1300 6530
rect -1360 6390 -1300 6450
rect -1360 6360 -1300 6370
rect -1360 6320 -1350 6360
rect -1350 6320 -1310 6360
rect -1310 6320 -1300 6360
rect -1360 6310 -1300 6320
rect -1000 6470 -940 6530
rect -1000 6390 -940 6450
rect -1000 6360 -940 6370
rect -1000 6320 -990 6360
rect -990 6320 -950 6360
rect -950 6320 -940 6360
rect -1000 6310 -940 6320
rect -640 6470 -580 6530
rect -640 6390 -580 6450
rect -640 6360 -580 6370
rect -640 6320 -630 6360
rect -630 6320 -590 6360
rect -590 6320 -580 6360
rect -640 6310 -580 6320
rect -280 6470 -220 6530
rect -280 6390 -220 6450
rect -280 6360 -220 6370
rect -280 6320 -270 6360
rect -270 6320 -230 6360
rect -230 6320 -220 6360
rect -280 6310 -220 6320
rect 80 6470 140 6530
rect 80 6390 140 6450
rect 80 6360 140 6370
rect 80 6320 90 6360
rect 90 6320 130 6360
rect 130 6320 140 6360
rect 80 6310 140 6320
rect 440 6470 500 6530
rect 440 6390 500 6450
rect 440 6360 500 6370
rect 440 6320 450 6360
rect 450 6320 490 6360
rect 490 6320 500 6360
rect 440 6310 500 6320
rect 800 6470 860 6530
rect 800 6390 860 6450
rect 800 6360 860 6370
rect 800 6320 810 6360
rect 810 6320 850 6360
rect 850 6320 860 6360
rect 800 6310 860 6320
rect 1160 6470 1220 6530
rect 1160 6390 1220 6450
rect 1160 6360 1220 6370
rect 1160 6320 1170 6360
rect 1170 6320 1210 6360
rect 1210 6320 1220 6360
rect 1160 6310 1220 6320
rect 1520 6470 1580 6530
rect 1520 6390 1580 6450
rect 1520 6360 1580 6370
rect 1520 6320 1530 6360
rect 1530 6320 1570 6360
rect 1570 6320 1580 6360
rect 1520 6310 1580 6320
rect 1880 6470 1940 6530
rect 1880 6390 1940 6450
rect 1880 6360 1940 6370
rect 1880 6320 1890 6360
rect 1890 6320 1930 6360
rect 1930 6320 1940 6360
rect 1880 6310 1940 6320
rect 2510 6470 2570 6530
rect 2510 6390 2570 6450
rect 2510 6310 2570 6370
rect 2950 6470 3010 6530
rect 2950 6390 3010 6450
rect 2950 6310 3010 6370
rect -1090 5620 -1030 5630
rect -1090 5580 -1080 5620
rect -1080 5580 -1040 5620
rect -1040 5580 -1030 5620
rect -1090 5570 -1030 5580
rect -910 5620 -850 5630
rect -910 5580 -900 5620
rect -900 5580 -860 5620
rect -860 5580 -850 5620
rect -910 5570 -850 5580
rect -730 5620 -670 5630
rect -730 5580 -720 5620
rect -720 5580 -680 5620
rect -680 5580 -670 5620
rect -730 5570 -670 5580
rect -550 5620 -490 5630
rect -550 5580 -540 5620
rect -540 5580 -500 5620
rect -500 5580 -490 5620
rect -550 5570 -490 5580
rect -370 5620 -310 5630
rect -370 5580 -360 5620
rect -360 5580 -320 5620
rect -320 5580 -310 5620
rect -370 5570 -310 5580
rect -190 5620 -130 5630
rect -190 5580 -180 5620
rect -180 5580 -140 5620
rect -140 5580 -130 5620
rect -190 5570 -130 5580
rect -10 5620 50 5630
rect -10 5580 0 5620
rect 0 5580 40 5620
rect 40 5580 50 5620
rect -10 5570 50 5580
rect 170 5620 230 5630
rect 170 5580 180 5620
rect 180 5580 220 5620
rect 220 5580 230 5620
rect 170 5570 230 5580
rect -100 5460 -40 5520
rect -460 5350 -400 5410
rect -820 5240 -760 5300
rect 350 5620 410 5630
rect 350 5580 360 5620
rect 360 5580 400 5620
rect 400 5580 410 5620
rect 350 5570 410 5580
rect 440 5570 500 5630
rect 530 5620 590 5630
rect 530 5580 540 5620
rect 540 5580 580 5620
rect 580 5580 590 5620
rect 530 5570 590 5580
rect -1180 5130 -1120 5190
rect 260 5130 320 5190
rect -2460 5020 -2400 5080
rect -2460 4940 -2400 5000
rect -2460 4860 -2400 4920
rect -2220 5020 -2160 5080
rect -2220 4940 -2160 5000
rect -2220 4860 -2160 4920
rect -1980 5020 -1920 5080
rect -1980 4940 -1920 5000
rect -1980 4860 -1920 4920
rect -1740 5020 -1680 5080
rect -1740 4940 -1680 5000
rect -1740 4860 -1680 4920
rect -1500 5020 -1440 5080
rect -1500 4940 -1440 5000
rect -1500 4860 -1440 4920
rect -1260 5020 -1200 5080
rect -1260 4940 -1200 5000
rect -1260 4860 -1200 4920
rect -1020 5020 -960 5080
rect -1020 4940 -960 5000
rect -1020 4860 -960 4920
rect -780 5020 -720 5080
rect -780 4940 -720 5000
rect -780 4860 -720 4920
rect -540 5020 -480 5080
rect -540 4940 -480 5000
rect -540 4860 -480 4920
rect -300 5020 -240 5080
rect -300 4940 -240 5000
rect -300 4860 -240 4920
rect -60 5020 0 5080
rect -60 4940 0 5000
rect -60 4860 0 4920
rect -2340 4750 -2280 4810
rect -2100 4460 -2040 4470
rect -2100 4420 -2090 4460
rect -2090 4420 -2050 4460
rect -2050 4420 -2040 4460
rect -2100 4410 -2040 4420
rect -1620 4750 -1560 4810
rect -1380 4460 -1320 4470
rect -1380 4420 -1370 4460
rect -1370 4420 -1330 4460
rect -1330 4420 -1320 4460
rect -1380 4410 -1320 4420
rect -2630 3580 -2570 3640
rect -2360 4290 -2300 4350
rect -2280 4290 -2220 4350
rect -1860 4290 -1800 4350
rect -1620 4290 -1560 4350
rect -1620 4020 -1560 4080
rect -900 4750 -840 4810
rect -660 4460 -600 4470
rect -660 4420 -650 4460
rect -650 4420 -610 4460
rect -610 4420 -600 4460
rect -660 4410 -600 4420
rect -180 4750 -120 4810
rect 80 4750 140 4810
rect 710 5620 770 5630
rect 710 5580 720 5620
rect 720 5580 760 5620
rect 760 5580 770 5620
rect 710 5570 770 5580
rect 890 5620 950 5630
rect 890 5580 900 5620
rect 900 5580 940 5620
rect 940 5580 950 5620
rect 890 5570 950 5580
rect 620 5460 680 5520
rect 1070 5620 1130 5630
rect 1070 5580 1080 5620
rect 1080 5580 1120 5620
rect 1120 5580 1130 5620
rect 1070 5570 1130 5580
rect 1250 5620 1310 5630
rect 1250 5580 1260 5620
rect 1260 5580 1300 5620
rect 1300 5580 1310 5620
rect 1250 5570 1310 5580
rect 980 5350 1040 5410
rect 1430 5620 1490 5630
rect 1430 5580 1440 5620
rect 1440 5580 1480 5620
rect 1480 5580 1490 5620
rect 1430 5570 1490 5580
rect 1610 5620 1670 5630
rect 1610 5580 1620 5620
rect 1620 5580 1660 5620
rect 1660 5580 1670 5620
rect 1610 5570 1670 5580
rect 1340 5240 1400 5300
rect 2260 6110 2320 6170
rect 2730 6160 2790 6170
rect 2730 6120 2740 6160
rect 2740 6120 2780 6160
rect 2780 6120 2790 6160
rect 2730 6110 2790 6120
rect 2610 5820 2670 5830
rect 2610 5780 2620 5820
rect 2620 5780 2660 5820
rect 2660 5780 2670 5820
rect 2610 5770 2670 5780
rect 2260 5350 2320 5410
rect 2850 5820 2910 5830
rect 2850 5780 2860 5820
rect 2860 5780 2900 5820
rect 2900 5780 2910 5820
rect 2850 5770 2910 5780
rect 2730 5240 2790 5300
rect 1700 5130 1760 5190
rect 580 5020 640 5080
rect 580 4940 640 5000
rect 580 4860 640 4920
rect 820 5020 880 5080
rect 820 4940 880 5000
rect 820 4860 880 4920
rect 1060 5020 1120 5080
rect 1060 4940 1120 5000
rect 1060 4860 1120 4920
rect 1300 5020 1360 5080
rect 1300 4940 1360 5000
rect 1300 4860 1360 4920
rect 1540 5020 1600 5080
rect 1540 4940 1600 5000
rect 1540 4860 1600 4920
rect 1780 5020 1840 5080
rect 1780 4940 1840 5000
rect 1780 4860 1840 4920
rect 2020 5020 2080 5080
rect 2020 4940 2080 5000
rect 2020 4860 2080 4920
rect 2260 5020 2320 5080
rect 2260 4940 2320 5000
rect 2260 4860 2320 4920
rect 2500 5020 2560 5080
rect 2500 4940 2560 5000
rect 2500 4860 2560 4920
rect 2740 5020 2800 5080
rect 2740 4940 2800 5000
rect 2740 4860 2800 4920
rect 440 4750 500 4810
rect -1140 4290 -1080 4350
rect -900 4290 -840 4350
rect -420 4290 -360 4350
rect -240 4290 -180 4350
rect -1140 4020 -1080 4080
rect -660 4020 -600 4080
rect -1380 3910 -1320 3970
rect -1454 3852 -1402 3860
rect -1454 3818 -1446 3852
rect -1446 3818 -1412 3852
rect -1412 3818 -1402 3852
rect -1454 3808 -1402 3818
rect -1296 3852 -1244 3860
rect -1296 3818 -1288 3852
rect -1288 3818 -1254 3852
rect -1254 3818 -1244 3852
rect -1296 3808 -1244 3818
rect -900 3910 -840 3970
rect -972 3852 -920 3860
rect -972 3818 -964 3852
rect -964 3818 -930 3852
rect -930 3818 -920 3852
rect -972 3808 -920 3818
rect -818 3852 -766 3860
rect -818 3818 -810 3852
rect -810 3818 -776 3852
rect -776 3818 -766 3852
rect -818 3808 -766 3818
rect -420 3910 -360 3970
rect -494 3852 -442 3860
rect -494 3818 -486 3852
rect -486 3818 -452 3852
rect -452 3818 -442 3852
rect -494 3808 -442 3818
rect -180 3810 -120 3820
rect -180 3770 -170 3810
rect -170 3770 -130 3810
rect -130 3770 -120 3810
rect -180 3760 -120 3770
rect -180 3730 -120 3740
rect -180 3690 -170 3730
rect -170 3690 -130 3730
rect -130 3690 -120 3730
rect -180 3680 -120 3690
rect -1557 3622 -1505 3632
rect -1557 3588 -1547 3622
rect -1547 3588 -1513 3622
rect -1513 3588 -1505 3622
rect -1557 3580 -1505 3588
rect -1197 3622 -1145 3632
rect -1197 3588 -1187 3622
rect -1187 3588 -1153 3622
rect -1153 3588 -1145 3622
rect -1197 3580 -1145 3588
rect -1077 3622 -1025 3632
rect -1077 3588 -1067 3622
rect -1067 3588 -1033 3622
rect -1033 3588 -1025 3622
rect -1077 3580 -1025 3588
rect -717 3622 -665 3632
rect -717 3588 -707 3622
rect -707 3588 -673 3622
rect -673 3588 -665 3622
rect -717 3580 -665 3588
rect -597 3622 -545 3632
rect -597 3588 -587 3622
rect -587 3588 -553 3622
rect -553 3588 -545 3622
rect -597 3580 -545 3588
rect -180 3650 -120 3660
rect -180 3610 -170 3650
rect -170 3610 -130 3650
rect -130 3610 -120 3650
rect -180 3600 -120 3610
rect -2240 3470 -2180 3530
rect -1490 3470 -1430 3530
rect -1270 3470 -1210 3530
rect -1010 3470 -950 3530
rect -790 3470 -730 3530
rect -530 3470 -470 3530
rect -2060 3360 -2000 3420
rect -2060 3280 -2000 3340
rect -2060 3250 -2000 3260
rect -2060 3210 -2050 3250
rect -2050 3210 -2010 3250
rect -2010 3210 -2000 3250
rect -2060 3200 -2000 3210
rect -1820 3360 -1760 3420
rect -1820 3280 -1760 3340
rect -1820 3250 -1760 3260
rect -1820 3210 -1810 3250
rect -1810 3210 -1770 3250
rect -1770 3210 -1760 3250
rect -1820 3200 -1760 3210
rect -1580 3360 -1520 3420
rect -1580 3280 -1520 3340
rect -1580 3250 -1520 3260
rect -1580 3210 -1570 3250
rect -1570 3210 -1530 3250
rect -1530 3210 -1520 3250
rect -1580 3200 -1520 3210
rect -1340 3360 -1280 3420
rect -1340 3280 -1280 3340
rect -1340 3250 -1280 3260
rect -1340 3210 -1330 3250
rect -1330 3210 -1290 3250
rect -1290 3210 -1280 3250
rect -1340 3200 -1280 3210
rect -700 3360 -640 3420
rect -700 3280 -640 3340
rect -700 3250 -640 3260
rect -700 3210 -690 3250
rect -690 3210 -650 3250
rect -650 3210 -640 3250
rect -700 3200 -640 3210
rect -460 3360 -400 3420
rect -460 3280 -400 3340
rect -460 3250 -400 3260
rect -460 3210 -450 3250
rect -450 3210 -410 3250
rect -410 3210 -400 3250
rect -460 3200 -400 3210
rect -220 3360 -160 3420
rect -220 3280 -160 3340
rect -220 3250 -160 3260
rect -220 3210 -210 3250
rect -210 3210 -170 3250
rect -170 3210 -160 3250
rect -220 3200 -160 3210
rect 180 3760 240 3820
rect 260 3760 320 3820
rect 340 3760 400 3820
rect 180 3680 240 3740
rect 260 3680 320 3740
rect 340 3680 400 3740
rect 180 3600 240 3660
rect 260 3600 320 3660
rect 340 3600 400 3660
rect -1080 2610 -1020 2620
rect -1080 2570 -1070 2610
rect -1070 2570 -1030 2610
rect -1030 2570 -1020 2610
rect -1080 2560 -1020 2570
rect -1080 2480 -1020 2540
rect -1080 2400 -1020 2460
rect 700 4750 760 4810
rect 1420 4750 1480 4810
rect 1180 4460 1240 4470
rect 1180 4420 1190 4460
rect 1190 4420 1230 4460
rect 1230 4420 1240 4460
rect 1180 4410 1240 4420
rect 2140 4750 2200 4810
rect 1900 4460 1960 4470
rect 1900 4420 1910 4460
rect 1910 4420 1950 4460
rect 1950 4420 1960 4460
rect 1900 4410 1960 4420
rect 760 4290 820 4350
rect 760 4210 820 4270
rect 760 4130 820 4190
rect 940 4290 1000 4350
rect 940 4210 1000 4270
rect 940 4130 1000 4190
rect 1180 4290 1240 4350
rect 1180 4210 1240 4270
rect 1180 4130 1240 4190
rect 1420 4290 1480 4350
rect 1420 4210 1480 4270
rect 1420 4130 1480 4190
rect 1660 4290 1720 4350
rect 1660 4210 1720 4270
rect 1660 4130 1720 4190
rect 1180 4020 1240 4080
rect 1660 4020 1720 4080
rect 940 3910 1000 3970
rect 700 3810 760 3820
rect 700 3770 710 3810
rect 710 3770 750 3810
rect 750 3770 760 3810
rect 700 3760 760 3770
rect 1022 3852 1074 3860
rect 1022 3818 1032 3852
rect 1032 3818 1066 3852
rect 1066 3818 1074 3852
rect 1022 3808 1074 3818
rect 1420 3910 1480 3970
rect 1346 3852 1398 3860
rect 1346 3818 1356 3852
rect 1356 3818 1390 3852
rect 1390 3818 1398 3852
rect 1346 3808 1398 3818
rect 1500 3852 1552 3860
rect 1500 3818 1510 3852
rect 1510 3818 1544 3852
rect 1544 3818 1552 3852
rect 1500 3808 1552 3818
rect 3170 5460 3230 5520
rect 2980 5020 3040 5080
rect 2980 4940 3040 5000
rect 2980 4860 3040 4920
rect 2860 4750 2920 4810
rect 2620 4460 2680 4470
rect 2620 4420 2630 4460
rect 2630 4420 2670 4460
rect 2670 4420 2680 4460
rect 2620 4410 2680 4420
rect 2140 4290 2200 4350
rect 2140 4210 2200 4270
rect 2140 4130 2200 4190
rect 2380 4290 2440 4350
rect 2380 4210 2440 4270
rect 2380 4130 2440 4190
rect 2800 4290 2860 4350
rect 2800 4210 2860 4270
rect 2800 4130 2860 4190
rect 2140 4020 2200 4080
rect 1900 3910 1960 3970
rect 1824 3852 1876 3860
rect 1824 3818 1834 3852
rect 1834 3818 1868 3852
rect 1868 3818 1876 3852
rect 1824 3808 1876 3818
rect 1982 3852 2034 3860
rect 1982 3818 1992 3852
rect 1992 3818 2026 3852
rect 2026 3818 2034 3852
rect 1982 3808 2034 3818
rect 700 3730 760 3740
rect 700 3690 710 3730
rect 710 3690 750 3730
rect 750 3690 760 3730
rect 700 3680 760 3690
rect 700 3650 760 3660
rect 700 3610 710 3650
rect 710 3610 750 3650
rect 750 3610 760 3650
rect 700 3600 760 3610
rect 1125 3622 1177 3632
rect 1125 3588 1133 3622
rect 1133 3588 1167 3622
rect 1167 3588 1177 3622
rect 1125 3580 1177 3588
rect 1245 3622 1297 3632
rect 1245 3588 1253 3622
rect 1253 3588 1287 3622
rect 1287 3588 1297 3622
rect 1245 3580 1297 3588
rect 1605 3622 1657 3632
rect 1605 3588 1613 3622
rect 1613 3588 1647 3622
rect 1647 3588 1657 3622
rect 1605 3580 1657 3588
rect 1725 3622 1777 3632
rect 1725 3588 1733 3622
rect 1733 3588 1767 3622
rect 1767 3588 1777 3622
rect 1725 3580 1777 3588
rect 3260 5350 3320 5410
rect 6760 9940 6820 10000
rect 6100 9290 6160 9350
rect 5260 9170 5320 9230
rect 7080 9940 7140 10000
rect 7400 9940 7460 10000
rect 7840 9940 7900 10000
rect 6540 9290 6600 9350
rect 6980 9290 7040 9350
rect 8280 9940 8340 10000
rect 6320 9170 6380 9230
rect 5900 8950 5960 9010
rect 5460 8100 5520 8160
rect 5680 8100 5740 8160
rect 6120 8100 6180 8160
rect 6440 8100 6500 8160
rect 7490 9310 7550 9320
rect 7490 9270 7500 9310
rect 7500 9270 7540 9310
rect 7540 9270 7550 9310
rect 7490 9260 7550 9270
rect 7620 9290 7680 9350
rect 8500 9940 8560 10000
rect 8060 9290 8120 9350
rect 7490 9060 7550 9120
rect 8190 9310 8250 9320
rect 8190 9270 8200 9310
rect 8200 9270 8240 9310
rect 8240 9270 8250 9310
rect 8190 9260 8250 9270
rect 8870 9270 8940 9340
rect 8060 9010 8120 9070
rect 7930 8810 7990 8820
rect 7930 8770 7940 8810
rect 7940 8770 7980 8810
rect 7980 8770 7990 8810
rect 7930 8760 7990 8770
rect 6760 8100 6820 8160
rect 7200 8100 7260 8160
rect 7520 8100 7580 8160
rect 12120 9010 12180 9070
rect 8190 8810 8250 8820
rect 8190 8770 8200 8810
rect 8200 8770 8240 8810
rect 8240 8770 8250 8810
rect 8190 8760 8250 8770
rect 8870 8740 8940 8810
rect 7840 8100 7900 8160
rect 8280 8100 8340 8160
rect 8500 8100 8560 8160
rect 9220 7950 9290 8020
rect 5260 7830 5320 7890
rect 12010 7830 12070 7890
rect 5040 5080 5100 5140
rect 5150 7720 5210 7780
rect 5150 7640 5210 7700
rect 5150 7560 5210 7620
rect 9340 7200 9400 7260
rect 9130 6730 9190 6740
rect 9130 6690 9140 6730
rect 9140 6690 9180 6730
rect 9180 6690 9190 6730
rect 9130 6680 9190 6690
rect 5150 4920 5210 4980
rect 5260 6340 5320 6350
rect 5260 6300 5270 6340
rect 5270 6300 5310 6340
rect 5310 6300 5320 6340
rect 5260 6290 5320 6300
rect 3490 4750 3550 4810
rect 3260 3810 3320 3870
rect 2085 3622 2137 3632
rect 2085 3588 2093 3622
rect 2093 3588 2127 3622
rect 2127 3588 2137 3622
rect 2085 3580 2137 3588
rect 3170 3580 3230 3640
rect 1050 3470 1110 3530
rect 1310 3470 1370 3530
rect 1530 3470 1590 3530
rect 1790 3470 1850 3530
rect 2010 3470 2070 3530
rect 2760 3470 2820 3530
rect 740 3360 800 3420
rect 740 3280 800 3340
rect 740 3250 800 3260
rect 740 3210 750 3250
rect 750 3210 790 3250
rect 790 3210 800 3250
rect 740 3200 800 3210
rect 980 3360 1040 3420
rect 980 3280 1040 3340
rect 980 3250 1040 3260
rect 980 3210 990 3250
rect 990 3210 1030 3250
rect 1030 3210 1040 3250
rect 980 3200 1040 3210
rect 1220 3360 1280 3420
rect 1220 3280 1280 3340
rect 1220 3250 1280 3260
rect 1220 3210 1230 3250
rect 1230 3210 1270 3250
rect 1270 3210 1280 3250
rect 1220 3200 1280 3210
rect 1860 3360 1920 3420
rect 1860 3280 1920 3340
rect 1860 3250 1920 3260
rect 1860 3210 1870 3250
rect 1870 3210 1910 3250
rect 1910 3210 1920 3250
rect 1860 3200 1920 3210
rect 2100 3360 2160 3420
rect 2100 3280 2160 3340
rect 2100 3250 2160 3260
rect 2100 3210 2110 3250
rect 2110 3210 2150 3250
rect 2150 3210 2160 3250
rect 2100 3200 2160 3210
rect 2340 3360 2400 3420
rect 2340 3280 2400 3340
rect 2340 3250 2400 3260
rect 2340 3210 2350 3250
rect 2350 3210 2390 3250
rect 2390 3210 2400 3250
rect 2340 3200 2400 3210
rect 2580 3360 2640 3420
rect 2580 3280 2640 3340
rect 2580 3250 2640 3260
rect 2580 3210 2590 3250
rect 2590 3210 2630 3250
rect 2630 3210 2640 3250
rect 2580 3200 2640 3210
rect 180 2560 240 2620
rect 260 2560 320 2620
rect 340 2560 400 2620
rect 180 2480 240 2540
rect 260 2480 320 2540
rect 340 2480 400 2540
rect 180 2400 240 2460
rect 260 2400 320 2460
rect 340 2400 400 2460
rect 1600 2610 1660 2620
rect 1600 2570 1610 2610
rect 1610 2570 1650 2610
rect 1650 2570 1660 2610
rect 1600 2560 1660 2570
rect 1600 2480 1660 2540
rect 1600 2400 1660 2460
rect -1820 2340 -1760 2350
rect -1820 2300 -1810 2340
rect -1810 2300 -1770 2340
rect -1770 2300 -1760 2340
rect -1820 2290 -1760 2300
rect -1660 2340 -1600 2350
rect -1660 2300 -1650 2340
rect -1650 2300 -1610 2340
rect -1610 2300 -1600 2340
rect -1660 2290 -1600 2300
rect -1500 2340 -1440 2350
rect -1500 2300 -1490 2340
rect -1490 2300 -1450 2340
rect -1450 2300 -1440 2340
rect -1500 2290 -1440 2300
rect -1340 2340 -1280 2350
rect -1340 2300 -1330 2340
rect -1330 2300 -1290 2340
rect -1290 2300 -1280 2340
rect -1340 2290 -1280 2300
rect -1180 2340 -1120 2350
rect -1180 2300 -1170 2340
rect -1170 2300 -1130 2340
rect -1130 2300 -1120 2340
rect -1180 2290 -1120 2300
rect -1020 2340 -960 2350
rect -1020 2300 -1010 2340
rect -1010 2300 -970 2340
rect -970 2300 -960 2340
rect -1020 2290 -960 2300
rect -860 2340 -800 2350
rect -860 2300 -850 2340
rect -850 2300 -810 2340
rect -810 2300 -800 2340
rect -860 2290 -800 2300
rect -700 2340 -640 2350
rect -700 2300 -690 2340
rect -690 2300 -650 2340
rect -650 2300 -640 2340
rect -700 2290 -640 2300
rect -540 2340 -480 2350
rect -540 2300 -530 2340
rect -530 2300 -490 2340
rect -490 2300 -480 2340
rect -540 2290 -480 2300
rect -380 2340 -320 2350
rect -380 2300 -370 2340
rect -370 2300 -330 2340
rect -330 2300 -320 2340
rect -380 2290 -320 2300
rect -220 2340 -160 2350
rect -220 2300 -210 2340
rect -210 2300 -170 2340
rect -170 2300 -160 2340
rect -220 2290 -160 2300
rect -60 2340 0 2350
rect -60 2300 -50 2340
rect -50 2300 -10 2340
rect -10 2300 0 2340
rect -60 2290 0 2300
rect 100 2340 160 2350
rect 100 2300 110 2340
rect 110 2300 150 2340
rect 150 2300 160 2340
rect 100 2290 160 2300
rect 260 2340 320 2350
rect 260 2300 270 2340
rect 270 2300 310 2340
rect 310 2300 320 2340
rect 260 2290 320 2300
rect 420 2340 480 2350
rect 420 2300 430 2340
rect 430 2300 470 2340
rect 470 2300 480 2340
rect 420 2290 480 2300
rect 580 2340 640 2350
rect 580 2300 590 2340
rect 590 2300 630 2340
rect 630 2300 640 2340
rect 580 2290 640 2300
rect 740 2340 800 2350
rect 740 2300 750 2340
rect 750 2300 790 2340
rect 790 2300 800 2340
rect 740 2290 800 2300
rect 900 2340 960 2350
rect 900 2300 910 2340
rect 910 2300 950 2340
rect 950 2300 960 2340
rect 900 2290 960 2300
rect 1060 2340 1120 2350
rect 1060 2300 1070 2340
rect 1070 2300 1110 2340
rect 1110 2300 1120 2340
rect 1060 2290 1120 2300
rect 1220 2340 1280 2350
rect 1220 2300 1230 2340
rect 1230 2300 1270 2340
rect 1270 2300 1280 2340
rect 1220 2290 1280 2300
rect 1380 2340 1440 2350
rect 1380 2300 1390 2340
rect 1390 2300 1430 2340
rect 1430 2300 1440 2340
rect 1380 2290 1440 2300
rect 1540 2340 1600 2350
rect 1540 2300 1550 2340
rect 1550 2300 1590 2340
rect 1590 2300 1600 2340
rect 1540 2290 1600 2300
rect 1700 2340 1760 2350
rect 1700 2300 1710 2340
rect 1710 2300 1750 2340
rect 1750 2300 1760 2340
rect 1700 2290 1760 2300
rect 1860 2340 1920 2350
rect 1860 2300 1870 2340
rect 1870 2300 1910 2340
rect 1910 2300 1920 2340
rect 1860 2290 1920 2300
rect 2020 2340 2080 2350
rect 2020 2300 2030 2340
rect 2030 2300 2070 2340
rect 2070 2300 2080 2340
rect 2020 2290 2080 2300
rect 2180 2340 2240 2350
rect 2180 2300 2190 2340
rect 2190 2300 2230 2340
rect 2230 2300 2240 2340
rect 2180 2290 2240 2300
rect -1900 2170 -1840 2180
rect -1900 2130 -1890 2170
rect -1890 2130 -1850 2170
rect -1850 2130 -1840 2170
rect -1900 2120 -1840 2130
rect 2490 2210 2550 2220
rect 2490 2170 2500 2210
rect 2500 2170 2540 2210
rect 2540 2170 2550 2210
rect 2490 2160 2550 2170
rect 2490 2130 2550 2140
rect 2490 2090 2500 2130
rect 2500 2090 2540 2130
rect 2540 2090 2550 2130
rect 2490 2080 2550 2090
rect -2360 1950 -2300 2010
rect -1950 1950 -1890 2010
rect -2630 1840 -2570 1900
rect -2310 1610 -2250 1670
rect -2310 -20 -2240 -10
rect -2310 -70 -2300 -20
rect -2300 -70 -2250 -20
rect -2250 -70 -2240 -20
rect -2310 -80 -2240 -70
rect -2860 -450 -2790 -440
rect -2860 -500 -2850 -450
rect -2850 -500 -2800 -450
rect -2800 -500 -2790 -450
rect -2740 -400 -2670 -390
rect -2740 -450 -2730 -400
rect -2730 -450 -2680 -400
rect -2680 -450 -2670 -400
rect -2740 -460 -2670 -450
rect -2860 -510 -2790 -500
rect -2860 -1798 -2790 -1788
rect -2860 -1848 -2850 -1798
rect -2850 -1848 -2800 -1798
rect -2800 -1848 -2790 -1798
rect -2860 -1858 -2790 -1848
rect -3030 -2590 -2970 -2530
rect -3030 -2670 -2970 -2610
rect -3030 -2750 -2970 -2690
rect -2500 -2008 -2430 -1998
rect -2500 -2058 -2490 -2008
rect -2490 -2058 -2440 -2008
rect -2440 -2058 -2430 -2008
rect -2500 -2068 -2430 -2058
rect -2490 -2590 -2430 -2530
rect -2490 -2670 -2430 -2610
rect -2490 -2750 -2430 -2690
rect -2070 -2158 -2000 -2148
rect -2070 -2208 -2060 -2158
rect -2060 -2208 -2010 -2158
rect -2010 -2208 -2000 -2158
rect -2070 -2218 -2000 -2208
rect -2060 -2590 -2000 -2530
rect -2060 -2670 -2000 -2610
rect -2060 -2750 -2000 -2690
rect -2860 -2860 -2800 -2800
rect 2830 1840 2890 1900
rect -1840 1720 -1780 1780
rect -438 1780 -368 1790
rect -438 1730 -428 1780
rect -428 1730 -378 1780
rect -378 1730 -368 1780
rect -438 1720 -368 1730
rect 960 1780 1030 1790
rect 960 1730 970 1780
rect 970 1730 1020 1780
rect 1020 1730 1030 1780
rect 960 1720 1030 1730
rect 970 1610 1030 1670
rect 2360 1530 2420 1590
rect 2710 1530 2770 1590
rect -1840 -480 -1780 -420
rect -1410 -480 -1350 -420
rect 260 -424 264 -420
rect 264 -424 320 -420
rect 260 -480 320 -424
rect 2700 -20 2770 -10
rect 2700 -70 2710 -20
rect 2710 -70 2760 -20
rect 2760 -70 2770 -20
rect 2700 -80 2770 -70
rect 2360 -480 2420 -420
rect 3170 1730 3230 1790
rect 3260 1530 3320 1590
rect 3600 4290 3660 4350
rect 3680 4290 3740 4350
rect 3760 4290 3820 4350
rect 3600 4210 3660 4270
rect 3680 4210 3740 4270
rect 3760 4210 3820 4270
rect 3600 4130 3660 4190
rect 3680 4130 3740 4190
rect 3760 4130 3820 4190
rect 5520 5560 5580 5620
rect 5720 5560 5780 5620
rect 5960 5610 6020 5620
rect 5960 5570 5970 5610
rect 5970 5570 6010 5610
rect 6010 5570 6020 5610
rect 5960 5560 6020 5570
rect 6120 5560 6180 5620
rect 6520 5560 6580 5620
rect 6920 5560 6980 5620
rect 7100 5720 7160 5730
rect 7100 5680 7110 5720
rect 7110 5680 7150 5720
rect 7150 5680 7160 5720
rect 7100 5670 7160 5680
rect 7320 5560 7380 5620
rect 7520 5560 7580 5620
rect 8240 5610 8300 5620
rect 8240 5570 8250 5610
rect 8250 5570 8290 5610
rect 8290 5570 8300 5610
rect 8240 5560 8300 5570
rect 7100 5500 7160 5510
rect 7100 5460 7110 5500
rect 7110 5460 7150 5500
rect 7150 5460 7160 5500
rect 7100 5450 7160 5460
rect 5740 4880 5800 4890
rect 5740 4840 5750 4880
rect 5750 4840 5790 4880
rect 5790 4840 5800 4880
rect 5740 4830 5800 4840
rect 6880 5220 6940 5230
rect 6880 5180 6890 5220
rect 6890 5180 6930 5220
rect 6930 5180 6940 5220
rect 6880 5170 6940 5180
rect 6180 5100 6240 5160
rect 6090 5000 6150 5060
rect 6840 4920 6900 4980
rect 7320 5220 7380 5230
rect 7320 5180 7330 5220
rect 7330 5180 7370 5220
rect 7370 5180 7380 5220
rect 7320 5170 7380 5180
rect 8860 5220 8920 5230
rect 8860 5180 8870 5220
rect 8870 5180 8910 5220
rect 8910 5180 8920 5220
rect 8860 5170 8920 5180
rect 9570 5260 9640 5330
rect 9340 5170 9400 5230
rect 8020 5100 8080 5110
rect 8020 5060 8030 5100
rect 8030 5060 8070 5100
rect 8070 5060 8080 5100
rect 8020 5050 8080 5060
rect 9730 5050 9790 5060
rect 9730 5010 9740 5050
rect 9740 5010 9780 5050
rect 9780 5010 9790 5050
rect 9730 5000 9790 5010
rect 12120 7720 12180 7780
rect 12120 7640 12180 7700
rect 12120 7560 12180 7620
rect 6180 4880 6240 4890
rect 6180 4840 6190 4880
rect 6190 4840 6230 4880
rect 6230 4840 6240 4880
rect 6180 4830 6240 4840
rect 7250 4850 7310 4910
rect 8020 4880 8080 4890
rect 8020 4840 8030 4880
rect 8030 4840 8070 4880
rect 8070 4840 8080 4880
rect 8020 4830 8080 4840
rect 8860 4880 8920 4890
rect 8860 4840 8870 4880
rect 8870 4840 8910 4880
rect 8910 4840 8920 4880
rect 8860 4830 8920 4840
rect 9340 4830 9400 4890
rect 6040 4500 6100 4510
rect 6040 4460 6050 4500
rect 6050 4460 6090 4500
rect 6090 4460 6100 4500
rect 6040 4450 6100 4460
rect 5640 4340 5700 4400
rect 5840 4340 5900 4400
rect 6040 4200 6100 4260
rect 6240 4340 6300 4400
rect 6640 4340 6700 4400
rect 5260 3540 5320 3600
rect 7040 4340 7100 4400
rect 7120 4390 7180 4400
rect 7120 4350 7130 4390
rect 7130 4350 7170 4390
rect 7170 4350 7180 4390
rect 7120 4340 7180 4350
rect 7440 4340 7500 4400
rect 6440 3590 6500 3600
rect 6440 3550 6450 3590
rect 6450 3550 6490 3590
rect 6490 3550 6500 3590
rect 6440 3540 6500 3550
rect 7240 4200 7300 4260
rect 7640 4340 7700 4400
rect 8240 4390 8300 4400
rect 8240 4350 8250 4390
rect 8250 4350 8290 4390
rect 8290 4350 8300 4390
rect 8240 4340 8300 4350
rect 9570 4750 9640 4820
rect 6840 3590 6900 3600
rect 6840 3550 6850 3590
rect 6850 3550 6890 3590
rect 6890 3550 6900 3590
rect 6840 3540 6900 3550
rect 9130 3200 9190 3210
rect 9130 3160 9140 3200
rect 9140 3160 9180 3200
rect 9180 3160 9190 3200
rect 9130 3150 9190 3160
rect 4190 2910 4250 2970
rect 4290 2910 4350 2970
rect 3600 980 3660 1040
rect 3680 980 3740 1040
rect 3760 980 3820 1040
rect 3990 1950 4050 2010
rect 3490 -420 3550 -360
rect 3870 280 3930 340
rect 3480 -662 3550 -652
rect 3480 -712 3490 -662
rect 3490 -712 3540 -662
rect 3540 -712 3550 -662
rect 3480 -722 3550 -712
rect 2820 -870 2890 -860
rect 2820 -920 2830 -870
rect 2830 -920 2880 -870
rect 2880 -920 2890 -870
rect 2820 -930 2890 -920
rect 2820 -2008 2890 -1998
rect 2820 -2058 2830 -2008
rect 2830 -2058 2880 -2008
rect 2880 -2058 2890 -2008
rect 2820 -2068 2890 -2058
rect 2460 -2158 2530 -2148
rect 2460 -2208 2470 -2158
rect 2470 -2208 2520 -2158
rect 2520 -2208 2530 -2158
rect 2460 -2218 2530 -2208
rect 260 -2540 320 -2530
rect 260 -2580 270 -2540
rect 270 -2580 310 -2540
rect 310 -2580 320 -2540
rect 260 -2590 320 -2580
rect 260 -2620 320 -2610
rect 260 -2660 270 -2620
rect 270 -2660 310 -2620
rect 310 -2660 320 -2620
rect 260 -2670 320 -2660
rect 260 -2700 320 -2690
rect 260 -2740 270 -2700
rect 270 -2740 310 -2700
rect 310 -2740 320 -2700
rect 260 -2750 320 -2740
rect 2460 -2590 2520 -2530
rect 2460 -2670 2520 -2610
rect 2460 -2750 2520 -2690
rect 2820 -2590 2880 -2530
rect 2820 -2670 2880 -2610
rect 2820 -2750 2880 -2690
rect 4110 980 4170 1040
rect 4110 -420 4170 -360
rect 9340 2820 9400 2880
rect 4240 -1120 4300 -1060
rect 3990 -1820 4050 -1760
rect 3480 -2008 3550 -1998
rect 3480 -2058 3490 -2008
rect 3490 -2058 3540 -2008
rect 3540 -2058 3550 -2008
rect 3480 -2068 3550 -2058
rect 3860 -2070 3930 -2000
rect 3000 -2590 3060 -2530
rect 3000 -2670 3060 -2610
rect 3000 -2750 3060 -2690
rect 4310 -2520 4370 -2460
rect 4310 -2860 4370 -2800
rect 2900 -2920 2960 -2910
rect 2900 -2960 2910 -2920
rect 2910 -2960 2950 -2920
rect 2950 -2960 2960 -2920
rect 2900 -2970 2960 -2960
rect 5350 -2920 5410 -2910
rect 5350 -2960 5360 -2920
rect 5360 -2960 5400 -2920
rect 5400 -2960 5410 -2920
rect 5350 -2970 5410 -2960
rect 12120 -2970 12180 -2910
<< metal2 >>
rect 8700 14320 8800 14360
rect 8700 14260 8720 14320
rect 8780 14280 8800 14320
rect 8780 14270 11020 14280
rect 8780 14260 9420 14270
rect 8700 14220 9420 14260
rect 8700 14160 8720 14220
rect 8780 14210 9420 14220
rect 9480 14210 9940 14270
rect 10000 14210 10460 14270
rect 10520 14210 10950 14270
rect 11010 14210 11020 14270
rect 8780 14200 11020 14210
rect 8780 14160 8800 14200
rect 8700 14120 8800 14160
rect 8920 14160 11510 14170
rect 8920 14100 8930 14160
rect 8990 14100 9010 14160
rect 9070 14100 9090 14160
rect 9150 14100 11280 14160
rect 11340 14100 11360 14160
rect 11420 14100 11440 14160
rect 11500 14100 11510 14160
rect 8920 14080 11510 14100
rect 8920 14020 8930 14080
rect 8990 14020 9010 14080
rect 9070 14020 9090 14080
rect 9150 14020 11280 14080
rect 11340 14020 11360 14080
rect 11420 14020 11440 14080
rect 11500 14020 11510 14080
rect 8920 14000 11510 14020
rect 8920 13940 8930 14000
rect 8990 13940 9010 14000
rect 9070 13940 9090 14000
rect 9150 13940 11280 14000
rect 11340 13940 11360 14000
rect 11420 13940 11440 14000
rect 11500 13940 11510 14000
rect 8920 13930 11510 13940
rect 9365 13552 12190 13560
rect 9365 13500 9370 13552
rect 9422 13500 9890 13552
rect 9942 13500 10410 13552
rect 10462 13500 10976 13552
rect 11028 13550 12190 13552
rect 11028 13500 12120 13550
rect 9365 13490 12120 13500
rect 12180 13490 12190 13550
rect 9420 13390 9700 13400
rect 9480 13330 9630 13390
rect 9690 13330 9700 13390
rect 9420 13290 9700 13330
rect 9480 13230 9630 13290
rect 9690 13230 9700 13290
rect 9420 13220 9700 13230
rect 9940 13390 10220 13400
rect 10000 13330 10150 13390
rect 10210 13330 10220 13390
rect 9940 13290 10220 13330
rect 10000 13230 10150 13290
rect 10210 13230 10220 13290
rect 9940 13220 10220 13230
rect 10460 13390 10740 13400
rect 10520 13330 10670 13390
rect 10730 13330 10740 13390
rect 10460 13290 10740 13330
rect 10520 13230 10670 13290
rect 10730 13230 10740 13290
rect 10460 13220 10740 13230
rect 9380 13172 9590 13180
rect -1670 13100 -1570 13140
rect 9380 13120 9384 13172
rect 9436 13170 9590 13172
rect 9436 13120 9520 13170
rect 9380 13110 9520 13120
rect 9580 13110 9590 13170
rect 9900 13172 10110 13180
rect 9900 13120 9904 13172
rect 9956 13170 10110 13172
rect 9956 13120 10040 13170
rect 9900 13110 10040 13120
rect 10100 13110 10110 13170
rect 10420 13172 10630 13180
rect 10420 13120 10424 13172
rect 10476 13170 10630 13172
rect 10476 13120 10560 13170
rect 10420 13110 10560 13120
rect 10620 13110 10630 13170
rect 9510 13100 9590 13110
rect 10030 13100 10110 13110
rect 10550 13100 10630 13110
rect -1670 13040 -1650 13100
rect -1590 13060 -1570 13100
rect -1590 13050 8730 13060
rect -1590 13040 -1340 13050
rect -1670 13000 -1340 13040
rect -1670 12940 -1650 13000
rect -1590 12990 -1340 13000
rect -1280 12990 -1120 13050
rect -1060 12990 -650 13050
rect -590 12990 -310 13050
rect -250 12990 -90 13050
rect -30 12990 350 13050
rect 410 12990 1030 13050
rect 1090 12990 1250 13050
rect 1310 12990 1720 13050
rect 1780 12990 2180 13050
rect 2240 12990 2530 13050
rect 2590 12990 2780 13050
rect 2840 12990 3000 13050
rect 3060 12990 3330 13050
rect 3390 12990 3990 13050
rect 4050 12990 4210 13050
rect 4270 12990 4780 13050
rect 4840 12990 5040 13050
rect 5100 12990 5290 13050
rect 5350 12990 5510 13050
rect 5570 12990 6060 13050
rect 6120 12990 6340 13050
rect 6400 12990 6590 13050
rect 6650 12990 6810 13050
rect 6870 12990 7360 13050
rect 7420 12990 7640 13050
rect 7700 12990 7890 13050
rect 7950 12990 8110 13050
rect 8170 12990 8660 13050
rect 8720 12990 8730 13050
rect -1590 12980 8730 12990
rect -1590 12940 -1570 12980
rect -1670 12900 -1570 12940
rect 8920 12760 9410 12770
rect 8920 12700 8930 12760
rect 8990 12700 9010 12760
rect 9070 12700 9090 12760
rect 9150 12700 9350 12760
rect 8920 12690 9410 12700
rect 8862 12680 9410 12690
rect -1780 12670 -1490 12680
rect -1780 12610 -1770 12670
rect -1710 12610 -1560 12670
rect -1500 12610 -1490 12670
rect 8862 12672 8930 12680
rect 8862 12620 8866 12672
rect 8918 12620 8930 12672
rect 8990 12620 9010 12680
rect 9070 12620 9090 12680
rect 9150 12620 9350 12680
rect 8862 12610 9410 12620
rect -1780 12600 -1490 12610
rect 8920 12600 9410 12610
rect 8920 12540 8930 12600
rect 8990 12540 9010 12600
rect 9070 12540 9090 12600
rect 9150 12540 9350 12600
rect 8920 12530 9410 12540
rect 9440 12760 9930 12770
rect 9500 12700 9870 12760
rect 9440 12680 9930 12700
rect 9500 12620 9870 12680
rect 9440 12600 9930 12620
rect 9500 12540 9870 12600
rect 9440 12530 9930 12540
rect 9960 12760 10450 12770
rect 10020 12700 10390 12760
rect 9960 12680 10450 12700
rect 10020 12620 10390 12680
rect 9960 12600 10450 12620
rect 10020 12540 10390 12600
rect 9960 12530 10450 12540
rect 10480 12760 11510 12770
rect 10540 12700 11280 12760
rect 11340 12700 11360 12760
rect 11420 12700 11440 12760
rect 11500 12700 11510 12760
rect 10480 12680 11510 12700
rect 10540 12620 11280 12680
rect 11340 12620 11360 12680
rect 11420 12620 11440 12680
rect 11500 12620 11510 12680
rect 10480 12600 11510 12620
rect 10540 12540 11280 12600
rect 11340 12540 11360 12600
rect 11420 12540 11440 12600
rect 11500 12540 11510 12600
rect 10480 12530 11510 12540
rect -1670 12320 -1570 12360
rect -1670 12260 -1650 12320
rect -1590 12280 -1570 12320
rect -1590 12270 8730 12280
rect -1590 12260 -1180 12270
rect -1670 12220 -1180 12260
rect -1670 12160 -1650 12220
rect -1590 12210 -1180 12220
rect -1120 12210 -760 12270
rect -700 12210 -90 12270
rect -30 12210 480 12270
rect 540 12210 1190 12270
rect 1250 12210 1620 12270
rect 1680 12210 2060 12270
rect 2120 12210 2310 12270
rect 2370 12210 2530 12270
rect 2590 12210 3000 12270
rect 3060 12210 3440 12270
rect 3500 12210 4060 12270
rect 4120 12210 4400 12270
rect 4460 12210 4760 12270
rect 4820 12210 5360 12270
rect 5420 12210 5700 12270
rect 5760 12210 6060 12270
rect 6120 12210 6660 12270
rect 6720 12210 7000 12270
rect 7060 12210 7360 12270
rect 7420 12210 7960 12270
rect 8020 12210 8300 12270
rect 8360 12210 8660 12270
rect 8720 12210 8730 12270
rect -1590 12200 8730 12210
rect -1590 12160 -1570 12200
rect -1670 12120 -1570 12160
rect 9620 12090 9700 12100
rect 10140 12090 10220 12100
rect 10660 12090 10740 12100
rect 9380 12082 9630 12090
rect 9380 12030 9384 12082
rect 9436 12030 9630 12082
rect 9690 12030 9700 12090
rect 9380 12020 9700 12030
rect 9900 12082 10150 12090
rect 9900 12030 9904 12082
rect 9956 12030 10150 12082
rect 10210 12030 10220 12090
rect 9900 12020 10220 12030
rect 10420 12082 10670 12090
rect 10420 12030 10424 12082
rect 10476 12030 10670 12082
rect 10730 12030 10740 12090
rect 10420 12020 10740 12030
rect 9420 11970 9590 11980
rect 9480 11910 9520 11970
rect 9580 11910 9590 11970
rect 9420 11900 9590 11910
rect 9940 11970 10110 11980
rect 10000 11910 10040 11970
rect 10100 11910 10110 11970
rect 9940 11900 10110 11910
rect 10460 11970 10630 11980
rect 10520 11910 10560 11970
rect 10620 11910 10630 11970
rect 10460 11900 10630 11910
rect 9410 11580 9760 11590
rect 9410 11520 9420 11580
rect 9480 11520 9690 11580
rect 9750 11520 9760 11580
rect 9410 11510 9760 11520
rect 9930 11580 10280 11590
rect 9930 11520 9940 11580
rect 10000 11520 10210 11580
rect 10270 11520 10280 11580
rect 9930 11510 10280 11520
rect 10450 11580 10800 11590
rect 10450 11520 10460 11580
rect 10520 11520 10730 11580
rect 10790 11520 10800 11580
rect 10450 11510 10800 11520
rect 9490 11400 11120 11410
rect 9490 11340 9500 11400
rect 9560 11340 10020 11400
rect 10080 11340 10540 11400
rect 10600 11340 10870 11400
rect 10930 11340 11060 11400
rect 9490 11330 11120 11340
rect 8700 10800 8800 10840
rect 8700 10740 8720 10800
rect 8780 10760 8800 10800
rect 8780 10750 11320 10760
rect 8780 10740 9690 10750
rect 8700 10700 9690 10740
rect 8700 10640 8720 10700
rect 8780 10690 9690 10700
rect 9750 10690 10210 10750
rect 10270 10690 10730 10750
rect 10790 10690 11250 10750
rect 11310 10690 11320 10750
rect 8780 10680 11320 10690
rect 8780 10640 8800 10680
rect 8700 10600 8800 10640
rect -980 10500 -880 10540
rect 9090 10520 9200 10540
rect -980 10440 -960 10500
rect -900 10460 -880 10500
rect 3800 10510 9110 10520
rect -900 10450 3360 10460
rect -900 10440 -630 10450
rect -980 10400 -630 10440
rect -980 10340 -960 10400
rect -900 10390 -630 10400
rect -570 10390 -410 10450
rect -350 10390 -110 10450
rect -50 10390 110 10450
rect 170 10390 270 10450
rect 330 10390 490 10450
rect 550 10390 790 10450
rect 850 10390 1010 10450
rect 1070 10390 1310 10450
rect 1370 10390 1750 10450
rect 1810 10390 2080 10450
rect 2140 10390 2510 10450
rect 2570 10390 2900 10450
rect 2960 10390 3290 10450
rect 3350 10390 3360 10450
rect 3800 10450 3810 10510
rect 3870 10450 9110 10510
rect 9180 10450 9200 10520
rect 3800 10440 9200 10450
rect 9090 10430 9200 10440
rect -900 10380 3360 10390
rect -900 10340 -880 10380
rect -980 10300 -880 10340
rect -230 10340 -150 10350
rect -230 10280 -220 10340
rect -160 10310 -150 10340
rect 1490 10340 1570 10350
rect 1490 10310 1500 10340
rect -160 10280 1500 10310
rect 1560 10310 1570 10340
rect 3570 10340 4590 10350
rect 2340 10320 2420 10330
rect 2340 10310 2350 10320
rect 1560 10280 2350 10310
rect -230 10270 2350 10280
rect 2340 10260 2350 10270
rect 2410 10260 2420 10320
rect 3570 10280 3580 10340
rect 3640 10280 4520 10340
rect 4580 10280 4590 10340
rect 3570 10270 4590 10280
rect 2340 10250 2420 10260
rect 4110 10000 4480 10010
rect 1140 9990 1220 10000
rect -1890 9960 -680 9970
rect -1890 9900 -750 9960
rect -690 9900 -680 9960
rect 1140 9930 1150 9990
rect 1210 9930 1220 9990
rect 1140 9920 1220 9930
rect 2230 9950 2310 9960
rect -1890 9890 -680 9900
rect 2230 9890 2240 9950
rect 2300 9890 2310 9950
rect 4110 9940 4120 10000
rect 4180 9940 4410 10000
rect 4470 9940 4480 10000
rect 4110 9930 4480 9940
rect 5350 10000 8570 10010
rect 5350 9940 5390 10000
rect 5450 9940 5490 10000
rect 5550 9940 5660 10000
rect 5720 9940 5880 10000
rect 5940 9940 6320 10000
rect 6380 9940 6760 10000
rect 6820 9940 7080 10000
rect 7140 9940 7400 10000
rect 7460 9940 7840 10000
rect 7900 9940 8280 10000
rect 8340 9940 8500 10000
rect 8560 9940 8570 10000
rect 5350 9930 8570 9940
rect 2230 9880 2310 9890
rect 3800 9920 3880 9930
rect 3800 9860 3810 9920
rect 3870 9860 3880 9920
rect 3800 9850 3880 9860
rect 1360 9380 1440 9390
rect -980 9320 -880 9360
rect 1360 9320 1370 9380
rect 1430 9320 1440 9380
rect 5030 9350 7050 9360
rect -980 9260 -960 9320
rect -900 9280 -880 9320
rect 5030 9290 5040 9350
rect 5100 9290 6100 9350
rect 6160 9290 6540 9350
rect 6600 9290 6980 9350
rect 7040 9290 7050 9350
rect 7610 9350 8130 9360
rect 5030 9280 7050 9290
rect 7480 9320 7560 9330
rect -900 9270 4040 9280
rect -900 9260 -630 9270
rect -980 9220 -630 9260
rect -980 9160 -960 9220
rect -900 9210 -630 9220
rect -570 9210 110 9270
rect 170 9210 270 9270
rect 330 9210 1010 9270
rect 1070 9210 1260 9270
rect 1320 9210 1450 9270
rect 1510 9210 1530 9270
rect 1590 9210 1740 9270
rect 1800 9210 2070 9270
rect 2130 9210 2510 9270
rect 2570 9210 2900 9270
rect 2960 9210 3110 9270
rect 3170 9210 3290 9270
rect 3350 9210 3970 9270
rect 4030 9210 4040 9270
rect 7480 9260 7490 9320
rect 7550 9260 7560 9320
rect 7610 9290 7620 9350
rect 7680 9290 8060 9350
rect 8120 9290 8130 9350
rect 8850 9340 8960 9360
rect 8850 9330 8870 9340
rect 7610 9280 8130 9290
rect 8180 9320 8870 9330
rect 7480 9250 7560 9260
rect 8180 9260 8190 9320
rect 8250 9270 8870 9320
rect 8940 9270 8960 9340
rect 8250 9260 8960 9270
rect 8180 9250 8960 9260
rect -900 9200 4040 9210
rect 4510 9230 6390 9240
rect -900 9160 -880 9200
rect 4510 9170 4520 9230
rect 4580 9170 5260 9230
rect 5320 9170 6320 9230
rect 6380 9170 6390 9230
rect -980 9120 -880 9160
rect -190 9160 -110 9170
rect -190 9100 -180 9160
rect -120 9150 -110 9160
rect 1340 9160 1420 9170
rect 3570 9160 4370 9170
rect 4510 9160 6390 9170
rect 1340 9150 1350 9160
rect -120 9110 1350 9150
rect -120 9100 -110 9110
rect -190 9090 -110 9100
rect 1340 9100 1350 9110
rect 1410 9140 1420 9160
rect 2340 9150 2420 9160
rect 2340 9140 2350 9150
rect 1410 9100 2350 9140
rect 1340 9090 1420 9100
rect 2340 9090 2350 9100
rect 2410 9090 2420 9150
rect 2760 9100 2770 9160
rect 2830 9150 2840 9160
rect 2930 9150 2940 9160
rect 2830 9110 2940 9150
rect 2830 9100 2840 9110
rect 2930 9100 2940 9110
rect 3000 9100 3010 9160
rect 2930 9090 3010 9100
rect 3570 9100 3580 9160
rect 3640 9100 4300 9160
rect 4360 9100 4370 9160
rect 3570 9090 4370 9100
rect 4400 9120 7560 9130
rect 2340 9080 2420 9090
rect 4400 9060 4410 9120
rect 4470 9060 7490 9120
rect 7550 9060 7560 9120
rect 4400 9050 7560 9060
rect 8050 9070 12190 9080
rect 4290 9010 5970 9020
rect 4290 8950 4300 9010
rect 4360 8950 4770 9010
rect 4830 8950 4850 9010
rect 4910 8950 4930 9010
rect 4990 8950 5900 9010
rect 5960 8950 5970 9010
rect 8050 9010 8060 9070
rect 8120 9010 12120 9070
rect 12180 9010 12190 9070
rect 8050 9000 12190 9010
rect 4290 8940 5970 8950
rect 4290 8900 8000 8910
rect 4290 8840 4300 8900
rect 4360 8840 8000 8900
rect 4290 8830 8000 8840
rect 7920 8820 8000 8830
rect 7920 8760 7930 8820
rect 7990 8760 8000 8820
rect 7920 8750 8000 8760
rect 8180 8820 8960 8830
rect 8180 8760 8190 8820
rect 8250 8810 8960 8820
rect 8250 8760 8870 8810
rect 8180 8750 8870 8760
rect 8850 8740 8870 8750
rect 8940 8740 8960 8810
rect 8850 8720 8960 8740
rect 1160 8590 1240 8600
rect -1780 8580 -680 8590
rect -1780 8520 -1770 8580
rect -1710 8520 -750 8580
rect -690 8520 -680 8580
rect 1160 8530 1170 8590
rect 1230 8530 1240 8590
rect 1160 8520 1240 8530
rect 2190 8590 2270 8600
rect 2190 8530 2200 8590
rect 2260 8530 2270 8590
rect 2190 8520 2270 8530
rect 4110 8540 4370 8550
rect -1780 8510 -680 8520
rect 4110 8480 4120 8540
rect 4180 8480 4300 8540
rect 4360 8480 4370 8540
rect 4110 8470 4370 8480
rect 3010 8200 3090 8210
rect -980 8140 -880 8180
rect -980 8080 -960 8140
rect -900 8100 -880 8140
rect 3010 8140 3020 8200
rect 3080 8140 3090 8200
rect 3010 8130 3090 8140
rect 3640 8200 4290 8210
rect 3640 8140 3650 8200
rect 3710 8140 4220 8200
rect 4280 8140 4290 8200
rect 3640 8130 4290 8140
rect 4450 8160 8570 8170
rect 4450 8100 4490 8160
rect 4550 8100 4590 8160
rect 4650 8100 5460 8160
rect 5520 8100 5680 8160
rect 5740 8100 6120 8160
rect 6180 8100 6440 8160
rect 6500 8100 6760 8160
rect 6820 8100 7200 8160
rect 7260 8100 7520 8160
rect 7580 8100 7840 8160
rect 7900 8100 8280 8160
rect 8340 8100 8500 8160
rect 8560 8100 8570 8160
rect -900 8090 4040 8100
rect 4450 8090 8570 8100
rect -900 8080 -630 8090
rect -980 8040 -630 8080
rect -980 7980 -960 8040
rect -900 8030 -630 8040
rect -570 8030 -410 8090
rect -350 8030 -110 8090
rect -50 8030 120 8090
rect 180 8030 270 8090
rect 330 8030 490 8090
rect 550 8030 790 8090
rect 850 8030 1010 8090
rect 1070 8030 1410 8090
rect 1470 8030 1740 8090
rect 1800 8030 2070 8090
rect 2130 8030 2510 8090
rect 2570 8030 2770 8090
rect 2830 8030 3290 8090
rect 3350 8030 3970 8090
rect 4030 8030 4040 8090
rect 9200 8030 9310 8040
rect -900 8020 4040 8030
rect 4210 8020 9310 8030
rect -900 7980 -880 8020
rect -980 7940 -880 7980
rect 4210 7960 4220 8020
rect 4280 7960 9220 8020
rect 4210 7950 9220 7960
rect 9290 7950 9310 8020
rect 9200 7930 9310 7950
rect 5250 7890 12080 7900
rect 5250 7830 5260 7890
rect 5320 7830 12010 7890
rect 12070 7830 12080 7890
rect 5250 7820 12080 7830
rect 5140 7780 12190 7790
rect 5140 7720 5150 7780
rect 5210 7720 12120 7780
rect 12180 7720 12190 7780
rect 5140 7700 12190 7720
rect 5140 7640 5150 7700
rect 5210 7640 12120 7700
rect 12180 7640 12190 7700
rect 5140 7620 12190 7640
rect 5140 7560 5150 7620
rect 5210 7560 12120 7620
rect 12180 7560 12190 7620
rect 5140 7550 12190 7560
rect 9320 7260 9420 7280
rect 650 7250 5000 7260
rect 650 7190 660 7250
rect 720 7190 880 7250
rect 940 7190 1100 7250
rect 1160 7190 1320 7250
rect 1380 7190 1540 7250
rect 1600 7190 1760 7250
rect 1820 7190 4770 7250
rect 4830 7190 4850 7250
rect 4910 7190 4930 7250
rect 4990 7190 5000 7250
rect 650 7170 5000 7190
rect 9320 7200 9340 7260
rect 9400 7200 9420 7260
rect 9320 7180 9420 7200
rect 650 7110 660 7170
rect 720 7110 880 7170
rect 940 7110 1100 7170
rect 1160 7110 1320 7170
rect 1380 7110 1540 7170
rect 1600 7110 1760 7170
rect 1820 7110 4770 7170
rect 4830 7110 4850 7170
rect 4910 7110 4930 7170
rect 4990 7110 5000 7170
rect 650 7090 5000 7110
rect -2640 7080 -70 7090
rect -2640 7020 -2630 7080
rect -2570 7020 -1240 7080
rect -1180 7020 -1020 7080
rect -960 7020 -800 7080
rect -740 7020 -580 7080
rect -520 7020 -360 7080
rect -300 7020 -140 7080
rect -80 7020 -70 7080
rect 650 7030 660 7090
rect 720 7030 880 7090
rect 940 7030 1100 7090
rect 1160 7030 1320 7090
rect 1380 7030 1540 7090
rect 1600 7030 1760 7090
rect 1820 7030 4770 7090
rect 4830 7030 4850 7090
rect 4910 7030 4930 7090
rect 4990 7030 5000 7090
rect 650 7020 5000 7030
rect -2640 7010 -70 7020
rect 4150 6980 4390 6990
rect -1360 6970 4390 6980
rect -1360 6910 -1350 6970
rect -1290 6910 -1130 6970
rect -1070 6910 -910 6970
rect -850 6910 -690 6970
rect -630 6910 -470 6970
rect -410 6910 -250 6970
rect -190 6910 -30 6970
rect 30 6910 550 6970
rect 610 6910 770 6970
rect 830 6910 990 6970
rect 1050 6910 1210 6970
rect 1270 6910 1430 6970
rect 1490 6910 1650 6970
rect 1710 6910 1870 6970
rect 1930 6910 4190 6970
rect 4250 6910 4290 6970
rect 4350 6910 4390 6970
rect -1360 6900 4390 6910
rect 4150 6890 4390 6900
rect 4450 6740 9200 6750
rect 4450 6680 4490 6740
rect 4550 6680 4590 6740
rect 4650 6680 9130 6740
rect 9190 6680 9200 6740
rect 4450 6670 9200 6680
rect -2870 6632 1764 6640
rect -2870 6630 -1182 6632
rect -2870 6570 -2860 6630
rect -2800 6580 -1182 6630
rect -1130 6580 -1072 6632
rect -1020 6580 -962 6632
rect -910 6580 -852 6632
rect -800 6580 -742 6632
rect -690 6580 -632 6632
rect -580 6580 -522 6632
rect -470 6580 -412 6632
rect -360 6580 -302 6632
rect -250 6580 -192 6632
rect -140 6580 718 6632
rect 770 6580 828 6632
rect 880 6580 938 6632
rect 990 6580 1048 6632
rect 1100 6580 1158 6632
rect 1210 6580 1268 6632
rect 1320 6580 1378 6632
rect 1430 6580 1488 6632
rect 1540 6580 1598 6632
rect 1650 6580 1708 6632
rect 1760 6580 1764 6632
rect -2800 6570 1764 6580
rect -1370 6530 4390 6540
rect -1370 6470 -1360 6530
rect -1300 6470 -1000 6530
rect -940 6470 -640 6530
rect -580 6470 -280 6530
rect -220 6470 80 6530
rect 140 6470 440 6530
rect 500 6470 800 6530
rect 860 6470 1160 6530
rect 1220 6470 1520 6530
rect 1580 6470 1880 6530
rect 1940 6470 2510 6530
rect 2570 6470 2950 6530
rect 3010 6500 4390 6530
rect 3010 6470 4190 6500
rect -1370 6450 4190 6470
rect -1370 6390 -1360 6450
rect -1300 6390 -1000 6450
rect -940 6390 -640 6450
rect -580 6390 -280 6450
rect -220 6390 80 6450
rect 140 6390 440 6450
rect 500 6390 800 6450
rect 860 6390 1160 6450
rect 1220 6390 1520 6450
rect 1580 6390 1880 6450
rect 1940 6390 2510 6450
rect 2570 6390 2950 6450
rect 3010 6440 4190 6450
rect 4250 6440 4290 6500
rect 4350 6440 4390 6500
rect 3010 6400 4390 6440
rect 3010 6390 4190 6400
rect -1370 6370 4190 6390
rect -1370 6310 -1360 6370
rect -1300 6310 -1000 6370
rect -940 6310 -640 6370
rect -580 6310 -280 6370
rect -220 6310 80 6370
rect 140 6310 440 6370
rect 500 6310 800 6370
rect 860 6310 1160 6370
rect 1220 6310 1520 6370
rect 1580 6310 1880 6370
rect 1940 6310 2510 6370
rect 2570 6310 2950 6370
rect 3010 6340 4190 6370
rect 4250 6340 4290 6400
rect 4350 6340 4390 6400
rect 3010 6310 4390 6340
rect -1370 6300 4390 6310
rect 5250 6350 5330 6360
rect 5250 6290 5260 6350
rect 5320 6290 5330 6350
rect 5250 6280 5330 6290
rect 2250 6170 2330 6180
rect 2250 6110 2260 6170
rect 2320 6160 2330 6170
rect 2720 6170 2800 6180
rect 2720 6160 2730 6170
rect 2320 6120 2730 6160
rect 2320 6110 2330 6120
rect 2250 6100 2330 6110
rect 2720 6110 2730 6120
rect 2790 6110 2800 6170
rect 2720 6100 2800 6110
rect 2600 5830 2920 5840
rect 2600 5770 2610 5830
rect 2670 5770 2850 5830
rect 2910 5770 2920 5830
rect 2600 5760 2920 5770
rect 7090 5730 7170 5740
rect 7090 5670 7100 5730
rect 7160 5670 7170 5730
rect 7090 5660 7170 5670
rect -1090 5630 1670 5640
rect -1030 5570 -910 5630
rect -850 5570 -730 5630
rect -670 5570 -550 5630
rect -490 5570 -370 5630
rect -310 5570 -190 5630
rect -130 5570 -10 5630
rect 50 5570 170 5630
rect 230 5570 350 5630
rect 410 5570 440 5630
rect 500 5570 530 5630
rect 590 5570 710 5630
rect 770 5570 890 5630
rect 950 5570 1070 5630
rect 1130 5570 1250 5630
rect 1310 5570 1430 5630
rect 1490 5570 1610 5630
rect -1090 5560 1670 5570
rect 4450 5630 4690 5640
rect 4450 5620 8310 5630
rect 4450 5560 4490 5620
rect 4550 5560 4590 5620
rect 4650 5560 5520 5620
rect 5580 5560 5720 5620
rect 5780 5560 5960 5620
rect 6020 5560 6120 5620
rect 6180 5560 6520 5620
rect 6580 5560 6920 5620
rect 6980 5560 7320 5620
rect 7380 5560 7520 5620
rect 7580 5560 8240 5620
rect 8300 5560 8310 5620
rect 4450 5550 8310 5560
rect 4450 5540 4690 5550
rect -110 5520 3240 5530
rect -110 5460 -100 5520
rect -40 5460 620 5520
rect 680 5460 3170 5520
rect 3230 5460 3240 5520
rect -110 5450 3240 5460
rect 7090 5510 7170 5520
rect 7090 5450 7100 5510
rect 7160 5450 7170 5510
rect 7090 5440 7170 5450
rect -470 5410 3330 5420
rect -470 5350 -460 5410
rect -400 5350 980 5410
rect 1040 5350 2260 5410
rect 2320 5350 3260 5410
rect 3320 5350 3330 5410
rect -470 5340 3330 5350
rect 9550 5330 9660 5350
rect -2980 5300 2800 5310
rect -2980 5240 -2970 5300
rect -2910 5240 -820 5300
rect -760 5240 1340 5300
rect 1400 5240 2730 5300
rect 2790 5240 2800 5300
rect 9550 5260 9570 5330
rect 9640 5260 9660 5330
rect 9550 5240 9660 5260
rect -2980 5230 2800 5240
rect 6870 5230 6950 5240
rect -2750 5190 1770 5200
rect -2750 5130 -2740 5190
rect -2680 5130 -1180 5190
rect -1120 5130 260 5190
rect 320 5130 1700 5190
rect 1760 5130 1770 5190
rect 6870 5170 6880 5230
rect 6940 5170 6950 5230
rect 6170 5160 6250 5170
rect 6870 5160 6950 5170
rect 7310 5230 7390 5240
rect 7310 5170 7320 5230
rect 7380 5170 7390 5230
rect -2750 5120 1770 5130
rect 5030 5140 5110 5150
rect -2470 5080 4390 5090
rect -2470 5020 -2460 5080
rect -2400 5020 -2220 5080
rect -2160 5020 -1980 5080
rect -1920 5020 -1740 5080
rect -1680 5020 -1500 5080
rect -1440 5020 -1260 5080
rect -1200 5020 -1020 5080
rect -960 5020 -780 5080
rect -720 5020 -540 5080
rect -480 5020 -300 5080
rect -240 5020 -60 5080
rect 0 5020 580 5080
rect 640 5020 820 5080
rect 880 5020 1060 5080
rect 1120 5020 1300 5080
rect 1360 5020 1540 5080
rect 1600 5020 1780 5080
rect 1840 5020 2020 5080
rect 2080 5020 2260 5080
rect 2320 5020 2500 5080
rect 2560 5020 2740 5080
rect 2800 5020 2980 5080
rect 3040 5050 4390 5080
rect 5030 5080 5040 5140
rect 5100 5130 5110 5140
rect 6170 5130 6180 5160
rect 5100 5100 6180 5130
rect 6240 5130 6250 5160
rect 7310 5130 7390 5170
rect 8850 5230 9410 5240
rect 8850 5170 8860 5230
rect 8920 5170 9340 5230
rect 9400 5170 9410 5230
rect 8850 5160 9410 5170
rect 6240 5100 7390 5130
rect 5100 5090 7390 5100
rect 8010 5110 8090 5120
rect 5100 5080 5110 5090
rect 5030 5070 5110 5080
rect 3040 5020 4190 5050
rect -2470 5000 4190 5020
rect -2470 4940 -2460 5000
rect -2400 4940 -2220 5000
rect -2160 4940 -1980 5000
rect -1920 4940 -1740 5000
rect -1680 4940 -1500 5000
rect -1440 4940 -1260 5000
rect -1200 4940 -1020 5000
rect -960 4940 -780 5000
rect -720 4940 -540 5000
rect -480 4940 -300 5000
rect -240 4940 -60 5000
rect 0 4940 580 5000
rect 640 4940 820 5000
rect 880 4940 1060 5000
rect 1120 4940 1300 5000
rect 1360 4940 1540 5000
rect 1600 4940 1780 5000
rect 1840 4940 2020 5000
rect 2080 4940 2260 5000
rect 2320 4940 2500 5000
rect 2560 4940 2740 5000
rect 2800 4940 2980 5000
rect 3040 4990 4190 5000
rect 4250 4990 4290 5050
rect 4350 4990 4390 5050
rect 6080 5000 6090 5060
rect 6150 5050 6160 5060
rect 8010 5050 8020 5110
rect 8080 5050 8090 5110
rect 6150 5010 8090 5050
rect 9720 5060 12130 5070
rect 6150 5000 6160 5010
rect 9720 5000 9730 5060
rect 9790 5000 12130 5060
rect 9720 4990 12130 5000
rect 3040 4950 4390 4990
rect 3040 4940 4190 4950
rect -2470 4920 4190 4940
rect -2470 4860 -2460 4920
rect -2400 4860 -2220 4920
rect -2160 4860 -1980 4920
rect -1920 4860 -1740 4920
rect -1680 4860 -1500 4920
rect -1440 4860 -1260 4920
rect -1200 4860 -1020 4920
rect -960 4860 -780 4920
rect -720 4860 -540 4920
rect -480 4860 -300 4920
rect -240 4860 -60 4920
rect 0 4860 580 4920
rect 640 4860 820 4920
rect 880 4860 1060 4920
rect 1120 4860 1300 4920
rect 1360 4860 1540 4920
rect 1600 4860 1780 4920
rect 1840 4860 2020 4920
rect 2080 4860 2260 4920
rect 2320 4860 2500 4920
rect 2560 4860 2740 4920
rect 2800 4860 2980 4920
rect 3040 4890 4190 4920
rect 4250 4890 4290 4950
rect 4350 4890 4390 4950
rect 5140 4980 5220 4990
rect 5140 4920 5150 4980
rect 5210 4970 5220 4980
rect 6830 4970 6840 4980
rect 5210 4930 6840 4970
rect 5210 4920 5220 4930
rect 5140 4910 5220 4920
rect 3040 4860 4390 4890
rect -2470 4850 4390 4860
rect 5730 4890 5810 4930
rect 6830 4920 6840 4930
rect 6900 4920 6910 4980
rect 7240 4910 7320 4920
rect 5730 4830 5740 4890
rect 5800 4830 5810 4890
rect 5730 4820 5810 4830
rect 6170 4890 6250 4900
rect 6170 4830 6180 4890
rect 6240 4830 6250 4890
rect 7240 4850 7250 4910
rect 7310 4900 7320 4910
rect 7310 4890 8090 4900
rect 7310 4860 8020 4890
rect 7310 4850 7320 4860
rect 7240 4840 7320 4850
rect 6170 4820 6250 4830
rect 8010 4830 8020 4860
rect 8080 4830 8090 4890
rect 8010 4820 8090 4830
rect 8850 4890 9410 4900
rect 8850 4830 8860 4890
rect 8920 4830 9340 4890
rect 9400 4830 9410 4890
rect 8850 4820 9410 4830
rect 9550 4820 9660 4840
rect -2870 4810 150 4820
rect -2870 4750 -2860 4810
rect -2800 4750 -2340 4810
rect -2280 4750 -1620 4810
rect -1560 4750 -900 4810
rect -840 4750 -180 4810
rect -120 4750 80 4810
rect 140 4750 150 4810
rect -2870 4740 150 4750
rect 430 4810 3560 4820
rect 430 4750 440 4810
rect 500 4750 700 4810
rect 760 4750 1420 4810
rect 1480 4750 2140 4810
rect 2200 4750 2860 4810
rect 2920 4750 3490 4810
rect 3550 4750 3560 4810
rect 430 4740 3560 4750
rect 9550 4750 9570 4820
rect 9640 4750 9660 4820
rect -1620 4710 -1560 4740
rect 2140 4700 2200 4740
rect 9550 4730 9660 4750
rect 6030 4510 6110 4520
rect -2110 4470 -2030 4480
rect -2110 4410 -2100 4470
rect -2040 4460 -2030 4470
rect -1390 4470 -1310 4480
rect -1390 4460 -1380 4470
rect -2040 4420 -1380 4460
rect -2040 4410 -2030 4420
rect -2110 4400 -2030 4410
rect -1390 4410 -1380 4420
rect -1320 4460 -1310 4470
rect -670 4470 -590 4480
rect -670 4460 -660 4470
rect -1320 4420 -660 4460
rect -1320 4410 -1310 4420
rect -1390 4400 -1310 4410
rect -670 4410 -660 4420
rect -600 4410 -590 4470
rect -670 4400 -590 4410
rect 1170 4470 1250 4480
rect 1170 4410 1180 4470
rect 1240 4460 1250 4470
rect 1890 4470 1970 4480
rect 1890 4460 1900 4470
rect 1240 4420 1900 4460
rect 1240 4410 1250 4420
rect 1170 4400 1250 4410
rect 1890 4410 1900 4420
rect 1960 4460 1970 4470
rect 2610 4470 2690 4480
rect 2610 4460 2620 4470
rect 1960 4420 2620 4460
rect 1960 4410 1970 4420
rect 1890 4400 1970 4410
rect 2610 4410 2620 4420
rect 2680 4410 2690 4470
rect 6030 4450 6040 4510
rect 6100 4450 6110 4510
rect 6030 4440 6110 4450
rect 2610 4400 2690 4410
rect 4150 4410 4390 4420
rect 4150 4400 8310 4410
rect -2370 4350 -170 4360
rect -2370 4290 -2360 4350
rect -2300 4290 -2280 4350
rect -2220 4290 -1860 4350
rect -1800 4290 -1620 4350
rect -1560 4290 -1140 4350
rect -1080 4290 -900 4350
rect -840 4290 -420 4350
rect -360 4290 -240 4350
rect -180 4290 -170 4350
rect -2370 4280 -170 4290
rect 750 4350 3830 4360
rect 750 4290 760 4350
rect 820 4290 940 4350
rect 1000 4290 1180 4350
rect 1240 4290 1420 4350
rect 1480 4290 1660 4350
rect 1720 4290 2140 4350
rect 2200 4290 2380 4350
rect 2440 4290 2800 4350
rect 2860 4290 3600 4350
rect 3660 4290 3680 4350
rect 3740 4290 3760 4350
rect 3820 4290 3830 4350
rect 4150 4340 4190 4400
rect 4250 4340 4290 4400
rect 4350 4340 5640 4400
rect 5700 4340 5840 4400
rect 5900 4340 6240 4400
rect 6300 4340 6640 4400
rect 6700 4340 7040 4400
rect 7100 4340 7120 4400
rect 7180 4340 7440 4400
rect 7500 4340 7640 4400
rect 7700 4340 8240 4400
rect 8300 4340 8310 4400
rect 4150 4330 8310 4340
rect 4150 4320 4390 4330
rect 750 4270 3830 4290
rect 750 4210 760 4270
rect 820 4210 940 4270
rect 1000 4210 1180 4270
rect 1240 4210 1420 4270
rect 1480 4210 1660 4270
rect 1720 4210 2140 4270
rect 2200 4210 2380 4270
rect 2440 4210 2800 4270
rect 2860 4210 3600 4270
rect 3660 4210 3680 4270
rect 3740 4210 3760 4270
rect 3820 4210 3830 4270
rect 750 4190 3830 4210
rect 6030 4260 7310 4270
rect 6030 4200 6040 4260
rect 6100 4200 7240 4260
rect 7300 4200 7310 4260
rect 6030 4190 7310 4200
rect 750 4130 760 4190
rect 820 4130 940 4190
rect 1000 4130 1180 4190
rect 1240 4130 1420 4190
rect 1480 4130 1660 4190
rect 1720 4130 2140 4190
rect 2200 4130 2380 4190
rect 2440 4130 2800 4190
rect 2860 4130 3600 4190
rect 3660 4130 3680 4190
rect 3740 4130 3760 4190
rect 3820 4130 3830 4190
rect 750 4120 3830 4130
rect -1630 4080 -590 4090
rect -1630 4020 -1620 4080
rect -1560 4020 -1140 4080
rect -1080 4020 -660 4080
rect -600 4020 -590 4080
rect -1630 4010 -590 4020
rect 1170 4080 2210 4090
rect 1170 4020 1180 4080
rect 1240 4020 1660 4080
rect 1720 4020 2140 4080
rect 2200 4020 2210 4080
rect 1170 4010 2210 4020
rect -1390 3970 -350 3980
rect -1390 3910 -1380 3970
rect -1320 3910 -900 3970
rect -840 3910 -420 3970
rect -360 3910 -350 3970
rect -1390 3900 -350 3910
rect 930 3970 1970 3980
rect 930 3910 940 3970
rect 1000 3910 1420 3970
rect 1480 3910 1900 3970
rect 1960 3910 1970 3970
rect 930 3900 1970 3910
rect -2750 3870 -2670 3880
rect 3250 3870 3330 3880
rect -2750 3810 -2740 3870
rect -2680 3860 -440 3870
rect -2680 3810 -1454 3860
rect -2750 3808 -1454 3810
rect -1402 3808 -1296 3860
rect -1244 3808 -972 3860
rect -920 3808 -818 3860
rect -766 3808 -494 3860
rect -442 3808 -440 3860
rect 1020 3860 3260 3870
rect -2750 3800 -440 3808
rect -190 3820 770 3830
rect -190 3760 -180 3820
rect -120 3760 180 3820
rect 240 3760 260 3820
rect 320 3760 340 3820
rect 400 3760 700 3820
rect 760 3760 770 3820
rect 1020 3808 1022 3860
rect 1074 3808 1346 3860
rect 1398 3808 1500 3860
rect 1552 3808 1824 3860
rect 1876 3808 1982 3860
rect 2034 3810 3260 3860
rect 3320 3810 3330 3870
rect 2034 3808 3330 3810
rect 1020 3800 3330 3808
rect -190 3740 770 3760
rect -190 3680 -180 3740
rect -120 3680 180 3740
rect 240 3680 260 3740
rect 320 3680 340 3740
rect 400 3680 700 3740
rect 760 3680 770 3740
rect -190 3660 770 3680
rect -2640 3640 -2560 3650
rect -2640 3580 -2630 3640
rect -2570 3632 -541 3640
rect -2570 3580 -1557 3632
rect -1505 3580 -1197 3632
rect -1145 3580 -1077 3632
rect -1025 3580 -717 3632
rect -665 3580 -597 3632
rect -545 3580 -541 3632
rect -190 3600 -180 3660
rect -120 3600 180 3660
rect 240 3600 260 3660
rect 320 3600 340 3660
rect 400 3600 700 3660
rect 760 3600 770 3660
rect 3160 3640 3240 3650
rect -190 3590 770 3600
rect 1121 3632 3170 3640
rect -2640 3570 -541 3580
rect 1121 3580 1125 3632
rect 1177 3580 1245 3632
rect 1297 3580 1605 3632
rect 1657 3580 1725 3632
rect 1777 3580 2085 3632
rect 2137 3580 3170 3632
rect 3230 3580 3240 3640
rect 1121 3570 3240 3580
rect 5250 3600 6910 3610
rect 5250 3540 5260 3600
rect 5320 3540 6440 3600
rect 6500 3540 6840 3600
rect 6900 3540 6910 3600
rect -2250 3530 -460 3540
rect -2250 3470 -2240 3530
rect -2180 3470 -1490 3530
rect -1430 3470 -1270 3530
rect -1210 3470 -1010 3530
rect -950 3470 -790 3530
rect -730 3470 -530 3530
rect -470 3470 -460 3530
rect -2250 3460 -460 3470
rect 1040 3530 2830 3540
rect 5250 3530 6910 3540
rect 1040 3470 1050 3530
rect 1110 3470 1310 3530
rect 1370 3470 1530 3530
rect 1590 3470 1790 3530
rect 1850 3470 2010 3530
rect 2070 3470 2760 3530
rect 2820 3470 2830 3530
rect 1040 3460 2830 3470
rect -2070 3420 4390 3430
rect -2070 3360 -2060 3420
rect -2000 3360 -1820 3420
rect -1760 3360 -1580 3420
rect -1520 3360 -1340 3420
rect -1280 3360 -700 3420
rect -640 3360 -460 3420
rect -400 3360 -220 3420
rect -160 3360 740 3420
rect 800 3360 980 3420
rect 1040 3360 1220 3420
rect 1280 3360 1860 3420
rect 1920 3360 2100 3420
rect 2160 3360 2340 3420
rect 2400 3360 2580 3420
rect 2640 3390 4390 3420
rect 2640 3360 4190 3390
rect -2070 3340 4190 3360
rect -2070 3280 -2060 3340
rect -2000 3280 -1820 3340
rect -1760 3280 -1580 3340
rect -1520 3280 -1340 3340
rect -1280 3280 -700 3340
rect -640 3280 -460 3340
rect -400 3280 -220 3340
rect -160 3280 740 3340
rect 800 3280 980 3340
rect 1040 3280 1220 3340
rect 1280 3280 1860 3340
rect 1920 3280 2100 3340
rect 2160 3280 2340 3340
rect 2400 3280 2580 3340
rect 2640 3330 4190 3340
rect 4250 3330 4290 3390
rect 4350 3330 4390 3390
rect 2640 3290 4390 3330
rect 2640 3280 4190 3290
rect -2070 3260 4190 3280
rect -2070 3200 -2060 3260
rect -2000 3200 -1820 3260
rect -1760 3200 -1580 3260
rect -1520 3200 -1340 3260
rect -1280 3200 -700 3260
rect -640 3200 -460 3260
rect -400 3200 -220 3260
rect -160 3200 740 3260
rect 800 3200 980 3260
rect 1040 3200 1220 3260
rect 1280 3200 1860 3260
rect 1920 3200 2100 3260
rect 2160 3200 2340 3260
rect 2400 3200 2580 3260
rect 2640 3230 4190 3260
rect 4250 3230 4290 3290
rect 4350 3230 4390 3290
rect 2640 3200 4390 3230
rect -2070 3190 4390 3200
rect 4450 3210 9200 3220
rect 4450 3150 4490 3210
rect 4550 3150 4590 3210
rect 4650 3150 9130 3210
rect 9190 3150 9200 3210
rect 4450 3140 9200 3150
rect 4150 2970 4390 2990
rect 4150 2910 4190 2970
rect 4250 2910 4290 2970
rect 4350 2910 4390 2970
rect 4150 2890 4390 2910
rect 9320 2880 9420 2900
rect 9320 2820 9340 2880
rect 9400 2820 9420 2880
rect 9320 2800 9420 2820
rect -1090 2620 4690 2630
rect -1090 2560 -1080 2620
rect -1020 2560 180 2620
rect 240 2560 260 2620
rect 320 2560 340 2620
rect 400 2560 1600 2620
rect 1660 2590 4690 2620
rect 1660 2560 4490 2590
rect -1090 2540 4490 2560
rect -1090 2480 -1080 2540
rect -1020 2480 180 2540
rect 240 2480 260 2540
rect 320 2480 340 2540
rect 400 2480 1600 2540
rect 1660 2530 4490 2540
rect 4550 2530 4590 2590
rect 4650 2530 4690 2590
rect 1660 2490 4690 2530
rect 1660 2480 4490 2490
rect -1090 2460 4490 2480
rect -1090 2400 -1080 2460
rect -1020 2400 180 2460
rect 240 2400 260 2460
rect 320 2400 340 2460
rect 400 2400 1600 2460
rect 1660 2430 4490 2460
rect 4550 2430 4590 2490
rect 4650 2430 4690 2490
rect 1660 2400 4690 2430
rect -1090 2390 4690 2400
rect -1830 2350 -1750 2360
rect -1830 2290 -1820 2350
rect -1760 2340 -1750 2350
rect -1670 2350 -1590 2360
rect -1670 2340 -1660 2350
rect -1760 2300 -1660 2340
rect -1760 2290 -1750 2300
rect -1830 2280 -1750 2290
rect -1670 2290 -1660 2300
rect -1600 2340 -1590 2350
rect -1510 2350 -1430 2360
rect -1510 2340 -1500 2350
rect -1600 2300 -1500 2340
rect -1600 2290 -1590 2300
rect -1670 2280 -1590 2290
rect -1510 2290 -1500 2300
rect -1440 2340 -1430 2350
rect -1350 2350 -1270 2360
rect -1350 2340 -1340 2350
rect -1440 2300 -1340 2340
rect -1440 2290 -1430 2300
rect -1510 2280 -1430 2290
rect -1350 2290 -1340 2300
rect -1280 2340 -1270 2350
rect -1190 2350 -1110 2360
rect -1190 2340 -1180 2350
rect -1280 2300 -1180 2340
rect -1280 2290 -1270 2300
rect -1350 2280 -1270 2290
rect -1190 2290 -1180 2300
rect -1120 2340 -1110 2350
rect -1030 2350 -950 2360
rect -1030 2340 -1020 2350
rect -1120 2300 -1020 2340
rect -1120 2290 -1110 2300
rect -1190 2280 -1110 2290
rect -1030 2290 -1020 2300
rect -960 2340 -950 2350
rect -870 2350 -790 2360
rect -870 2340 -860 2350
rect -960 2300 -860 2340
rect -960 2290 -950 2300
rect -1030 2280 -950 2290
rect -870 2290 -860 2300
rect -800 2340 -790 2350
rect -710 2350 -630 2360
rect -710 2340 -700 2350
rect -800 2300 -700 2340
rect -800 2290 -790 2300
rect -870 2280 -790 2290
rect -710 2290 -700 2300
rect -640 2340 -630 2350
rect -550 2350 -470 2360
rect -550 2340 -540 2350
rect -640 2300 -540 2340
rect -640 2290 -630 2300
rect -710 2280 -630 2290
rect -550 2290 -540 2300
rect -480 2340 -470 2350
rect -390 2350 -310 2360
rect -390 2340 -380 2350
rect -480 2300 -380 2340
rect -480 2290 -470 2300
rect -550 2280 -470 2290
rect -390 2290 -380 2300
rect -320 2340 -310 2350
rect -230 2350 -150 2360
rect -230 2340 -220 2350
rect -320 2300 -220 2340
rect -320 2290 -310 2300
rect -390 2280 -310 2290
rect -230 2290 -220 2300
rect -160 2340 -150 2350
rect -70 2350 10 2360
rect -70 2340 -60 2350
rect -160 2300 -60 2340
rect -160 2290 -150 2300
rect -230 2280 -150 2290
rect -70 2290 -60 2300
rect 0 2340 10 2350
rect 90 2350 170 2360
rect 90 2340 100 2350
rect 0 2300 100 2340
rect 0 2290 10 2300
rect -70 2280 10 2290
rect 90 2290 100 2300
rect 160 2290 170 2350
rect 90 2280 170 2290
rect 250 2350 330 2360
rect 250 2290 260 2350
rect 320 2340 330 2350
rect 410 2350 490 2360
rect 410 2340 420 2350
rect 320 2300 420 2340
rect 320 2290 330 2300
rect 250 2280 330 2290
rect 410 2290 420 2300
rect 480 2340 490 2350
rect 570 2350 650 2360
rect 570 2340 580 2350
rect 480 2300 580 2340
rect 480 2290 490 2300
rect 410 2280 490 2290
rect 570 2290 580 2300
rect 640 2340 650 2350
rect 730 2350 810 2360
rect 730 2340 740 2350
rect 640 2300 740 2340
rect 640 2290 650 2300
rect 570 2280 650 2290
rect 730 2290 740 2300
rect 800 2340 810 2350
rect 890 2350 970 2360
rect 890 2340 900 2350
rect 800 2300 900 2340
rect 800 2290 810 2300
rect 730 2280 810 2290
rect 890 2290 900 2300
rect 960 2340 970 2350
rect 1050 2350 1130 2360
rect 1050 2340 1060 2350
rect 960 2300 1060 2340
rect 960 2290 970 2300
rect 890 2280 970 2290
rect 1050 2290 1060 2300
rect 1120 2340 1130 2350
rect 1210 2350 1290 2360
rect 1210 2340 1220 2350
rect 1120 2300 1220 2340
rect 1120 2290 1130 2300
rect 1050 2280 1130 2290
rect 1210 2290 1220 2300
rect 1280 2340 1290 2350
rect 1370 2350 1450 2360
rect 1370 2340 1380 2350
rect 1280 2300 1380 2340
rect 1280 2290 1290 2300
rect 1210 2280 1290 2290
rect 1370 2290 1380 2300
rect 1440 2340 1450 2350
rect 1530 2350 1610 2360
rect 1530 2340 1540 2350
rect 1440 2300 1540 2340
rect 1440 2290 1450 2300
rect 1370 2280 1450 2290
rect 1530 2290 1540 2300
rect 1600 2340 1610 2350
rect 1690 2350 1770 2360
rect 1690 2340 1700 2350
rect 1600 2300 1700 2340
rect 1600 2290 1610 2300
rect 1530 2280 1610 2290
rect 1690 2290 1700 2300
rect 1760 2340 1770 2350
rect 1850 2350 1930 2360
rect 1850 2340 1860 2350
rect 1760 2300 1860 2340
rect 1760 2290 1770 2300
rect 1690 2280 1770 2290
rect 1850 2290 1860 2300
rect 1920 2340 1930 2350
rect 2010 2350 2090 2360
rect 2010 2340 2020 2350
rect 1920 2300 2020 2340
rect 1920 2290 1930 2300
rect 1850 2280 1930 2290
rect 2010 2290 2020 2300
rect 2080 2340 2090 2350
rect 2170 2350 2250 2360
rect 2170 2340 2180 2350
rect 2080 2300 2180 2340
rect 2080 2290 2090 2300
rect 2010 2280 2090 2290
rect 2170 2290 2180 2300
rect 2240 2290 2250 2350
rect 2170 2280 2250 2290
rect 2480 2220 4690 2230
rect -2980 2180 -1830 2190
rect -2980 2120 -2970 2180
rect -2910 2120 -1900 2180
rect -1840 2120 -1830 2180
rect -2980 2110 -1830 2120
rect 2480 2160 2490 2220
rect 2550 2180 4690 2220
rect 2550 2160 4490 2180
rect 2480 2140 4490 2160
rect 2480 2080 2490 2140
rect 2550 2120 4490 2140
rect 4550 2120 4590 2180
rect 4650 2120 4690 2180
rect 2550 2080 4690 2120
rect 2480 2070 4690 2080
rect -2370 2010 4060 2020
rect -2370 1950 -2360 2010
rect -2300 1950 -1950 2010
rect -1890 1950 3990 2010
rect 4050 1950 4060 2010
rect -2370 1940 4060 1950
rect -2640 1900 2900 1910
rect -2640 1840 -2630 1900
rect -2570 1840 2830 1900
rect 2890 1840 2900 1900
rect -2640 1830 2900 1840
rect 3160 1790 3240 1800
rect -1850 1780 -438 1790
rect -1850 1720 -1840 1780
rect -1780 1720 -438 1780
rect -368 1720 -358 1790
rect 950 1720 960 1790
rect 1030 1780 1040 1790
rect 3160 1780 3170 1790
rect 1030 1740 3170 1780
rect 1030 1720 1040 1740
rect 3160 1730 3170 1740
rect 3230 1730 3240 1790
rect 3160 1720 3240 1730
rect -1850 1710 -440 1720
rect -2320 1670 1040 1680
rect -2320 1610 -2310 1670
rect -2250 1610 970 1670
rect 1030 1610 1040 1670
rect -2320 1600 1040 1610
rect 2350 1590 2430 1600
rect 2350 1530 2360 1590
rect 2420 1580 2430 1590
rect 2700 1590 2780 1600
rect 2700 1580 2710 1590
rect 2420 1540 2710 1580
rect 2420 1530 2430 1540
rect 2350 1520 2430 1530
rect 2700 1530 2710 1540
rect 2770 1580 2780 1590
rect 3250 1590 3330 1600
rect 3250 1580 3260 1590
rect 2770 1540 3260 1580
rect 2770 1530 2780 1540
rect 2700 1520 2780 1530
rect 3250 1530 3260 1540
rect 3320 1530 3330 1590
rect 3250 1520 3330 1530
rect 3590 1040 4190 1060
rect 3590 980 3600 1040
rect 3660 980 3680 1040
rect 3740 980 3760 1040
rect 3820 980 4110 1040
rect 4170 980 4190 1040
rect 3590 960 4190 980
rect 3860 340 4380 350
rect 3860 280 3870 340
rect 3930 280 4310 340
rect 4370 280 4380 340
rect 3860 270 4380 280
rect -2310 -10 -2240 0
rect -2310 -90 -2240 -80
rect 2700 -10 2770 0
rect 2700 -90 2770 -80
rect 3480 -360 4190 -340
rect -2740 -390 -2670 -380
rect -2860 -440 -2790 -430
rect -2740 -470 -2670 -460
rect -1850 -420 -1340 -410
rect -1850 -480 -1840 -420
rect -1780 -480 -1410 -420
rect -1350 -480 -1340 -420
rect -1850 -490 -1340 -480
rect 250 -420 2430 -410
rect 250 -480 260 -420
rect 320 -480 2360 -420
rect 2420 -480 2430 -420
rect 3480 -420 3490 -360
rect 3550 -420 4110 -360
rect 4170 -420 4190 -360
rect 3480 -440 4190 -420
rect 250 -490 2430 -480
rect -2860 -530 -2790 -510
rect 3480 -652 3550 -640
rect 3480 -732 3550 -722
rect 2820 -860 2890 -850
rect 2820 -940 2890 -930
rect 4230 -1060 4310 -1050
rect 4230 -1120 4240 -1060
rect 4300 -1120 4310 -1060
rect 4230 -1130 4310 -1120
rect 3970 -1760 4070 -1740
rect -2860 -1788 -2790 -1778
rect 3970 -1820 3990 -1760
rect 4050 -1820 4070 -1760
rect 3970 -1840 4070 -1820
rect -2860 -1868 -2790 -1858
rect -2850 -1870 -2810 -1868
rect -2500 -1998 -2430 -1988
rect -2500 -2078 -2430 -2068
rect 2820 -1998 2890 -1988
rect 2820 -2078 2890 -2068
rect 3480 -1990 3550 -1988
rect 3480 -1998 3940 -1990
rect 3550 -2000 3940 -1998
rect 3550 -2068 3860 -2000
rect 3480 -2070 3860 -2068
rect 3930 -2070 3940 -2000
rect -2480 -2080 -2440 -2078
rect 2830 -2080 2870 -2078
rect 3480 -2080 3940 -2070
rect -2070 -2148 -2000 -2138
rect -2070 -2228 -2000 -2218
rect 2460 -2148 2530 -2138
rect 2460 -2228 2530 -2218
rect -2050 -2230 -2010 -2228
rect 2470 -2230 2510 -2228
rect 4300 -2460 4380 -2450
rect 4300 -2520 4310 -2460
rect 4370 -2520 4380 -2460
rect -3040 -2530 3070 -2520
rect 4300 -2530 4380 -2520
rect -3040 -2590 -3030 -2530
rect -2970 -2590 -2490 -2530
rect -2430 -2590 -2060 -2530
rect -2000 -2590 260 -2530
rect 320 -2590 2460 -2530
rect 2520 -2590 2820 -2530
rect 2880 -2590 3000 -2530
rect 3060 -2590 3070 -2530
rect -3040 -2610 3070 -2590
rect -3040 -2670 -3030 -2610
rect -2970 -2670 -2490 -2610
rect -2430 -2670 -2060 -2610
rect -2000 -2670 260 -2610
rect 320 -2670 2460 -2610
rect 2520 -2670 2820 -2610
rect 2880 -2670 3000 -2610
rect 3060 -2670 3070 -2610
rect -3040 -2690 3070 -2670
rect -3040 -2750 -3030 -2690
rect -2970 -2750 -2490 -2690
rect -2430 -2750 -2060 -2690
rect -2000 -2750 260 -2690
rect 320 -2750 2460 -2690
rect 2520 -2750 2820 -2690
rect 2880 -2750 3000 -2690
rect 3060 -2750 3070 -2690
rect -3040 -2760 3070 -2750
rect -2870 -2800 4380 -2790
rect -2870 -2860 -2860 -2800
rect -2800 -2860 4310 -2800
rect 4370 -2860 4380 -2800
rect -2870 -2870 4380 -2860
rect -3070 -2900 -2970 -2890
rect 14000 -2900 14100 -2890
rect -3070 -2910 2970 -2900
rect -3070 -2970 -3050 -2910
rect -2990 -2970 2900 -2910
rect 2960 -2970 2970 -2910
rect -3070 -2980 2970 -2970
rect 5340 -2910 14100 -2900
rect 5340 -2970 5350 -2910
rect 5410 -2970 12120 -2910
rect 12180 -2970 14020 -2910
rect 14080 -2970 14100 -2910
rect 5340 -2980 14100 -2970
rect -3070 -2990 -2970 -2980
rect 14000 -2990 14100 -2980
rect -4270 -3290 11420 -3270
rect -4270 -3360 10830 -3290
rect 10900 -3360 11330 -3290
rect 11400 -3360 11420 -3290
rect -4270 -3380 11420 -3360
<< via2 >>
rect 8720 14260 8780 14320
rect 8720 14160 8780 14220
rect -1650 13040 -1590 13100
rect -1650 12940 -1590 13000
rect -1650 12260 -1590 12320
rect -1650 12160 -1590 12220
rect 8720 10740 8780 10800
rect 8720 10640 8780 10700
rect -960 10440 -900 10500
rect -960 10340 -900 10400
rect 9110 10450 9180 10520
rect 5390 9940 5450 10000
rect 5490 9940 5550 10000
rect -960 9260 -900 9320
rect -960 9160 -900 9220
rect 8870 9270 8940 9340
rect 8870 8740 8940 8810
rect -960 8080 -900 8140
rect 4490 8100 4550 8160
rect 4590 8100 4650 8160
rect -960 7980 -900 8040
rect 9220 7950 9290 8020
rect 9340 7200 9400 7260
rect 4190 6910 4250 6970
rect 4290 6910 4350 6970
rect 4490 6680 4550 6740
rect 4590 6680 4650 6740
rect 4190 6440 4250 6500
rect 4290 6440 4350 6500
rect 4190 6340 4250 6400
rect 4290 6340 4350 6400
rect 4490 5560 4550 5620
rect 4590 5560 4650 5620
rect 9570 5260 9640 5330
rect 4190 4990 4250 5050
rect 4290 4990 4350 5050
rect 4190 4890 4250 4950
rect 4290 4890 4350 4950
rect 9570 4750 9640 4820
rect 4190 4340 4250 4400
rect 4290 4340 4350 4400
rect 4190 3330 4250 3390
rect 4290 3330 4350 3390
rect 4190 3230 4250 3290
rect 4290 3230 4350 3290
rect 4490 3150 4550 3210
rect 4590 3150 4650 3210
rect 4190 2910 4250 2970
rect 4290 2910 4350 2970
rect 9340 2820 9400 2880
rect 4490 2530 4550 2590
rect 4590 2530 4650 2590
rect 4490 2430 4550 2490
rect 4590 2430 4650 2490
rect 4490 2120 4550 2180
rect 4590 2120 4650 2180
rect 4110 980 4170 1040
rect 4310 280 4370 340
rect 4110 -420 4170 -360
rect 4240 -1120 4300 -1060
rect 3990 -1820 4050 -1760
rect 4310 -2520 4370 -2460
rect -3050 -2970 -2990 -2910
rect 14020 -2970 14080 -2910
rect 10830 -3360 10900 -3290
rect 11330 -3360 11400 -3290
<< metal3 >>
rect -4270 14320 8800 14360
rect -4270 14260 8720 14320
rect 8780 14260 8800 14320
rect -4270 14220 8800 14260
rect -4270 14160 8720 14220
rect 8780 14160 8800 14220
rect -4270 14120 8800 14160
rect -4270 13100 -1570 13140
rect -4270 13040 -1650 13100
rect -1590 13040 -1570 13100
rect -4270 13000 -1570 13040
rect -4270 12940 -1650 13000
rect -1590 12940 -1570 13000
rect -4270 12900 -1570 12940
rect -4270 12320 -1570 12360
rect -4270 12260 -1650 12320
rect -1590 12260 -1570 12320
rect -4270 12220 -1570 12260
rect -4270 12160 -1650 12220
rect -1590 12160 -1570 12220
rect -4270 12120 -1570 12160
rect -4270 10800 8800 10840
rect -4270 10740 8720 10800
rect 8780 10740 8800 10800
rect -4270 10700 8800 10740
rect -4270 10640 8720 10700
rect 8780 10640 8800 10700
rect -4270 10600 8800 10640
rect -4270 10500 -880 10540
rect -4270 10440 -960 10500
rect -900 10440 -880 10500
rect -4270 10400 -880 10440
rect -4270 10340 -960 10400
rect -900 10340 -880 10400
rect -4270 10300 -880 10340
rect 5350 10000 5590 10600
rect 9090 10520 10300 10540
rect 9090 10450 9110 10520
rect 9180 10450 10300 10520
rect 9090 10430 10300 10450
rect 5350 9940 5390 10000
rect 5450 9940 5490 10000
rect 5550 9940 5590 10000
rect 5350 9930 5590 9940
rect -4270 9320 -880 9360
rect -4270 9260 -960 9320
rect -900 9260 -880 9320
rect -4270 9220 -880 9260
rect 8850 9340 8960 9360
rect 8850 9270 8870 9340
rect 8940 9270 8960 9340
rect 8850 9250 8960 9270
rect 9200 9220 10300 10430
rect -4270 9160 -960 9220
rect -900 9160 -880 9220
rect -4270 9120 -880 9160
rect 8850 8810 8960 8830
rect 8850 8740 8870 8810
rect 8940 8740 8960 8810
rect 8850 8720 8960 8740
rect -4270 8140 -880 8180
rect -4270 8080 -960 8140
rect -900 8080 -880 8140
rect -4270 8040 -880 8080
rect -4270 7980 -960 8040
rect -900 7980 -880 8040
rect -4270 7940 -880 7980
rect 4450 8160 4690 8170
rect 4450 8100 4490 8160
rect 4550 8100 4590 8160
rect 4650 8100 4690 8160
rect 4450 7830 4690 8100
rect 9200 8040 9800 8860
rect 9200 8020 9310 8040
rect 9200 7950 9220 8020
rect 9290 7950 9310 8020
rect 9200 7930 9310 7950
rect -4270 7590 4690 7830
rect -4270 7290 4390 7530
rect 4150 6970 4390 7290
rect 4150 6910 4190 6970
rect 4250 6910 4290 6970
rect 4350 6910 4390 6970
rect 4150 6500 4390 6910
rect 4150 6440 4190 6500
rect 4250 6440 4290 6500
rect 4350 6440 4390 6500
rect 4150 6400 4390 6440
rect 4150 6340 4190 6400
rect 4250 6340 4290 6400
rect 4350 6340 4390 6400
rect 4150 5050 4390 6340
rect 4150 4990 4190 5050
rect 4250 4990 4290 5050
rect 4350 4990 4390 5050
rect 4150 4950 4390 4990
rect 4150 4890 4190 4950
rect 4250 4890 4290 4950
rect 4350 4890 4390 4950
rect 4150 4400 4390 4890
rect 4150 4340 4190 4400
rect 4250 4340 4290 4400
rect 4350 4340 4390 4400
rect 4150 3390 4390 4340
rect 4150 3330 4190 3390
rect 4250 3330 4290 3390
rect 4350 3330 4390 3390
rect 4150 3290 4390 3330
rect 4150 3230 4190 3290
rect 4250 3230 4290 3290
rect 4350 3230 4390 3290
rect 4150 2970 4390 3230
rect 4150 2910 4190 2970
rect 4250 2910 4290 2970
rect 4350 2910 4390 2970
rect 4150 2890 4390 2910
rect 4450 6740 4690 7590
rect 9320 7270 9420 7280
rect 9320 7260 11960 7270
rect 9320 7200 9340 7260
rect 9400 7200 11960 7260
rect 9320 7180 11960 7200
rect 4450 6680 4490 6740
rect 4550 6680 4590 6740
rect 4650 6680 4690 6740
rect 4450 5620 4690 6680
rect 4450 5560 4490 5620
rect 4550 5560 4590 5620
rect 4650 5560 4690 5620
rect 4450 3210 4690 5560
rect 9550 5330 9660 5350
rect 9550 5260 9570 5330
rect 9640 5260 9660 5330
rect 9550 5240 9660 5260
rect 9900 5210 11960 7180
rect 9550 4820 9660 4840
rect 9550 4750 9570 4820
rect 9640 4750 9660 4820
rect 9550 4730 9660 4750
rect 4450 3150 4490 3210
rect 4550 3150 4590 3210
rect 4650 3150 4690 3210
rect 4450 2590 4690 3150
rect 9900 2900 11960 4870
rect 9320 2880 11960 2900
rect 9320 2820 9340 2880
rect 9400 2820 11960 2880
rect 9320 2810 11960 2820
rect 9320 2800 9420 2810
rect 4450 2530 4490 2590
rect 4550 2530 4590 2590
rect 4650 2530 4690 2590
rect 4450 2490 4690 2530
rect 4450 2430 4490 2490
rect 4550 2430 4590 2490
rect 4650 2430 4690 2490
rect 4450 2180 4690 2430
rect 4450 2120 4490 2180
rect 4550 2120 4590 2180
rect 4650 2120 4690 2180
rect 4450 2070 4690 2120
rect 4430 1060 4890 1250
rect 5130 1060 5590 1250
rect 5830 1060 6290 1250
rect 6530 1060 6990 1250
rect 7230 1060 7690 1250
rect 7930 1060 8390 1250
rect 8630 1060 9090 1250
rect 9330 1060 9790 1250
rect 10030 1060 10490 1250
rect 10730 1060 11190 1250
rect 4090 1050 4190 1060
rect 4090 970 4100 1050
rect 4180 970 4190 1050
rect 4090 960 4190 970
rect 4430 960 11190 1060
rect 4430 790 4890 960
rect 5130 790 5590 960
rect 5830 790 6290 960
rect 6530 790 6990 960
rect 7230 790 7690 960
rect 7930 790 8390 960
rect 8630 790 9090 960
rect 9330 790 9790 960
rect 10030 790 10490 960
rect 10730 790 11190 960
rect 10910 550 11010 790
rect 4430 360 4890 550
rect 5130 360 5590 550
rect 5830 360 6290 550
rect 6530 360 6990 550
rect 7230 360 7690 550
rect 7930 360 8390 550
rect 8630 360 9090 550
rect 9330 360 9790 550
rect 10030 360 10490 550
rect 10730 360 11190 550
rect 4430 350 11190 360
rect 4300 340 11190 350
rect 4300 280 4310 340
rect 4370 280 11190 340
rect 4300 270 11190 280
rect 4430 260 11190 270
rect 4430 90 4890 260
rect 5130 90 5590 260
rect 5830 90 6290 260
rect 6530 90 6990 260
rect 7230 90 7690 260
rect 7930 90 8390 260
rect 8630 90 9090 260
rect 9330 90 9790 260
rect 10030 90 10490 260
rect 10730 90 11190 260
rect 4430 -340 4890 -150
rect 5130 -340 5590 -150
rect 5830 -340 6290 -150
rect 6530 -340 6990 -150
rect 7230 -340 7690 -150
rect 7930 -340 8390 -150
rect 8630 -340 9090 -150
rect 9330 -340 9790 -150
rect 10030 -340 10490 -150
rect 10730 -340 11190 -150
rect 4090 -350 4190 -340
rect 4090 -430 4100 -350
rect 4180 -430 4190 -350
rect 4090 -440 4190 -430
rect 4430 -440 11190 -340
rect 4430 -610 4890 -440
rect 5130 -610 5590 -440
rect 5830 -610 6290 -440
rect 6530 -610 6990 -440
rect 7230 -610 7690 -440
rect 7930 -610 8390 -440
rect 8630 -610 9090 -440
rect 9330 -610 9790 -440
rect 10030 -610 10490 -440
rect 10730 -610 11190 -440
rect 10910 -850 11010 -610
rect 4430 -1040 4890 -850
rect 5130 -1040 5590 -850
rect 5830 -1040 6290 -850
rect 6530 -1040 6990 -850
rect 7230 -1040 7690 -850
rect 7930 -1040 8390 -850
rect 8630 -1040 9090 -850
rect 9330 -1040 9790 -850
rect 10030 -1040 10490 -850
rect 10730 -1040 11190 -850
rect 4430 -1050 11190 -1040
rect 4230 -1060 11190 -1050
rect 4230 -1120 4240 -1060
rect 4300 -1120 11190 -1060
rect 4230 -1130 11190 -1120
rect 4430 -1140 11190 -1130
rect 4430 -1310 4890 -1140
rect 5130 -1310 5590 -1140
rect 5830 -1310 6290 -1140
rect 6530 -1310 6990 -1140
rect 7230 -1310 7690 -1140
rect 7930 -1310 8390 -1140
rect 8630 -1310 9090 -1140
rect 9330 -1310 9790 -1140
rect 10030 -1310 10490 -1140
rect 10730 -1310 11190 -1140
rect 4430 -1740 4890 -1550
rect 5130 -1740 5590 -1550
rect 5830 -1740 6290 -1550
rect 6530 -1740 6990 -1550
rect 7230 -1740 7690 -1550
rect 7930 -1740 8390 -1550
rect 8630 -1740 9090 -1550
rect 9330 -1740 9790 -1550
rect 10030 -1740 10490 -1550
rect 10730 -1740 11190 -1550
rect 3970 -1750 4070 -1740
rect 3970 -1830 3980 -1750
rect 4060 -1830 4070 -1750
rect 3970 -1840 4070 -1830
rect 4430 -1840 11190 -1740
rect 4430 -2010 4890 -1840
rect 5130 -2010 5590 -1840
rect 5830 -2010 6290 -1840
rect 6530 -2010 6990 -1840
rect 7230 -2010 7690 -1840
rect 7930 -2010 8390 -1840
rect 8630 -2010 9090 -1840
rect 9330 -2010 9790 -1840
rect 10030 -2010 10490 -1840
rect 10730 -2010 11190 -1840
rect 10910 -2250 11010 -2010
rect 4430 -2440 4890 -2250
rect 5130 -2440 5590 -2250
rect 5830 -2440 6290 -2250
rect 6530 -2440 6990 -2250
rect 7230 -2440 7690 -2250
rect 7930 -2440 8390 -2250
rect 8630 -2440 9090 -2250
rect 9330 -2440 9790 -2250
rect 10030 -2440 10490 -2250
rect 10730 -2440 11190 -2250
rect 4430 -2450 11190 -2440
rect 4300 -2460 11190 -2450
rect 4300 -2520 4310 -2460
rect 4370 -2520 11190 -2460
rect 4300 -2530 11190 -2520
rect 4430 -2540 11190 -2530
rect 4430 -2710 4890 -2540
rect 5130 -2710 5590 -2540
rect 5830 -2710 6290 -2540
rect 6530 -2710 6990 -2540
rect 7230 -2710 7690 -2540
rect 7930 -2710 8390 -2540
rect 8630 -2710 9090 -2540
rect 9330 -2710 9790 -2540
rect 10030 -2710 10490 -2540
rect 10730 -2710 11190 -2540
rect -3070 -2910 -2970 -2890
rect -3070 -2970 -3050 -2910
rect -2990 -2970 -2970 -2910
rect -3070 -3620 -2970 -2970
rect 14000 -2910 14100 -2890
rect 14000 -2970 14020 -2910
rect 14080 -2970 14100 -2910
rect 10810 -3290 10920 -3270
rect 10810 -3360 10830 -3290
rect 10900 -3360 10920 -3290
rect 10810 -3380 10920 -3360
rect 11310 -3290 11420 -3270
rect 11310 -3360 11330 -3290
rect 11400 -3360 11420 -3290
rect 11310 -3380 11420 -3360
rect 14000 -3620 14100 -2970
rect -3070 -15680 10950 -3620
rect 11280 -15680 14100 -3620
<< via3 >>
rect 8870 9270 8940 9340
rect 8870 8740 8940 8810
rect 9570 5260 9640 5330
rect 9570 4750 9640 4820
rect 4100 1040 4180 1050
rect 4100 980 4110 1040
rect 4110 980 4170 1040
rect 4170 980 4180 1040
rect 4100 970 4180 980
rect 4100 -360 4180 -350
rect 4100 -420 4110 -360
rect 4110 -420 4170 -360
rect 4170 -420 4180 -360
rect 4100 -430 4180 -420
rect 3980 -1760 4060 -1750
rect 3980 -1820 3990 -1760
rect 3990 -1820 4050 -1760
rect 4050 -1820 4060 -1760
rect 3980 -1830 4060 -1820
rect 10830 -3360 10900 -3290
rect 11330 -3360 11400 -3290
<< mimcap >>
rect 9230 9340 10270 10510
rect 9230 9270 9250 9340
rect 9320 9270 10270 9340
rect 9230 9250 10270 9270
rect 9230 8810 9770 8830
rect 9230 8740 9250 8810
rect 9320 8740 9770 8810
rect 9230 8070 9770 8740
rect 9930 5330 11930 7240
rect 9930 5260 9950 5330
rect 10020 5260 11930 5330
rect 9930 5240 11930 5260
rect 9930 4820 11930 4840
rect 9930 4750 9950 4820
rect 10020 4750 11930 4820
rect 9930 2840 11930 4750
rect 4460 1050 4860 1220
rect 4460 970 4630 1050
rect 4710 970 4860 1050
rect 4460 820 4860 970
rect 5160 1050 5560 1220
rect 5160 970 5320 1050
rect 5400 970 5560 1050
rect 5160 820 5560 970
rect 5860 1050 6260 1220
rect 5860 970 6020 1050
rect 6100 970 6260 1050
rect 5860 820 6260 970
rect 6560 1050 6960 1220
rect 6560 970 6720 1050
rect 6800 970 6960 1050
rect 6560 820 6960 970
rect 7260 1050 7660 1220
rect 7260 970 7420 1050
rect 7500 970 7660 1050
rect 7260 820 7660 970
rect 7960 1050 8360 1220
rect 7960 970 8120 1050
rect 8200 970 8360 1050
rect 7960 820 8360 970
rect 8660 1050 9060 1220
rect 8660 970 8820 1050
rect 8900 970 9060 1050
rect 8660 820 9060 970
rect 9360 1050 9760 1220
rect 9360 970 9520 1050
rect 9600 970 9760 1050
rect 9360 820 9760 970
rect 10060 1050 10460 1220
rect 10060 970 10220 1050
rect 10300 970 10460 1050
rect 10060 820 10460 970
rect 10760 1050 11160 1220
rect 10760 970 10920 1050
rect 11000 970 11160 1050
rect 10760 820 11160 970
rect 4460 350 4860 520
rect 4460 270 4630 350
rect 4710 270 4860 350
rect 4460 120 4860 270
rect 5160 350 5560 520
rect 5160 270 5320 350
rect 5400 270 5560 350
rect 5160 120 5560 270
rect 5860 350 6260 520
rect 5860 270 6020 350
rect 6100 270 6260 350
rect 5860 120 6260 270
rect 6560 350 6960 520
rect 6560 270 6720 350
rect 6800 270 6960 350
rect 6560 120 6960 270
rect 7260 350 7660 520
rect 7260 270 7420 350
rect 7500 270 7660 350
rect 7260 120 7660 270
rect 7960 350 8360 520
rect 7960 270 8120 350
rect 8200 270 8360 350
rect 7960 120 8360 270
rect 8660 350 9060 520
rect 8660 270 8820 350
rect 8900 270 9060 350
rect 8660 120 9060 270
rect 9360 350 9760 520
rect 9360 270 9520 350
rect 9600 270 9760 350
rect 9360 120 9760 270
rect 10060 350 10460 520
rect 10060 270 10220 350
rect 10300 270 10460 350
rect 10060 120 10460 270
rect 10760 350 11160 520
rect 10760 270 10920 350
rect 11000 270 11160 350
rect 10760 120 11160 270
rect 4460 -350 4860 -180
rect 4460 -430 4630 -350
rect 4710 -430 4860 -350
rect 4460 -580 4860 -430
rect 5160 -350 5560 -180
rect 5160 -430 5320 -350
rect 5400 -430 5560 -350
rect 5160 -580 5560 -430
rect 5860 -350 6260 -180
rect 5860 -430 6020 -350
rect 6100 -430 6260 -350
rect 5860 -580 6260 -430
rect 6560 -350 6960 -180
rect 6560 -430 6720 -350
rect 6800 -430 6960 -350
rect 6560 -580 6960 -430
rect 7260 -350 7660 -180
rect 7260 -430 7420 -350
rect 7500 -430 7660 -350
rect 7260 -580 7660 -430
rect 7960 -350 8360 -180
rect 7960 -430 8120 -350
rect 8200 -430 8360 -350
rect 7960 -580 8360 -430
rect 8660 -350 9060 -180
rect 8660 -430 8820 -350
rect 8900 -430 9060 -350
rect 8660 -580 9060 -430
rect 9360 -350 9760 -180
rect 9360 -430 9520 -350
rect 9600 -430 9760 -350
rect 9360 -580 9760 -430
rect 10060 -350 10460 -180
rect 10060 -430 10220 -350
rect 10300 -430 10460 -350
rect 10060 -580 10460 -430
rect 10760 -350 11160 -180
rect 10760 -430 10920 -350
rect 11000 -430 11160 -350
rect 10760 -580 11160 -430
rect 4460 -1050 4860 -880
rect 4460 -1130 4630 -1050
rect 4710 -1130 4860 -1050
rect 4460 -1280 4860 -1130
rect 5160 -1050 5560 -880
rect 5160 -1130 5320 -1050
rect 5400 -1130 5560 -1050
rect 5160 -1280 5560 -1130
rect 5860 -1050 6260 -880
rect 5860 -1130 6020 -1050
rect 6100 -1130 6260 -1050
rect 5860 -1280 6260 -1130
rect 6560 -1050 6960 -880
rect 6560 -1130 6720 -1050
rect 6800 -1130 6960 -1050
rect 6560 -1280 6960 -1130
rect 7260 -1050 7660 -880
rect 7260 -1130 7420 -1050
rect 7500 -1130 7660 -1050
rect 7260 -1280 7660 -1130
rect 7960 -1050 8360 -880
rect 7960 -1130 8120 -1050
rect 8200 -1130 8360 -1050
rect 7960 -1280 8360 -1130
rect 8660 -1050 9060 -880
rect 8660 -1130 8820 -1050
rect 8900 -1130 9060 -1050
rect 8660 -1280 9060 -1130
rect 9360 -1050 9760 -880
rect 9360 -1130 9520 -1050
rect 9600 -1130 9760 -1050
rect 9360 -1280 9760 -1130
rect 10060 -1050 10460 -880
rect 10060 -1130 10220 -1050
rect 10300 -1130 10460 -1050
rect 10060 -1280 10460 -1130
rect 10760 -1050 11160 -880
rect 10760 -1130 10920 -1050
rect 11000 -1130 11160 -1050
rect 10760 -1280 11160 -1130
rect 4460 -1750 4860 -1580
rect 4460 -1830 4630 -1750
rect 4710 -1830 4860 -1750
rect 4460 -1980 4860 -1830
rect 5160 -1750 5560 -1580
rect 5160 -1830 5320 -1750
rect 5400 -1830 5560 -1750
rect 5160 -1980 5560 -1830
rect 5860 -1750 6260 -1580
rect 5860 -1830 6020 -1750
rect 6100 -1830 6260 -1750
rect 5860 -1980 6260 -1830
rect 6560 -1750 6960 -1580
rect 6560 -1830 6720 -1750
rect 6800 -1830 6960 -1750
rect 6560 -1980 6960 -1830
rect 7260 -1750 7660 -1580
rect 7260 -1830 7420 -1750
rect 7500 -1830 7660 -1750
rect 7260 -1980 7660 -1830
rect 7960 -1750 8360 -1580
rect 7960 -1830 8120 -1750
rect 8200 -1830 8360 -1750
rect 7960 -1980 8360 -1830
rect 8660 -1750 9060 -1580
rect 8660 -1830 8820 -1750
rect 8900 -1830 9060 -1750
rect 8660 -1980 9060 -1830
rect 9360 -1750 9760 -1580
rect 9360 -1830 9520 -1750
rect 9600 -1830 9760 -1750
rect 9360 -1980 9760 -1830
rect 10060 -1750 10460 -1580
rect 10060 -1830 10220 -1750
rect 10300 -1830 10460 -1750
rect 10060 -1980 10460 -1830
rect 10760 -1750 11160 -1580
rect 10760 -1830 10920 -1750
rect 11000 -1830 11160 -1750
rect 10760 -1980 11160 -1830
rect 4460 -2450 4860 -2280
rect 4460 -2530 4630 -2450
rect 4710 -2530 4860 -2450
rect 4460 -2680 4860 -2530
rect 5160 -2450 5560 -2280
rect 5160 -2530 5320 -2450
rect 5400 -2530 5560 -2450
rect 5160 -2680 5560 -2530
rect 5860 -2450 6260 -2280
rect 5860 -2530 6020 -2450
rect 6100 -2530 6260 -2450
rect 5860 -2680 6260 -2530
rect 6560 -2450 6960 -2280
rect 6560 -2530 6720 -2450
rect 6800 -2530 6960 -2450
rect 6560 -2680 6960 -2530
rect 7260 -2450 7660 -2280
rect 7260 -2530 7420 -2450
rect 7500 -2530 7660 -2450
rect 7260 -2680 7660 -2530
rect 7960 -2450 8360 -2280
rect 7960 -2530 8120 -2450
rect 8200 -2530 8360 -2450
rect 7960 -2680 8360 -2530
rect 8660 -2450 9060 -2280
rect 8660 -2530 8820 -2450
rect 8900 -2530 9060 -2450
rect 8660 -2680 9060 -2530
rect 9360 -2450 9760 -2280
rect 9360 -2530 9520 -2450
rect 9600 -2530 9760 -2450
rect 9360 -2680 9760 -2530
rect 10060 -2450 10460 -2280
rect 10060 -2530 10220 -2450
rect 10300 -2530 10460 -2450
rect 10060 -2680 10460 -2530
rect 10760 -2450 11160 -2280
rect 10760 -2530 10920 -2450
rect 11000 -2530 11160 -2450
rect 10760 -2680 11160 -2530
rect -3040 -3670 10920 -3650
rect -3040 -3740 10830 -3670
rect 10900 -3740 10920 -3670
rect -3040 -15650 10920 -3740
rect 11310 -3670 14070 -3650
rect 11310 -3740 11330 -3670
rect 11400 -3740 14070 -3670
rect 11310 -15650 14070 -3740
<< mimcapcontact >>
rect 9250 9270 9320 9340
rect 9250 8740 9320 8810
rect 9950 5260 10020 5330
rect 9950 4750 10020 4820
rect 4630 970 4710 1050
rect 5320 970 5400 1050
rect 6020 970 6100 1050
rect 6720 970 6800 1050
rect 7420 970 7500 1050
rect 8120 970 8200 1050
rect 8820 970 8900 1050
rect 9520 970 9600 1050
rect 10220 970 10300 1050
rect 10920 970 11000 1050
rect 4630 270 4710 350
rect 5320 270 5400 350
rect 6020 270 6100 350
rect 6720 270 6800 350
rect 7420 270 7500 350
rect 8120 270 8200 350
rect 8820 270 8900 350
rect 9520 270 9600 350
rect 10220 270 10300 350
rect 10920 270 11000 350
rect 4630 -430 4710 -350
rect 5320 -430 5400 -350
rect 6020 -430 6100 -350
rect 6720 -430 6800 -350
rect 7420 -430 7500 -350
rect 8120 -430 8200 -350
rect 8820 -430 8900 -350
rect 9520 -430 9600 -350
rect 10220 -430 10300 -350
rect 10920 -430 11000 -350
rect 4630 -1130 4710 -1050
rect 5320 -1130 5400 -1050
rect 6020 -1130 6100 -1050
rect 6720 -1130 6800 -1050
rect 7420 -1130 7500 -1050
rect 8120 -1130 8200 -1050
rect 8820 -1130 8900 -1050
rect 9520 -1130 9600 -1050
rect 10220 -1130 10300 -1050
rect 10920 -1130 11000 -1050
rect 4630 -1830 4710 -1750
rect 5320 -1830 5400 -1750
rect 6020 -1830 6100 -1750
rect 6720 -1830 6800 -1750
rect 7420 -1830 7500 -1750
rect 8120 -1830 8200 -1750
rect 8820 -1830 8900 -1750
rect 9520 -1830 9600 -1750
rect 10220 -1830 10300 -1750
rect 10920 -1830 11000 -1750
rect 4630 -2530 4710 -2450
rect 5320 -2530 5400 -2450
rect 6020 -2530 6100 -2450
rect 6720 -2530 6800 -2450
rect 7420 -2530 7500 -2450
rect 8120 -2530 8200 -2450
rect 8820 -2530 8900 -2450
rect 9520 -2530 9600 -2450
rect 10220 -2530 10300 -2450
rect 10920 -2530 11000 -2450
rect 10830 -3740 10900 -3670
rect 11330 -3740 11400 -3670
<< metal4 >>
rect 8850 9340 9340 9360
rect 8850 9270 8870 9340
rect 8940 9270 9250 9340
rect 9320 9270 9340 9340
rect 8850 9250 9340 9270
rect 8850 8810 9340 8830
rect 8850 8740 8870 8810
rect 8940 8740 9250 8810
rect 9320 8740 9340 8810
rect 8850 8720 9340 8740
rect 9550 5330 10030 5350
rect 9550 5260 9570 5330
rect 9640 5260 9950 5330
rect 10020 5260 10030 5330
rect 9550 5240 10030 5260
rect 9550 4820 10030 4840
rect 9550 4750 9570 4820
rect 9640 4750 9950 4820
rect 10020 4750 10030 4820
rect 9550 4730 10030 4750
rect 4090 1050 11010 1060
rect 4090 970 4100 1050
rect 4180 970 4630 1050
rect 4710 970 5320 1050
rect 5400 970 6020 1050
rect 6100 970 6720 1050
rect 6800 970 7420 1050
rect 7500 970 8120 1050
rect 8200 970 8820 1050
rect 8900 970 9520 1050
rect 9600 970 10220 1050
rect 10300 970 10920 1050
rect 11000 970 11010 1050
rect 4090 960 11010 970
rect 10910 360 11010 960
rect 4620 350 11010 360
rect 4620 270 4630 350
rect 4710 270 5320 350
rect 5400 270 6020 350
rect 6100 270 6720 350
rect 6800 270 7420 350
rect 7500 270 8120 350
rect 8200 270 8820 350
rect 8900 270 9520 350
rect 9600 270 10220 350
rect 10300 270 10920 350
rect 11000 270 11010 350
rect 4620 260 11010 270
rect 4090 -350 11010 -340
rect 4090 -430 4100 -350
rect 4180 -430 4630 -350
rect 4710 -430 5320 -350
rect 5400 -430 6020 -350
rect 6100 -430 6720 -350
rect 6800 -430 7420 -350
rect 7500 -430 8120 -350
rect 8200 -430 8820 -350
rect 8900 -430 9520 -350
rect 9600 -430 10220 -350
rect 10300 -430 10920 -350
rect 11000 -430 11010 -350
rect 4090 -440 11010 -430
rect 10910 -1040 11010 -440
rect 4620 -1050 11010 -1040
rect 4620 -1130 4630 -1050
rect 4710 -1130 5320 -1050
rect 5400 -1130 6020 -1050
rect 6100 -1130 6720 -1050
rect 6800 -1130 7420 -1050
rect 7500 -1130 8120 -1050
rect 8200 -1130 8820 -1050
rect 8900 -1130 9520 -1050
rect 9600 -1130 10220 -1050
rect 10300 -1130 10920 -1050
rect 11000 -1130 11010 -1050
rect 4620 -1140 11010 -1130
rect 3970 -1750 11010 -1740
rect 3970 -1830 3980 -1750
rect 4060 -1830 4630 -1750
rect 4710 -1830 5320 -1750
rect 5400 -1830 6020 -1750
rect 6100 -1830 6720 -1750
rect 6800 -1830 7420 -1750
rect 7500 -1830 8120 -1750
rect 8200 -1830 8820 -1750
rect 8900 -1830 9520 -1750
rect 9600 -1830 10220 -1750
rect 10300 -1830 10920 -1750
rect 11000 -1830 11010 -1750
rect 3970 -1840 11010 -1830
rect 10910 -2440 11010 -1840
rect 4620 -2450 11010 -2440
rect 4620 -2530 4630 -2450
rect 4710 -2530 5320 -2450
rect 5400 -2530 6020 -2450
rect 6100 -2530 6720 -2450
rect 6800 -2530 7420 -2450
rect 7500 -2530 8120 -2450
rect 8200 -2530 8820 -2450
rect 8900 -2530 9520 -2450
rect 9600 -2530 10220 -2450
rect 10300 -2530 10920 -2450
rect 11000 -2530 11010 -2450
rect 4620 -2540 11010 -2530
rect 10810 -3290 10920 -3270
rect 10810 -3360 10830 -3290
rect 10900 -3360 10920 -3290
rect 10810 -3670 10920 -3360
rect 10810 -3740 10830 -3670
rect 10900 -3740 10920 -3670
rect 10810 -3750 10920 -3740
rect 11310 -3290 11420 -3270
rect 11310 -3360 11330 -3290
rect 11400 -3360 11420 -3290
rect 11310 -3670 11420 -3360
rect 11310 -3740 11330 -3670
rect 11400 -3740 11420 -3670
rect 11310 -3750 11420 -3740
use sky130_fd_pr__res_xhigh_po_0p35_CKJJH6  sky130_fd_pr__res_xhigh_po_0p35_CKJJH6_0
timestamp 0
transform 1 0 9369 0 1 6204
box -262 -677 262 677
use sky130_fd_pr__res_xhigh_po_0p35_Y4K2XU  sky130_fd_pr__res_xhigh_po_0p35_Y4K2XU_0
timestamp 0
transform 1 0 9369 0 1 3712
box -262 -705 262 705
<< end >>
