magic
tech sky130A
magscale 1 2
timestamp 1756886911
<< nwell >>
rect 330 12730 10780 12940
rect 11060 10760 13370 12990
rect 1140 8620 6120 9860
rect 7400 9250 10620 9830
rect -480 6630 1160 6910
rect 1420 6630 3060 6910
rect -490 5630 3070 6310
rect 3370 5830 4140 6110
rect 11007 5527 11531 6881
rect -1590 4470 1140 4750
rect 1440 4470 4170 4750
rect 7310 3530 10750 4840
rect 11007 3007 11531 4417
rect -3763 -2303 -3239 -711
rect -2976 -2306 -2120 -312
rect -1863 -2303 -1007 219
rect 3457 -2303 4313 219
rect 4570 -2300 5094 -918
rect 5357 -2303 5881 -711
rect 2827 -3403 5513 -2879
<< pwell >>
rect 11060 13070 13180 14490
rect -740 1427 600 1580
rect -740 393 -587 1427
rect 447 393 600 1427
rect -740 240 600 393
rect 620 1427 1960 1580
rect 620 393 773 1427
rect 1807 393 1960 1427
rect 620 240 1960 393
rect 1980 1427 3320 1580
rect 1980 393 2133 1427
rect 3167 393 3320 1427
rect 1980 240 3320 393
rect -740 67 600 220
rect -740 -967 -587 67
rect 447 -967 600 67
rect -740 -1120 600 -967
rect 620 67 1960 220
rect 620 -967 773 67
rect 1807 -967 1960 67
rect 620 -1120 1960 -967
rect 1980 67 3320 220
rect 1980 -967 2133 67
rect 3167 -967 3320 67
rect 1980 -1120 3320 -967
rect -740 -1293 600 -1140
rect -740 -2327 -587 -1293
rect 447 -2327 600 -1293
rect -740 -2480 600 -2327
rect 620 -1293 1960 -1140
rect 620 -2327 773 -1293
rect 1807 -2327 1960 -1293
rect 620 -2480 1960 -2327
rect 1980 -1293 3320 -1140
rect 1980 -2327 2133 -1293
rect 3167 -2327 3320 -1293
rect 1980 -2480 3320 -2327
rect 1250 -2760 1330 -2480
<< nbase >>
rect -587 393 447 1427
rect 773 393 1807 1427
rect 2133 393 3167 1427
rect -587 -967 447 67
rect 773 -967 1807 67
rect 2133 -967 3167 67
rect -587 -2327 447 -1293
rect 773 -2327 1807 -1293
rect 2133 -2327 3167 -1293
<< nmos >>
rect 11290 14150 11320 14350
rect 11810 14150 11840 14350
rect 12330 14150 12360 14350
rect 12930 14150 12960 14350
rect 11290 13670 11320 13970
rect 11810 13670 11840 13970
rect 12330 13670 12360 13970
rect 520 13120 550 13220
rect 630 13120 660 13220
rect 740 13120 770 13220
rect 850 13120 880 13220
rect 1100 13120 1130 13220
rect 1210 13120 1240 13220
rect 1550 13120 1580 13220
rect 1660 13120 1690 13220
rect 1770 13120 1800 13220
rect 1880 13120 1910 13220
rect 2210 13120 2240 13220
rect 2320 13120 2350 13220
rect 2430 13120 2460 13220
rect 2540 13120 2570 13220
rect 2890 13120 2920 13220
rect 3000 13120 3030 13220
rect 3110 13120 3140 13220
rect 3220 13120 3250 13220
rect 3470 13120 3500 13220
rect 3580 13120 3610 13220
rect 4030 13120 4060 13220
rect 4390 13120 4420 13220
rect 4640 13120 4670 13220
rect 4750 13120 4780 13220
rect 4860 13120 4890 13220
rect 4970 13120 5000 13220
rect 5300 13120 5330 13220
rect 5410 13120 5440 13220
rect 5520 13120 5550 13220
rect 5850 13120 5880 13220
rect 5960 13120 5990 13220
rect 6070 13120 6100 13220
rect 6180 13120 6210 13220
rect 6510 13120 6540 13220
rect 6620 13120 6650 13220
rect 6730 13120 6760 13220
rect 7150 13210 7180 13310
rect 7260 13210 7290 13310
rect 7370 13210 7400 13310
rect 7480 13210 7510 13310
rect 7810 13210 7840 13310
rect 7920 13210 7950 13310
rect 8030 13210 8060 13310
rect 8450 13210 8480 13310
rect 8560 13210 8590 13310
rect 8670 13210 8700 13310
rect 8780 13210 8810 13310
rect 9110 13210 9140 13310
rect 9220 13210 9250 13310
rect 9330 13210 9360 13310
rect 9750 13210 9780 13310
rect 9860 13210 9890 13310
rect 9970 13210 10000 13310
rect 10080 13210 10110 13310
rect 10410 13210 10440 13310
rect 10520 13210 10550 13310
rect 10630 13210 10660 13310
rect 11288 13290 11320 13490
rect 11808 13290 11840 13490
rect 12328 13290 12360 13490
rect 1340 10040 1370 10240
rect 1450 10040 1480 10240
rect 1860 10040 1890 10240
rect 1970 10040 2000 10240
rect 2240 10040 2270 10240
rect 2350 10040 2380 10240
rect 2760 10040 2790 10240
rect 2870 10040 2900 10240
rect 3280 10040 3310 10240
rect 3390 10040 3420 10240
rect 3720 10040 3750 10240
rect 4050 10040 4080 10240
rect 4490 10040 4520 10240
rect 4880 10040 4910 10240
rect 5270 10040 5300 10240
rect 5560 10040 5590 10240
rect 1340 8240 1370 8440
rect 1450 8240 1480 8440
rect 1860 8240 1890 8440
rect 1970 8240 2000 8440
rect 2240 8240 2270 8440
rect 2350 8240 2380 8440
rect 2760 8240 2790 8440
rect 2870 8240 2900 8440
rect 3270 8240 3300 8440
rect 3600 8240 3630 8440
rect 3930 8240 3960 8440
rect 4490 8240 4520 8440
rect 4880 8240 4910 8440
rect 5270 8240 5300 8440
rect 5560 8240 5590 8440
rect 5950 8240 5980 8440
rect 7440 8290 7560 8690
rect 7660 8290 7780 8690
rect 7880 8290 8000 8690
rect 8100 8290 8220 8690
rect 8520 8290 8640 8690
rect 8740 8290 8860 8690
rect 8960 8290 9080 8690
rect 9180 8290 9300 8690
rect 9600 8290 9720 8690
rect 9820 8290 9940 8690
rect 10040 8290 10160 8690
rect 10260 8290 10380 8690
rect 7500 5810 7600 6060
rect 7700 5810 7800 6060
rect 7900 5810 8000 6060
rect 8100 5810 8200 6060
rect 8300 5810 8400 6060
rect 8500 5810 8600 6060
rect 8700 5810 8800 6060
rect 8900 5810 9000 6060
rect 9100 5810 9200 6060
rect 9300 5810 9400 6060
rect 7550 5270 7580 5370
rect 7680 5270 7710 5370
rect 7810 5270 7840 5370
rect 7940 5270 7970 5370
rect 8070 5270 8100 5370
rect 8200 5270 8230 5370
rect 8690 5270 8720 5370
rect 8820 5270 8850 5370
rect 8950 5270 8980 5370
rect 9080 5270 9110 5370
rect 9210 5270 9240 5370
rect 9340 5270 9370 5370
rect 9830 5270 9860 5370
rect 9960 5270 9990 5370
rect 10090 5270 10120 5370
rect 10220 5270 10250 5370
rect 10350 5270 10380 5370
rect 10480 5270 10510 5370
rect -550 3670 -510 3770
rect -430 3670 -390 3770
rect -310 3670 -270 3770
rect -190 3670 -150 3770
rect -70 3670 -30 3770
rect 50 3670 90 3770
rect 170 3670 210 3770
rect 290 3670 330 3770
rect 410 3670 450 3770
rect 530 3670 570 3770
rect 2010 3670 2050 3770
rect 2130 3670 2170 3770
rect 2250 3670 2290 3770
rect 2370 3670 2410 3770
rect 2490 3670 2530 3770
rect 2610 3670 2650 3770
rect 2730 3670 2770 3770
rect 2850 3670 2890 3770
rect 2970 3670 3010 3770
rect 3090 3670 3130 3770
rect -1170 2660 -170 3160
rect 70 2660 1070 3160
rect 1510 2660 2510 3160
rect 2750 2660 3750 3160
rect -750 2050 1250 2250
rect 1330 2050 3330 2250
<< pmos >>
rect 680 12800 710 12900
rect 1100 12800 1130 12900
rect 1210 12800 1240 12900
rect 1770 12800 1800 12900
rect 1880 12800 1910 12900
rect 2210 12800 2240 12900
rect 2320 12800 2350 12900
rect 2430 12800 2460 12900
rect 3050 12800 3080 12900
rect 3470 12800 3500 12900
rect 3580 12800 3610 12900
rect 3920 12800 3950 12900
rect 4030 12800 4060 12900
rect 4280 12800 4310 12900
rect 4390 12800 4420 12900
rect 4860 12800 4890 12900
rect 4970 12800 5000 12900
rect 5300 12800 5330 12900
rect 5410 12800 5440 12900
rect 5920 12800 5950 12900
rect 6260 12800 6290 12900
rect 6370 12800 6400 12900
rect 6620 12800 6650 12900
rect 6730 12800 6760 12900
rect 7220 12800 7250 12900
rect 7560 12800 7590 12900
rect 7670 12800 7700 12900
rect 7920 12800 7950 12900
rect 8030 12800 8060 12900
rect 8520 12800 8550 12900
rect 8860 12800 8890 12900
rect 8970 12800 9000 12900
rect 9220 12800 9250 12900
rect 9330 12800 9360 12900
rect 9820 12800 9850 12900
rect 10160 12800 10190 12900
rect 10270 12800 10300 12900
rect 10520 12800 10550 12900
rect 10630 12800 10660 12900
rect 11288 12370 11320 12770
rect 11808 12370 11840 12770
rect 12328 12370 12360 12770
rect 11290 11590 11320 12190
rect 11810 11590 11840 12190
rect 12330 11590 12360 12190
rect 11290 10900 11590 11300
rect 11810 10900 12110 11300
rect 12330 10900 12630 11300
rect 12850 10900 13150 11300
rect 1340 9420 1370 9820
rect 1450 9420 1480 9820
rect 1860 9420 1890 9820
rect 1970 9420 2000 9820
rect 2240 9420 2270 9820
rect 2350 9420 2380 9820
rect 2760 9420 2790 9820
rect 2870 9420 2900 9820
rect 3280 9420 3310 9820
rect 3390 9420 3420 9820
rect 3720 9420 3750 9820
rect 4050 9420 4080 9820
rect 4490 9420 4520 9820
rect 4880 9420 4910 9820
rect 5270 9420 5300 9820
rect 5560 9420 5590 9820
rect 5950 9420 5980 9820
rect 7640 9390 7760 9790
rect 7860 9390 7980 9790
rect 8080 9390 8200 9790
rect 8300 9390 8420 9790
rect 8520 9390 8640 9790
rect 8740 9390 8860 9790
rect 9160 9390 9280 9790
rect 9380 9390 9500 9790
rect 9600 9390 9720 9790
rect 9820 9390 9940 9790
rect 10040 9390 10160 9790
rect 10260 9390 10380 9790
rect 1340 8660 1370 9060
rect 1450 8660 1480 9060
rect 1860 8660 1890 9060
rect 1970 8660 2000 9060
rect 2240 8660 2270 9060
rect 2350 8660 2380 9060
rect 2760 8660 2790 9060
rect 2870 8660 2900 9060
rect 3270 8660 3300 9060
rect 3600 8660 3630 9060
rect 3930 8660 3960 9060
rect 4490 8660 4520 9060
rect 4880 8660 4910 9060
rect 5270 8660 5300 9060
rect 5560 8660 5590 9060
rect -280 6670 -250 6870
rect -170 6670 -140 6870
rect -60 6670 -30 6870
rect 50 6670 80 6870
rect 160 6670 190 6870
rect 270 6670 300 6870
rect 380 6670 410 6870
rect 490 6670 520 6870
rect 600 6670 630 6870
rect 710 6670 740 6870
rect 820 6670 850 6870
rect 930 6670 960 6870
rect 1620 6670 1650 6870
rect 1730 6670 1760 6870
rect 1840 6670 1870 6870
rect 1950 6670 1980 6870
rect 2060 6670 2090 6870
rect 2170 6670 2200 6870
rect 2280 6670 2310 6870
rect 2390 6670 2420 6870
rect 2500 6670 2530 6870
rect 2610 6670 2640 6870
rect 2720 6670 2750 6870
rect 2830 6670 2860 6870
rect -290 5670 -190 6270
rect -110 5670 -10 6270
rect 70 5670 170 6270
rect 250 5670 350 6270
rect 430 5670 530 6270
rect 610 5670 710 6270
rect 790 5670 890 6270
rect 970 5670 1070 6270
rect 1150 5670 1250 6270
rect 1330 5670 1430 6270
rect 1510 5670 1610 6270
rect 1690 5670 1790 6270
rect 1870 5670 1970 6270
rect 2050 5670 2150 6270
rect 2230 5670 2330 6270
rect 2410 5670 2510 6270
rect 2590 5670 2690 6270
rect 2770 5670 2870 6270
rect 3580 5870 3610 6070
rect 3690 5870 3720 6070
rect 3800 5870 3830 6070
rect 3910 5870 3940 6070
rect -1390 4510 -1350 4710
rect -1270 4510 -1230 4710
rect -1150 4510 -1110 4710
rect -1030 4510 -990 4710
rect -910 4510 -870 4710
rect -790 4510 -750 4710
rect -670 4510 -630 4710
rect -550 4510 -510 4710
rect -430 4510 -390 4710
rect -310 4510 -270 4710
rect -190 4510 -150 4710
rect -70 4510 -30 4710
rect 50 4510 90 4710
rect 170 4510 210 4710
rect 290 4510 330 4710
rect 410 4510 450 4710
rect 530 4510 570 4710
rect 650 4510 690 4710
rect 770 4510 810 4710
rect 890 4510 930 4710
rect 1650 4510 1690 4710
rect 1770 4510 1810 4710
rect 1890 4510 1930 4710
rect 2010 4510 2050 4710
rect 2130 4510 2170 4710
rect 2250 4510 2290 4710
rect 2370 4510 2410 4710
rect 2490 4510 2530 4710
rect 2610 4510 2650 4710
rect 2730 4510 2770 4710
rect 2850 4510 2890 4710
rect 2970 4510 3010 4710
rect 3090 4510 3130 4710
rect 3210 4510 3250 4710
rect 3330 4510 3370 4710
rect 3450 4510 3490 4710
rect 3570 4510 3610 4710
rect 3690 4510 3730 4710
rect 3810 4510 3850 4710
rect 3930 4510 3970 4710
rect 7550 4590 7580 4790
rect 7680 4590 7710 4790
rect 7810 4590 7840 4790
rect 7940 4590 7970 4790
rect 8070 4590 8100 4790
rect 8200 4590 8230 4790
rect 8690 4590 8720 4790
rect 8820 4590 8850 4790
rect 8950 4590 8980 4790
rect 9080 4590 9110 4790
rect 9210 4590 9240 4790
rect 9340 4590 9370 4790
rect 9830 4590 9860 4790
rect 9960 4590 9990 4790
rect 10090 4590 10120 4790
rect 10220 4590 10250 4790
rect 10350 4590 10380 4790
rect 10480 4590 10510 4790
rect 7620 3640 7720 4140
rect 7820 3640 7920 4140
rect 8020 3640 8120 4140
rect 8220 3640 8320 4140
rect 8420 3640 8520 4140
rect 8620 3640 8720 4140
rect 8820 3640 8920 4140
rect 9020 3640 9120 4140
rect 9220 3640 9320 4140
rect 9420 3640 9520 4140
<< ndiff >>
rect 11210 14320 11290 14350
rect 11210 14280 11230 14320
rect 11270 14280 11290 14320
rect 11210 14220 11290 14280
rect 11210 14180 11230 14220
rect 11270 14180 11290 14220
rect 11210 14150 11290 14180
rect 11320 14320 11400 14350
rect 11320 14280 11340 14320
rect 11380 14280 11400 14320
rect 11320 14220 11400 14280
rect 11320 14180 11340 14220
rect 11380 14180 11400 14220
rect 11320 14150 11400 14180
rect 11730 14320 11810 14350
rect 11730 14280 11750 14320
rect 11790 14280 11810 14320
rect 11730 14220 11810 14280
rect 11730 14180 11750 14220
rect 11790 14180 11810 14220
rect 11730 14150 11810 14180
rect 11840 14320 11920 14350
rect 11840 14280 11860 14320
rect 11900 14280 11920 14320
rect 11840 14220 11920 14280
rect 11840 14180 11860 14220
rect 11900 14180 11920 14220
rect 11840 14150 11920 14180
rect 12250 14320 12330 14350
rect 12250 14280 12270 14320
rect 12310 14280 12330 14320
rect 12250 14220 12330 14280
rect 12250 14180 12270 14220
rect 12310 14180 12330 14220
rect 12250 14150 12330 14180
rect 12360 14320 12440 14350
rect 12360 14280 12380 14320
rect 12420 14280 12440 14320
rect 12360 14220 12440 14280
rect 12360 14180 12380 14220
rect 12420 14180 12440 14220
rect 12360 14150 12440 14180
rect 12850 14320 12930 14350
rect 12850 14280 12870 14320
rect 12910 14280 12930 14320
rect 12850 14220 12930 14280
rect 12850 14180 12870 14220
rect 12910 14180 12930 14220
rect 12850 14150 12930 14180
rect 12960 14320 13040 14350
rect 12960 14280 12980 14320
rect 13020 14280 13040 14320
rect 12960 14220 13040 14280
rect 12960 14180 12980 14220
rect 13020 14180 13040 14220
rect 12960 14150 13040 14180
rect 11210 13940 11290 13970
rect 11210 13900 11230 13940
rect 11270 13900 11290 13940
rect 11210 13840 11290 13900
rect 11210 13800 11230 13840
rect 11270 13800 11290 13840
rect 11210 13740 11290 13800
rect 11210 13700 11230 13740
rect 11270 13700 11290 13740
rect 11210 13670 11290 13700
rect 11320 13940 11400 13970
rect 11320 13900 11340 13940
rect 11380 13900 11400 13940
rect 11320 13840 11400 13900
rect 11320 13800 11340 13840
rect 11380 13800 11400 13840
rect 11320 13740 11400 13800
rect 11320 13700 11340 13740
rect 11380 13700 11400 13740
rect 11320 13670 11400 13700
rect 11730 13940 11810 13970
rect 11730 13900 11750 13940
rect 11790 13900 11810 13940
rect 11730 13840 11810 13900
rect 11730 13800 11750 13840
rect 11790 13800 11810 13840
rect 11730 13740 11810 13800
rect 11730 13700 11750 13740
rect 11790 13700 11810 13740
rect 11730 13670 11810 13700
rect 11840 13940 11920 13970
rect 11840 13900 11860 13940
rect 11900 13900 11920 13940
rect 11840 13840 11920 13900
rect 11840 13800 11860 13840
rect 11900 13800 11920 13840
rect 11840 13740 11920 13800
rect 11840 13700 11860 13740
rect 11900 13700 11920 13740
rect 11840 13670 11920 13700
rect 12250 13940 12330 13970
rect 12250 13900 12270 13940
rect 12310 13900 12330 13940
rect 12250 13840 12330 13900
rect 12250 13800 12270 13840
rect 12310 13800 12330 13840
rect 12250 13740 12330 13800
rect 12250 13700 12270 13740
rect 12310 13700 12330 13740
rect 12250 13670 12330 13700
rect 12360 13940 12440 13970
rect 12360 13900 12380 13940
rect 12420 13900 12440 13940
rect 12360 13840 12440 13900
rect 12360 13800 12380 13840
rect 12420 13800 12440 13840
rect 12360 13740 12440 13800
rect 12360 13700 12380 13740
rect 12420 13700 12440 13740
rect 12360 13670 12440 13700
rect 440 13190 520 13220
rect 440 13150 460 13190
rect 500 13150 520 13190
rect 440 13120 520 13150
rect 550 13190 630 13220
rect 550 13150 570 13190
rect 610 13150 630 13190
rect 550 13120 630 13150
rect 660 13190 740 13220
rect 660 13150 680 13190
rect 720 13150 740 13190
rect 660 13120 740 13150
rect 770 13190 850 13220
rect 770 13150 790 13190
rect 830 13150 850 13190
rect 770 13120 850 13150
rect 880 13190 960 13220
rect 880 13150 900 13190
rect 940 13150 960 13190
rect 880 13120 960 13150
rect 1020 13190 1100 13220
rect 1020 13150 1040 13190
rect 1080 13150 1100 13190
rect 1020 13120 1100 13150
rect 1130 13190 1210 13220
rect 1130 13150 1150 13190
rect 1190 13150 1210 13190
rect 1130 13120 1210 13150
rect 1240 13190 1320 13220
rect 1240 13150 1260 13190
rect 1300 13150 1320 13190
rect 1240 13120 1320 13150
rect 1470 13190 1550 13220
rect 1470 13150 1490 13190
rect 1530 13150 1550 13190
rect 1470 13120 1550 13150
rect 1580 13190 1660 13220
rect 1580 13150 1600 13190
rect 1640 13150 1660 13190
rect 1580 13120 1660 13150
rect 1690 13190 1770 13220
rect 1690 13150 1710 13190
rect 1750 13150 1770 13190
rect 1690 13120 1770 13150
rect 1800 13190 1880 13220
rect 1800 13150 1820 13190
rect 1860 13150 1880 13190
rect 1800 13120 1880 13150
rect 1910 13190 1990 13220
rect 1910 13150 1930 13190
rect 1970 13150 1990 13190
rect 1910 13120 1990 13150
rect 2130 13190 2210 13220
rect 2130 13150 2150 13190
rect 2190 13150 2210 13190
rect 2130 13120 2210 13150
rect 2240 13190 2320 13220
rect 2240 13150 2260 13190
rect 2300 13150 2320 13190
rect 2240 13120 2320 13150
rect 2350 13190 2430 13220
rect 2350 13150 2370 13190
rect 2410 13150 2430 13190
rect 2350 13120 2430 13150
rect 2460 13190 2540 13220
rect 2460 13150 2480 13190
rect 2520 13150 2540 13190
rect 2460 13120 2540 13150
rect 2570 13190 2650 13220
rect 2570 13150 2590 13190
rect 2630 13150 2650 13190
rect 2570 13120 2650 13150
rect 2810 13190 2890 13220
rect 2810 13150 2830 13190
rect 2870 13150 2890 13190
rect 2810 13120 2890 13150
rect 2920 13190 3000 13220
rect 2920 13150 2940 13190
rect 2980 13150 3000 13190
rect 2920 13120 3000 13150
rect 3030 13190 3110 13220
rect 3030 13150 3050 13190
rect 3090 13150 3110 13190
rect 3030 13120 3110 13150
rect 3140 13190 3220 13220
rect 3140 13150 3160 13190
rect 3200 13150 3220 13190
rect 3140 13120 3220 13150
rect 3250 13190 3330 13220
rect 3250 13150 3270 13190
rect 3310 13150 3330 13190
rect 3250 13120 3330 13150
rect 3390 13190 3470 13220
rect 3390 13150 3410 13190
rect 3450 13150 3470 13190
rect 3390 13120 3470 13150
rect 3500 13190 3580 13220
rect 3500 13150 3520 13190
rect 3560 13150 3580 13190
rect 3500 13120 3580 13150
rect 3610 13190 3690 13220
rect 3610 13150 3630 13190
rect 3670 13150 3690 13190
rect 3610 13120 3690 13150
rect 3950 13190 4030 13220
rect 3950 13150 3970 13190
rect 4010 13150 4030 13190
rect 3950 13120 4030 13150
rect 4060 13190 4140 13220
rect 4060 13150 4080 13190
rect 4120 13150 4140 13190
rect 4060 13120 4140 13150
rect 4310 13190 4390 13220
rect 4310 13150 4330 13190
rect 4370 13150 4390 13190
rect 4310 13120 4390 13150
rect 4420 13190 4500 13220
rect 4420 13150 4440 13190
rect 4480 13150 4500 13190
rect 4420 13120 4500 13150
rect 4560 13190 4640 13220
rect 4560 13150 4580 13190
rect 4620 13150 4640 13190
rect 4560 13120 4640 13150
rect 4670 13190 4750 13220
rect 4670 13150 4690 13190
rect 4730 13150 4750 13190
rect 4670 13120 4750 13150
rect 4780 13190 4860 13220
rect 4780 13150 4800 13190
rect 4840 13150 4860 13190
rect 4780 13120 4860 13150
rect 4890 13190 4970 13220
rect 4890 13150 4910 13190
rect 4950 13150 4970 13190
rect 4890 13120 4970 13150
rect 5000 13190 5080 13220
rect 5000 13150 5020 13190
rect 5060 13150 5080 13190
rect 5000 13120 5080 13150
rect 5220 13190 5300 13220
rect 5220 13150 5240 13190
rect 5280 13150 5300 13190
rect 5220 13120 5300 13150
rect 5330 13190 5410 13220
rect 5330 13150 5350 13190
rect 5390 13150 5410 13190
rect 5330 13120 5410 13150
rect 5440 13190 5520 13220
rect 5440 13150 5460 13190
rect 5500 13150 5520 13190
rect 5440 13120 5520 13150
rect 5550 13190 5630 13220
rect 5550 13150 5570 13190
rect 5610 13150 5630 13190
rect 5550 13120 5630 13150
rect 5770 13190 5850 13220
rect 5770 13150 5790 13190
rect 5830 13150 5850 13190
rect 5770 13120 5850 13150
rect 5880 13190 5960 13220
rect 5880 13150 5900 13190
rect 5940 13150 5960 13190
rect 5880 13120 5960 13150
rect 5990 13190 6070 13220
rect 5990 13150 6010 13190
rect 6050 13150 6070 13190
rect 5990 13120 6070 13150
rect 6100 13190 6180 13220
rect 6100 13150 6120 13190
rect 6160 13150 6180 13190
rect 6100 13120 6180 13150
rect 6210 13190 6290 13220
rect 6210 13150 6230 13190
rect 6270 13150 6290 13190
rect 6210 13120 6290 13150
rect 6430 13190 6510 13220
rect 6430 13150 6450 13190
rect 6490 13150 6510 13190
rect 6430 13120 6510 13150
rect 6540 13190 6620 13220
rect 6540 13150 6560 13190
rect 6600 13150 6620 13190
rect 6540 13120 6620 13150
rect 6650 13190 6730 13220
rect 6650 13150 6670 13190
rect 6710 13150 6730 13190
rect 6650 13120 6730 13150
rect 6760 13190 6840 13220
rect 7070 13280 7150 13310
rect 7070 13240 7090 13280
rect 7130 13240 7150 13280
rect 7070 13210 7150 13240
rect 7180 13280 7260 13310
rect 7180 13240 7200 13280
rect 7240 13240 7260 13280
rect 7180 13210 7260 13240
rect 7290 13280 7370 13310
rect 7290 13240 7310 13280
rect 7350 13240 7370 13280
rect 7290 13210 7370 13240
rect 7400 13280 7480 13310
rect 7400 13240 7420 13280
rect 7460 13240 7480 13280
rect 7400 13210 7480 13240
rect 7510 13280 7590 13310
rect 7510 13240 7530 13280
rect 7570 13240 7590 13280
rect 7510 13210 7590 13240
rect 7730 13280 7810 13310
rect 7730 13240 7750 13280
rect 7790 13240 7810 13280
rect 7730 13210 7810 13240
rect 7840 13280 7920 13310
rect 7840 13240 7860 13280
rect 7900 13240 7920 13280
rect 7840 13210 7920 13240
rect 7950 13280 8030 13310
rect 7950 13240 7970 13280
rect 8010 13240 8030 13280
rect 7950 13210 8030 13240
rect 8060 13280 8140 13310
rect 8060 13240 8080 13280
rect 8120 13240 8140 13280
rect 8060 13210 8140 13240
rect 8370 13280 8450 13310
rect 8370 13240 8390 13280
rect 8430 13240 8450 13280
rect 8370 13210 8450 13240
rect 8480 13280 8560 13310
rect 8480 13240 8500 13280
rect 8540 13240 8560 13280
rect 8480 13210 8560 13240
rect 8590 13280 8670 13310
rect 8590 13240 8610 13280
rect 8650 13240 8670 13280
rect 8590 13210 8670 13240
rect 8700 13280 8780 13310
rect 8700 13240 8720 13280
rect 8760 13240 8780 13280
rect 8700 13210 8780 13240
rect 8810 13280 8890 13310
rect 8810 13240 8830 13280
rect 8870 13240 8890 13280
rect 8810 13210 8890 13240
rect 9030 13280 9110 13310
rect 9030 13240 9050 13280
rect 9090 13240 9110 13280
rect 9030 13210 9110 13240
rect 9140 13280 9220 13310
rect 9140 13240 9160 13280
rect 9200 13240 9220 13280
rect 9140 13210 9220 13240
rect 9250 13280 9330 13310
rect 9250 13240 9270 13280
rect 9310 13240 9330 13280
rect 9250 13210 9330 13240
rect 9360 13280 9440 13310
rect 9360 13240 9380 13280
rect 9420 13240 9440 13280
rect 9360 13210 9440 13240
rect 9670 13280 9750 13310
rect 9670 13240 9690 13280
rect 9730 13240 9750 13280
rect 9670 13210 9750 13240
rect 9780 13280 9860 13310
rect 9780 13240 9800 13280
rect 9840 13240 9860 13280
rect 9780 13210 9860 13240
rect 9890 13280 9970 13310
rect 9890 13240 9910 13280
rect 9950 13240 9970 13280
rect 9890 13210 9970 13240
rect 10000 13280 10080 13310
rect 10000 13240 10020 13280
rect 10060 13240 10080 13280
rect 10000 13210 10080 13240
rect 10110 13280 10190 13310
rect 10110 13240 10130 13280
rect 10170 13240 10190 13280
rect 10110 13210 10190 13240
rect 10330 13280 10410 13310
rect 10330 13240 10350 13280
rect 10390 13240 10410 13280
rect 10330 13210 10410 13240
rect 10440 13280 10520 13310
rect 10440 13240 10460 13280
rect 10500 13240 10520 13280
rect 10440 13210 10520 13240
rect 10550 13280 10630 13310
rect 10550 13240 10570 13280
rect 10610 13240 10630 13280
rect 10550 13210 10630 13240
rect 10660 13280 10740 13310
rect 10660 13240 10680 13280
rect 10720 13240 10740 13280
rect 10660 13210 10740 13240
rect 6760 13150 6780 13190
rect 6820 13150 6840 13190
rect 6760 13120 6840 13150
rect 11208 13460 11288 13490
rect 11208 13420 11228 13460
rect 11268 13420 11288 13460
rect 11208 13360 11288 13420
rect 11208 13320 11228 13360
rect 11268 13320 11288 13360
rect 11208 13290 11288 13320
rect 11320 13460 11400 13490
rect 11320 13420 11340 13460
rect 11380 13420 11400 13460
rect 11320 13360 11400 13420
rect 11320 13320 11340 13360
rect 11380 13320 11400 13360
rect 11320 13290 11400 13320
rect 11728 13460 11808 13490
rect 11728 13420 11748 13460
rect 11788 13420 11808 13460
rect 11728 13360 11808 13420
rect 11728 13320 11748 13360
rect 11788 13320 11808 13360
rect 11728 13290 11808 13320
rect 11840 13460 11920 13490
rect 11840 13420 11860 13460
rect 11900 13420 11920 13460
rect 11840 13360 11920 13420
rect 11840 13320 11860 13360
rect 11900 13320 11920 13360
rect 11840 13290 11920 13320
rect 12248 13460 12328 13490
rect 12248 13420 12268 13460
rect 12308 13420 12328 13460
rect 12248 13360 12328 13420
rect 12248 13320 12268 13360
rect 12308 13320 12328 13360
rect 12248 13290 12328 13320
rect 12360 13460 12440 13490
rect 12360 13420 12380 13460
rect 12420 13420 12440 13460
rect 12360 13360 12440 13420
rect 12360 13320 12380 13360
rect 12420 13320 12440 13360
rect 12360 13290 12440 13320
rect 1260 10210 1340 10240
rect 1260 10170 1280 10210
rect 1320 10170 1340 10210
rect 1260 10110 1340 10170
rect 1260 10070 1280 10110
rect 1320 10070 1340 10110
rect 1260 10040 1340 10070
rect 1370 10210 1450 10240
rect 1370 10170 1390 10210
rect 1430 10170 1450 10210
rect 1370 10110 1450 10170
rect 1370 10070 1390 10110
rect 1430 10070 1450 10110
rect 1370 10040 1450 10070
rect 1480 10210 1560 10240
rect 1480 10170 1500 10210
rect 1540 10170 1560 10210
rect 1480 10110 1560 10170
rect 1480 10070 1500 10110
rect 1540 10070 1560 10110
rect 1480 10040 1560 10070
rect 1780 10210 1860 10240
rect 1780 10170 1800 10210
rect 1840 10170 1860 10210
rect 1780 10110 1860 10170
rect 1780 10070 1800 10110
rect 1840 10070 1860 10110
rect 1780 10040 1860 10070
rect 1890 10210 1970 10240
rect 1890 10170 1910 10210
rect 1950 10170 1970 10210
rect 1890 10110 1970 10170
rect 1890 10070 1910 10110
rect 1950 10070 1970 10110
rect 1890 10040 1970 10070
rect 2000 10210 2080 10240
rect 2160 10210 2240 10240
rect 2000 10170 2020 10210
rect 2060 10170 2080 10210
rect 2160 10170 2180 10210
rect 2220 10170 2240 10210
rect 2000 10110 2080 10170
rect 2160 10110 2240 10170
rect 2000 10070 2020 10110
rect 2060 10070 2080 10110
rect 2160 10070 2180 10110
rect 2220 10070 2240 10110
rect 2000 10040 2080 10070
rect 2160 10040 2240 10070
rect 2270 10210 2350 10240
rect 2270 10170 2290 10210
rect 2330 10170 2350 10210
rect 2270 10110 2350 10170
rect 2270 10070 2290 10110
rect 2330 10070 2350 10110
rect 2270 10040 2350 10070
rect 2380 10210 2460 10240
rect 2380 10170 2400 10210
rect 2440 10170 2460 10210
rect 2380 10110 2460 10170
rect 2380 10070 2400 10110
rect 2440 10070 2460 10110
rect 2380 10040 2460 10070
rect 2680 10210 2760 10240
rect 2680 10170 2700 10210
rect 2740 10170 2760 10210
rect 2680 10110 2760 10170
rect 2680 10070 2700 10110
rect 2740 10070 2760 10110
rect 2680 10040 2760 10070
rect 2790 10210 2870 10240
rect 2790 10170 2810 10210
rect 2850 10170 2870 10210
rect 2790 10110 2870 10170
rect 2790 10070 2810 10110
rect 2850 10070 2870 10110
rect 2790 10040 2870 10070
rect 2900 10210 2980 10240
rect 2900 10170 2920 10210
rect 2960 10170 2980 10210
rect 2900 10110 2980 10170
rect 2900 10070 2920 10110
rect 2960 10070 2980 10110
rect 2900 10040 2980 10070
rect 3200 10210 3280 10240
rect 3200 10170 3220 10210
rect 3260 10170 3280 10210
rect 3200 10110 3280 10170
rect 3200 10070 3220 10110
rect 3260 10070 3280 10110
rect 3200 10040 3280 10070
rect 3310 10210 3390 10240
rect 3310 10170 3330 10210
rect 3370 10170 3390 10210
rect 3310 10110 3390 10170
rect 3310 10070 3330 10110
rect 3370 10070 3390 10110
rect 3310 10040 3390 10070
rect 3420 10210 3500 10240
rect 3420 10170 3440 10210
rect 3480 10170 3500 10210
rect 3420 10110 3500 10170
rect 3420 10070 3440 10110
rect 3480 10070 3500 10110
rect 3420 10040 3500 10070
rect 3640 10210 3720 10240
rect 3640 10170 3660 10210
rect 3700 10170 3720 10210
rect 3640 10110 3720 10170
rect 3640 10070 3660 10110
rect 3700 10070 3720 10110
rect 3640 10040 3720 10070
rect 3750 10210 3830 10240
rect 3750 10170 3770 10210
rect 3810 10170 3830 10210
rect 3750 10110 3830 10170
rect 3750 10070 3770 10110
rect 3810 10070 3830 10110
rect 3750 10040 3830 10070
rect 3970 10210 4050 10240
rect 3970 10170 3990 10210
rect 4030 10170 4050 10210
rect 3970 10110 4050 10170
rect 3970 10070 3990 10110
rect 4030 10070 4050 10110
rect 3970 10040 4050 10070
rect 4080 10210 4160 10240
rect 4080 10170 4100 10210
rect 4140 10170 4160 10210
rect 4080 10110 4160 10170
rect 4080 10070 4100 10110
rect 4140 10070 4160 10110
rect 4080 10040 4160 10070
rect 4390 10210 4490 10240
rect 4390 10170 4420 10210
rect 4460 10170 4490 10210
rect 4390 10110 4490 10170
rect 4390 10070 4420 10110
rect 4460 10070 4490 10110
rect 4390 10040 4490 10070
rect 4520 10210 4620 10240
rect 4520 10170 4550 10210
rect 4590 10170 4620 10210
rect 4520 10110 4620 10170
rect 4520 10070 4550 10110
rect 4590 10070 4620 10110
rect 4520 10040 4620 10070
rect 4780 10210 4880 10240
rect 4780 10170 4810 10210
rect 4850 10170 4880 10210
rect 4780 10110 4880 10170
rect 4780 10070 4810 10110
rect 4850 10070 4880 10110
rect 4780 10040 4880 10070
rect 4910 10210 5010 10240
rect 4910 10170 4940 10210
rect 4980 10170 5010 10210
rect 4910 10110 5010 10170
rect 4910 10070 4940 10110
rect 4980 10070 5010 10110
rect 4910 10040 5010 10070
rect 5170 10210 5270 10240
rect 5170 10170 5200 10210
rect 5240 10170 5270 10210
rect 5170 10110 5270 10170
rect 5170 10070 5200 10110
rect 5240 10070 5270 10110
rect 5170 10040 5270 10070
rect 5300 10210 5400 10240
rect 5300 10170 5330 10210
rect 5370 10170 5400 10210
rect 5300 10110 5400 10170
rect 5300 10070 5330 10110
rect 5370 10070 5400 10110
rect 5300 10040 5400 10070
rect 5460 10210 5560 10240
rect 5460 10170 5490 10210
rect 5530 10170 5560 10210
rect 5460 10110 5560 10170
rect 5460 10070 5490 10110
rect 5530 10070 5560 10110
rect 5460 10040 5560 10070
rect 5590 10210 5690 10240
rect 5590 10170 5620 10210
rect 5660 10170 5690 10210
rect 5590 10110 5690 10170
rect 5590 10070 5620 10110
rect 5660 10070 5690 10110
rect 5590 10040 5690 10070
rect 7340 8660 7440 8690
rect 7340 8620 7370 8660
rect 7410 8620 7440 8660
rect 7340 8560 7440 8620
rect 7340 8520 7370 8560
rect 7410 8520 7440 8560
rect 7340 8460 7440 8520
rect 1260 8410 1340 8440
rect 1260 8370 1280 8410
rect 1320 8370 1340 8410
rect 1260 8310 1340 8370
rect 1260 8270 1280 8310
rect 1320 8270 1340 8310
rect 1260 8240 1340 8270
rect 1370 8410 1450 8440
rect 1370 8370 1390 8410
rect 1430 8370 1450 8410
rect 1370 8310 1450 8370
rect 1370 8270 1390 8310
rect 1430 8270 1450 8310
rect 1370 8240 1450 8270
rect 1480 8410 1560 8440
rect 1480 8370 1500 8410
rect 1540 8370 1560 8410
rect 1480 8310 1560 8370
rect 1480 8270 1500 8310
rect 1540 8270 1560 8310
rect 1480 8240 1560 8270
rect 1780 8410 1860 8440
rect 1780 8370 1800 8410
rect 1840 8370 1860 8410
rect 1780 8310 1860 8370
rect 1780 8270 1800 8310
rect 1840 8270 1860 8310
rect 1780 8240 1860 8270
rect 1890 8410 1970 8440
rect 1890 8370 1910 8410
rect 1950 8370 1970 8410
rect 1890 8310 1970 8370
rect 1890 8270 1910 8310
rect 1950 8270 1970 8310
rect 1890 8240 1970 8270
rect 2000 8410 2080 8440
rect 2160 8410 2240 8440
rect 2000 8370 2020 8410
rect 2060 8370 2080 8410
rect 2160 8370 2180 8410
rect 2220 8370 2240 8410
rect 2000 8310 2080 8370
rect 2160 8310 2240 8370
rect 2000 8270 2020 8310
rect 2060 8270 2080 8310
rect 2160 8270 2180 8310
rect 2220 8270 2240 8310
rect 2000 8240 2080 8270
rect 2160 8240 2240 8270
rect 2270 8410 2350 8440
rect 2270 8370 2290 8410
rect 2330 8370 2350 8410
rect 2270 8310 2350 8370
rect 2270 8270 2290 8310
rect 2330 8270 2350 8310
rect 2270 8240 2350 8270
rect 2380 8410 2460 8440
rect 2380 8370 2400 8410
rect 2440 8370 2460 8410
rect 2380 8310 2460 8370
rect 2380 8270 2400 8310
rect 2440 8270 2460 8310
rect 2380 8240 2460 8270
rect 2680 8410 2760 8440
rect 2680 8370 2700 8410
rect 2740 8370 2760 8410
rect 2680 8310 2760 8370
rect 2680 8270 2700 8310
rect 2740 8270 2760 8310
rect 2680 8240 2760 8270
rect 2790 8410 2870 8440
rect 2790 8370 2810 8410
rect 2850 8370 2870 8410
rect 2790 8310 2870 8370
rect 2790 8270 2810 8310
rect 2850 8270 2870 8310
rect 2790 8240 2870 8270
rect 2900 8410 2980 8440
rect 2900 8370 2920 8410
rect 2960 8370 2980 8410
rect 2900 8310 2980 8370
rect 2900 8270 2920 8310
rect 2960 8270 2980 8310
rect 2900 8240 2980 8270
rect 3190 8410 3270 8440
rect 3190 8370 3210 8410
rect 3250 8370 3270 8410
rect 3190 8310 3270 8370
rect 3190 8270 3210 8310
rect 3250 8270 3270 8310
rect 3190 8240 3270 8270
rect 3300 8410 3380 8440
rect 3300 8370 3320 8410
rect 3360 8370 3380 8410
rect 3300 8310 3380 8370
rect 3300 8270 3320 8310
rect 3360 8270 3380 8310
rect 3300 8240 3380 8270
rect 3520 8410 3600 8440
rect 3520 8370 3540 8410
rect 3580 8370 3600 8410
rect 3520 8310 3600 8370
rect 3520 8270 3540 8310
rect 3580 8270 3600 8310
rect 3520 8240 3600 8270
rect 3630 8410 3710 8440
rect 3630 8370 3650 8410
rect 3690 8370 3710 8410
rect 3630 8310 3710 8370
rect 3630 8270 3650 8310
rect 3690 8270 3710 8310
rect 3630 8240 3710 8270
rect 3850 8410 3930 8440
rect 3850 8370 3870 8410
rect 3910 8370 3930 8410
rect 3850 8310 3930 8370
rect 3850 8270 3870 8310
rect 3910 8270 3930 8310
rect 3850 8240 3930 8270
rect 3960 8410 4040 8440
rect 3960 8370 3980 8410
rect 4020 8370 4040 8410
rect 3960 8310 4040 8370
rect 3960 8270 3980 8310
rect 4020 8270 4040 8310
rect 3960 8240 4040 8270
rect 4390 8410 4490 8440
rect 4390 8370 4420 8410
rect 4460 8370 4490 8410
rect 4390 8310 4490 8370
rect 4390 8270 4420 8310
rect 4460 8270 4490 8310
rect 4390 8240 4490 8270
rect 4520 8410 4620 8440
rect 4520 8370 4550 8410
rect 4590 8370 4620 8410
rect 4520 8310 4620 8370
rect 4520 8270 4550 8310
rect 4590 8270 4620 8310
rect 4520 8240 4620 8270
rect 4780 8410 4880 8440
rect 4780 8370 4810 8410
rect 4850 8370 4880 8410
rect 4780 8310 4880 8370
rect 4780 8270 4810 8310
rect 4850 8270 4880 8310
rect 4780 8240 4880 8270
rect 4910 8410 5010 8440
rect 4910 8370 4940 8410
rect 4980 8370 5010 8410
rect 4910 8310 5010 8370
rect 4910 8270 4940 8310
rect 4980 8270 5010 8310
rect 4910 8240 5010 8270
rect 5170 8410 5270 8440
rect 5170 8370 5200 8410
rect 5240 8370 5270 8410
rect 5170 8310 5270 8370
rect 5170 8270 5200 8310
rect 5240 8270 5270 8310
rect 5170 8240 5270 8270
rect 5300 8410 5400 8440
rect 5300 8370 5330 8410
rect 5370 8370 5400 8410
rect 5300 8310 5400 8370
rect 5300 8270 5330 8310
rect 5370 8270 5400 8310
rect 5300 8240 5400 8270
rect 5460 8410 5560 8440
rect 5460 8370 5490 8410
rect 5530 8370 5560 8410
rect 5460 8310 5560 8370
rect 5460 8270 5490 8310
rect 5530 8270 5560 8310
rect 5460 8240 5560 8270
rect 5590 8410 5690 8440
rect 5590 8370 5620 8410
rect 5660 8370 5690 8410
rect 5590 8310 5690 8370
rect 5590 8270 5620 8310
rect 5660 8270 5690 8310
rect 5590 8240 5690 8270
rect 5850 8410 5950 8440
rect 5850 8370 5880 8410
rect 5920 8370 5950 8410
rect 5850 8310 5950 8370
rect 5850 8270 5880 8310
rect 5920 8270 5950 8310
rect 5850 8240 5950 8270
rect 5980 8410 6080 8440
rect 5980 8370 6010 8410
rect 6050 8370 6080 8410
rect 5980 8310 6080 8370
rect 5980 8270 6010 8310
rect 6050 8270 6080 8310
rect 7340 8420 7370 8460
rect 7410 8420 7440 8460
rect 7340 8360 7440 8420
rect 7340 8320 7370 8360
rect 7410 8320 7440 8360
rect 7340 8290 7440 8320
rect 7560 8660 7660 8690
rect 7560 8620 7590 8660
rect 7630 8620 7660 8660
rect 7560 8560 7660 8620
rect 7560 8520 7590 8560
rect 7630 8520 7660 8560
rect 7560 8460 7660 8520
rect 7560 8420 7590 8460
rect 7630 8420 7660 8460
rect 7560 8360 7660 8420
rect 7560 8320 7590 8360
rect 7630 8320 7660 8360
rect 7560 8290 7660 8320
rect 7780 8660 7880 8690
rect 7780 8620 7810 8660
rect 7850 8620 7880 8660
rect 7780 8560 7880 8620
rect 7780 8520 7810 8560
rect 7850 8520 7880 8560
rect 7780 8460 7880 8520
rect 7780 8420 7810 8460
rect 7850 8420 7880 8460
rect 7780 8360 7880 8420
rect 7780 8320 7810 8360
rect 7850 8320 7880 8360
rect 7780 8290 7880 8320
rect 8000 8660 8100 8690
rect 8000 8620 8030 8660
rect 8070 8620 8100 8660
rect 8000 8560 8100 8620
rect 8000 8520 8030 8560
rect 8070 8520 8100 8560
rect 8000 8460 8100 8520
rect 8000 8420 8030 8460
rect 8070 8420 8100 8460
rect 8000 8360 8100 8420
rect 8000 8320 8030 8360
rect 8070 8320 8100 8360
rect 8000 8290 8100 8320
rect 8220 8660 8320 8690
rect 8420 8660 8520 8690
rect 8220 8620 8250 8660
rect 8290 8620 8320 8660
rect 8420 8620 8450 8660
rect 8490 8620 8520 8660
rect 8220 8560 8320 8620
rect 8420 8560 8520 8620
rect 8220 8520 8250 8560
rect 8290 8520 8320 8560
rect 8420 8520 8450 8560
rect 8490 8520 8520 8560
rect 8220 8460 8320 8520
rect 8420 8460 8520 8520
rect 8220 8420 8250 8460
rect 8290 8420 8320 8460
rect 8420 8420 8450 8460
rect 8490 8420 8520 8460
rect 8220 8360 8320 8420
rect 8420 8360 8520 8420
rect 8220 8320 8250 8360
rect 8290 8320 8320 8360
rect 8420 8320 8450 8360
rect 8490 8320 8520 8360
rect 8220 8290 8320 8320
rect 8420 8290 8520 8320
rect 8640 8660 8740 8690
rect 8640 8620 8670 8660
rect 8710 8620 8740 8660
rect 8640 8560 8740 8620
rect 8640 8520 8670 8560
rect 8710 8520 8740 8560
rect 8640 8460 8740 8520
rect 8640 8420 8670 8460
rect 8710 8420 8740 8460
rect 8640 8360 8740 8420
rect 8640 8320 8670 8360
rect 8710 8320 8740 8360
rect 8640 8290 8740 8320
rect 8860 8660 8960 8690
rect 8860 8620 8890 8660
rect 8930 8620 8960 8660
rect 8860 8560 8960 8620
rect 8860 8520 8890 8560
rect 8930 8520 8960 8560
rect 8860 8460 8960 8520
rect 8860 8420 8890 8460
rect 8930 8420 8960 8460
rect 8860 8360 8960 8420
rect 8860 8320 8890 8360
rect 8930 8320 8960 8360
rect 8860 8290 8960 8320
rect 9080 8660 9180 8690
rect 9080 8620 9110 8660
rect 9150 8620 9180 8660
rect 9080 8560 9180 8620
rect 9080 8520 9110 8560
rect 9150 8520 9180 8560
rect 9080 8460 9180 8520
rect 9080 8420 9110 8460
rect 9150 8420 9180 8460
rect 9080 8360 9180 8420
rect 9080 8320 9110 8360
rect 9150 8320 9180 8360
rect 9080 8290 9180 8320
rect 9300 8660 9400 8690
rect 9500 8660 9600 8690
rect 9300 8620 9330 8660
rect 9370 8620 9400 8660
rect 9500 8620 9530 8660
rect 9570 8620 9600 8660
rect 9300 8560 9400 8620
rect 9500 8560 9600 8620
rect 9300 8520 9330 8560
rect 9370 8520 9400 8560
rect 9500 8520 9530 8560
rect 9570 8520 9600 8560
rect 9300 8460 9400 8520
rect 9500 8460 9600 8520
rect 9300 8420 9330 8460
rect 9370 8420 9400 8460
rect 9500 8420 9530 8460
rect 9570 8420 9600 8460
rect 9300 8360 9400 8420
rect 9500 8360 9600 8420
rect 9300 8320 9330 8360
rect 9370 8320 9400 8360
rect 9500 8320 9530 8360
rect 9570 8320 9600 8360
rect 9300 8290 9400 8320
rect 9500 8290 9600 8320
rect 9720 8660 9820 8690
rect 9720 8620 9750 8660
rect 9790 8620 9820 8660
rect 9720 8560 9820 8620
rect 9720 8520 9750 8560
rect 9790 8520 9820 8560
rect 9720 8460 9820 8520
rect 9720 8420 9750 8460
rect 9790 8420 9820 8460
rect 9720 8360 9820 8420
rect 9720 8320 9750 8360
rect 9790 8320 9820 8360
rect 9720 8290 9820 8320
rect 9940 8660 10040 8690
rect 9940 8620 9970 8660
rect 10010 8620 10040 8660
rect 9940 8560 10040 8620
rect 9940 8520 9970 8560
rect 10010 8520 10040 8560
rect 9940 8460 10040 8520
rect 9940 8420 9970 8460
rect 10010 8420 10040 8460
rect 9940 8360 10040 8420
rect 9940 8320 9970 8360
rect 10010 8320 10040 8360
rect 9940 8290 10040 8320
rect 10160 8660 10260 8690
rect 10160 8620 10190 8660
rect 10230 8620 10260 8660
rect 10160 8560 10260 8620
rect 10160 8520 10190 8560
rect 10230 8520 10260 8560
rect 10160 8460 10260 8520
rect 10160 8420 10190 8460
rect 10230 8420 10260 8460
rect 10160 8360 10260 8420
rect 10160 8320 10190 8360
rect 10230 8320 10260 8360
rect 10160 8290 10260 8320
rect 10380 8660 10480 8690
rect 10380 8620 10410 8660
rect 10450 8620 10480 8660
rect 10380 8560 10480 8620
rect 10380 8520 10410 8560
rect 10450 8520 10480 8560
rect 10380 8460 10480 8520
rect 10380 8420 10410 8460
rect 10450 8420 10480 8460
rect 10380 8360 10480 8420
rect 10380 8320 10410 8360
rect 10450 8320 10480 8360
rect 10380 8290 10480 8320
rect 5980 8240 6080 8270
rect 7400 6030 7500 6060
rect 7400 5980 7430 6030
rect 7470 5980 7500 6030
rect 7400 5890 7500 5980
rect 7400 5840 7430 5890
rect 7470 5840 7500 5890
rect 7400 5810 7500 5840
rect 7600 6030 7700 6060
rect 7600 5980 7630 6030
rect 7670 5980 7700 6030
rect 7600 5890 7700 5980
rect 7600 5840 7630 5890
rect 7670 5840 7700 5890
rect 7600 5810 7700 5840
rect 7800 6030 7900 6060
rect 7800 5980 7830 6030
rect 7870 5980 7900 6030
rect 7800 5890 7900 5980
rect 7800 5840 7830 5890
rect 7870 5840 7900 5890
rect 7800 5810 7900 5840
rect 8000 6030 8100 6060
rect 8000 5980 8030 6030
rect 8070 5980 8100 6030
rect 8000 5890 8100 5980
rect 8000 5840 8030 5890
rect 8070 5840 8100 5890
rect 8000 5810 8100 5840
rect 8200 6030 8300 6060
rect 8200 5980 8230 6030
rect 8270 5980 8300 6030
rect 8200 5890 8300 5980
rect 8200 5840 8230 5890
rect 8270 5840 8300 5890
rect 8200 5810 8300 5840
rect 8400 6030 8500 6060
rect 8400 5980 8430 6030
rect 8470 5980 8500 6030
rect 8400 5890 8500 5980
rect 8400 5840 8430 5890
rect 8470 5840 8500 5890
rect 8400 5810 8500 5840
rect 8600 6030 8700 6060
rect 8600 5980 8630 6030
rect 8670 5980 8700 6030
rect 8600 5890 8700 5980
rect 8600 5840 8630 5890
rect 8670 5840 8700 5890
rect 8600 5810 8700 5840
rect 8800 6030 8900 6060
rect 8800 5980 8830 6030
rect 8870 5980 8900 6030
rect 8800 5890 8900 5980
rect 8800 5840 8830 5890
rect 8870 5840 8900 5890
rect 8800 5810 8900 5840
rect 9000 6030 9100 6060
rect 9000 5980 9030 6030
rect 9070 5980 9100 6030
rect 9000 5890 9100 5980
rect 9000 5840 9030 5890
rect 9070 5840 9100 5890
rect 9000 5810 9100 5840
rect 9200 6030 9300 6060
rect 9200 5980 9230 6030
rect 9270 5980 9300 6030
rect 9200 5890 9300 5980
rect 9200 5840 9230 5890
rect 9270 5840 9300 5890
rect 9200 5810 9300 5840
rect 9400 6030 9500 6060
rect 9400 5980 9430 6030
rect 9470 5980 9500 6030
rect 9400 5890 9500 5980
rect 9400 5840 9430 5890
rect 9470 5840 9500 5890
rect 9400 5810 9500 5840
rect 7450 5340 7550 5370
rect 7450 5300 7480 5340
rect 7520 5300 7550 5340
rect 7450 5270 7550 5300
rect 7580 5340 7680 5370
rect 7580 5300 7610 5340
rect 7650 5300 7680 5340
rect 7580 5270 7680 5300
rect 7710 5340 7810 5370
rect 7710 5300 7740 5340
rect 7780 5300 7810 5340
rect 7710 5270 7810 5300
rect 7840 5340 7940 5370
rect 7840 5300 7870 5340
rect 7910 5300 7940 5340
rect 7840 5270 7940 5300
rect 7970 5340 8070 5370
rect 7970 5300 8000 5340
rect 8040 5300 8070 5340
rect 7970 5270 8070 5300
rect 8100 5340 8200 5370
rect 8100 5300 8130 5340
rect 8170 5300 8200 5340
rect 8100 5270 8200 5300
rect 8230 5340 8330 5370
rect 8230 5300 8260 5340
rect 8300 5300 8330 5340
rect 8230 5270 8330 5300
rect 8590 5340 8690 5370
rect 8590 5300 8620 5340
rect 8660 5300 8690 5340
rect 8590 5270 8690 5300
rect 8720 5340 8820 5370
rect 8720 5300 8750 5340
rect 8790 5300 8820 5340
rect 8720 5270 8820 5300
rect 8850 5340 8950 5370
rect 8850 5300 8880 5340
rect 8920 5300 8950 5340
rect 8850 5270 8950 5300
rect 8980 5340 9080 5370
rect 8980 5300 9010 5340
rect 9050 5300 9080 5340
rect 8980 5270 9080 5300
rect 9110 5340 9210 5370
rect 9110 5300 9140 5340
rect 9180 5300 9210 5340
rect 9110 5270 9210 5300
rect 9240 5340 9340 5370
rect 9240 5300 9270 5340
rect 9310 5300 9340 5340
rect 9240 5270 9340 5300
rect 9370 5340 9470 5370
rect 9370 5300 9400 5340
rect 9440 5300 9470 5340
rect 9370 5270 9470 5300
rect 9730 5340 9830 5370
rect 9730 5300 9760 5340
rect 9800 5300 9830 5340
rect 9730 5270 9830 5300
rect 9860 5340 9960 5370
rect 9860 5300 9890 5340
rect 9930 5300 9960 5340
rect 9860 5270 9960 5300
rect 9990 5340 10090 5370
rect 9990 5300 10020 5340
rect 10060 5300 10090 5340
rect 9990 5270 10090 5300
rect 10120 5340 10220 5370
rect 10120 5300 10150 5340
rect 10190 5300 10220 5340
rect 10120 5270 10220 5300
rect 10250 5340 10350 5370
rect 10250 5300 10280 5340
rect 10320 5300 10350 5340
rect 10250 5270 10350 5300
rect 10380 5340 10480 5370
rect 10380 5300 10410 5340
rect 10450 5300 10480 5340
rect 10380 5270 10480 5300
rect 10510 5340 10610 5370
rect 10510 5300 10540 5340
rect 10580 5300 10610 5340
rect 10510 5270 10610 5300
rect -630 3740 -550 3770
rect -630 3700 -610 3740
rect -570 3700 -550 3740
rect -630 3670 -550 3700
rect -510 3740 -430 3770
rect -510 3700 -490 3740
rect -450 3700 -430 3740
rect -510 3670 -430 3700
rect -390 3740 -310 3770
rect -390 3700 -370 3740
rect -330 3700 -310 3740
rect -390 3670 -310 3700
rect -270 3740 -190 3770
rect -270 3700 -250 3740
rect -210 3700 -190 3740
rect -270 3670 -190 3700
rect -150 3740 -70 3770
rect -150 3700 -130 3740
rect -90 3700 -70 3740
rect -150 3670 -70 3700
rect -30 3740 50 3770
rect -30 3700 -10 3740
rect 30 3700 50 3740
rect -30 3670 50 3700
rect 90 3740 170 3770
rect 90 3700 110 3740
rect 150 3700 170 3740
rect 90 3670 170 3700
rect 210 3740 290 3770
rect 210 3700 230 3740
rect 270 3700 290 3740
rect 210 3670 290 3700
rect 330 3740 410 3770
rect 330 3700 350 3740
rect 390 3700 410 3740
rect 330 3670 410 3700
rect 450 3740 530 3770
rect 450 3700 470 3740
rect 510 3700 530 3740
rect 450 3670 530 3700
rect 570 3740 650 3770
rect 570 3700 590 3740
rect 630 3700 650 3740
rect 570 3670 650 3700
rect 1930 3740 2010 3770
rect 1930 3700 1950 3740
rect 1990 3700 2010 3740
rect 1930 3670 2010 3700
rect 2050 3740 2130 3770
rect 2050 3700 2070 3740
rect 2110 3700 2130 3740
rect 2050 3670 2130 3700
rect 2170 3740 2250 3770
rect 2170 3700 2190 3740
rect 2230 3700 2250 3740
rect 2170 3670 2250 3700
rect 2290 3740 2370 3770
rect 2290 3700 2310 3740
rect 2350 3700 2370 3740
rect 2290 3670 2370 3700
rect 2410 3740 2490 3770
rect 2410 3700 2430 3740
rect 2470 3700 2490 3740
rect 2410 3670 2490 3700
rect 2530 3740 2610 3770
rect 2530 3700 2550 3740
rect 2590 3700 2610 3740
rect 2530 3670 2610 3700
rect 2650 3740 2730 3770
rect 2650 3700 2670 3740
rect 2710 3700 2730 3740
rect 2650 3670 2730 3700
rect 2770 3740 2850 3770
rect 2770 3700 2790 3740
rect 2830 3700 2850 3740
rect 2770 3670 2850 3700
rect 2890 3740 2970 3770
rect 2890 3700 2910 3740
rect 2950 3700 2970 3740
rect 2890 3670 2970 3700
rect 3010 3740 3090 3770
rect 3010 3700 3030 3740
rect 3070 3700 3090 3740
rect 3010 3670 3090 3700
rect 3130 3740 3210 3770
rect 3130 3700 3150 3740
rect 3190 3700 3210 3740
rect 3130 3670 3210 3700
rect -1250 3130 -1170 3160
rect -1250 3090 -1230 3130
rect -1190 3090 -1170 3130
rect -1250 3030 -1170 3090
rect -1250 2990 -1230 3030
rect -1190 2990 -1170 3030
rect -1250 2930 -1170 2990
rect -1250 2890 -1230 2930
rect -1190 2890 -1170 2930
rect -1250 2830 -1170 2890
rect -1250 2790 -1230 2830
rect -1190 2790 -1170 2830
rect -1250 2730 -1170 2790
rect -1250 2690 -1230 2730
rect -1190 2690 -1170 2730
rect -1250 2660 -1170 2690
rect -170 3130 -90 3160
rect -10 3130 70 3160
rect -170 3090 -150 3130
rect -110 3090 -90 3130
rect -10 3090 10 3130
rect 50 3090 70 3130
rect -170 3030 -90 3090
rect -10 3030 70 3090
rect -170 2990 -150 3030
rect -110 2990 -90 3030
rect -10 2990 10 3030
rect 50 2990 70 3030
rect -170 2930 -90 2990
rect -10 2930 70 2990
rect -170 2890 -150 2930
rect -110 2890 -90 2930
rect -10 2890 10 2930
rect 50 2890 70 2930
rect -170 2830 -90 2890
rect -10 2830 70 2890
rect -170 2790 -150 2830
rect -110 2790 -90 2830
rect -10 2790 10 2830
rect 50 2790 70 2830
rect -170 2730 -90 2790
rect -10 2730 70 2790
rect -170 2690 -150 2730
rect -110 2690 -90 2730
rect -10 2690 10 2730
rect 50 2690 70 2730
rect -170 2660 -90 2690
rect -10 2660 70 2690
rect 1070 3130 1150 3160
rect 1070 3090 1090 3130
rect 1130 3090 1150 3130
rect 1070 3030 1150 3090
rect 1070 2990 1090 3030
rect 1130 2990 1150 3030
rect 1070 2930 1150 2990
rect 1070 2890 1090 2930
rect 1130 2890 1150 2930
rect 1070 2830 1150 2890
rect 1070 2790 1090 2830
rect 1130 2790 1150 2830
rect 1070 2730 1150 2790
rect 1070 2690 1090 2730
rect 1130 2690 1150 2730
rect 1070 2660 1150 2690
rect 1430 3130 1510 3160
rect 1430 3090 1450 3130
rect 1490 3090 1510 3130
rect 1430 3030 1510 3090
rect 1430 2990 1450 3030
rect 1490 2990 1510 3030
rect 1430 2930 1510 2990
rect 1430 2890 1450 2930
rect 1490 2890 1510 2930
rect 1430 2830 1510 2890
rect 1430 2790 1450 2830
rect 1490 2790 1510 2830
rect 1430 2730 1510 2790
rect 1430 2690 1450 2730
rect 1490 2690 1510 2730
rect 1430 2660 1510 2690
rect 2510 3130 2590 3160
rect 2670 3130 2750 3160
rect 2510 3090 2530 3130
rect 2570 3090 2590 3130
rect 2670 3090 2690 3130
rect 2730 3090 2750 3130
rect 2510 3030 2590 3090
rect 2670 3030 2750 3090
rect 2510 2990 2530 3030
rect 2570 2990 2590 3030
rect 2670 2990 2690 3030
rect 2730 2990 2750 3030
rect 2510 2930 2590 2990
rect 2670 2930 2750 2990
rect 2510 2890 2530 2930
rect 2570 2890 2590 2930
rect 2670 2890 2690 2930
rect 2730 2890 2750 2930
rect 2510 2830 2590 2890
rect 2670 2830 2750 2890
rect 2510 2790 2530 2830
rect 2570 2790 2590 2830
rect 2670 2790 2690 2830
rect 2730 2790 2750 2830
rect 2510 2730 2590 2790
rect 2670 2730 2750 2790
rect 2510 2690 2530 2730
rect 2570 2690 2590 2730
rect 2670 2690 2690 2730
rect 2730 2690 2750 2730
rect 2510 2670 2590 2690
rect 2670 2670 2750 2690
rect 2510 2660 2750 2670
rect 3750 3130 3830 3160
rect 3750 3090 3770 3130
rect 3810 3090 3830 3130
rect 3750 3030 3830 3090
rect 3750 2990 3770 3030
rect 3810 2990 3830 3030
rect 3750 2930 3830 2990
rect 3750 2890 3770 2930
rect 3810 2890 3830 2930
rect 3750 2830 3830 2890
rect 3750 2790 3770 2830
rect 3810 2790 3830 2830
rect 3750 2730 3830 2790
rect 3750 2690 3770 2730
rect 3810 2690 3830 2730
rect 3750 2660 3830 2690
rect -830 2220 -750 2250
rect -830 2180 -810 2220
rect -770 2180 -750 2220
rect -830 2120 -750 2180
rect -830 2080 -810 2120
rect -770 2080 -750 2120
rect -830 2050 -750 2080
rect 1250 2220 1330 2250
rect 1250 2180 1270 2220
rect 1310 2180 1330 2220
rect 1250 2120 1330 2180
rect 1250 2080 1270 2120
rect 1310 2080 1330 2120
rect 1250 2050 1330 2080
rect 3330 2220 3410 2250
rect 3330 2180 3350 2220
rect 3390 2180 3410 2220
rect 3330 2120 3410 2180
rect 3330 2080 3350 2120
rect 3390 2080 3410 2120
rect 3330 2050 3410 2080
<< pdiff >>
rect 600 12870 680 12900
rect 600 12830 620 12870
rect 660 12830 680 12870
rect 600 12800 680 12830
rect 710 12870 790 12900
rect 710 12830 730 12870
rect 770 12830 790 12870
rect 710 12800 790 12830
rect 1020 12870 1100 12900
rect 1020 12830 1040 12870
rect 1080 12830 1100 12870
rect 1020 12800 1100 12830
rect 1130 12870 1210 12900
rect 1130 12830 1150 12870
rect 1190 12830 1210 12870
rect 1130 12800 1210 12830
rect 1240 12870 1320 12900
rect 1240 12830 1260 12870
rect 1300 12830 1320 12870
rect 1240 12800 1320 12830
rect 1690 12870 1770 12900
rect 1690 12830 1710 12870
rect 1750 12830 1770 12870
rect 1690 12800 1770 12830
rect 1800 12870 1880 12900
rect 1800 12830 1820 12870
rect 1860 12830 1880 12870
rect 1800 12800 1880 12830
rect 1910 12870 1990 12900
rect 1910 12830 1930 12870
rect 1970 12830 1990 12870
rect 1910 12800 1990 12830
rect 2130 12870 2210 12900
rect 2130 12830 2150 12870
rect 2190 12830 2210 12870
rect 2130 12800 2210 12830
rect 2240 12870 2320 12900
rect 2240 12830 2260 12870
rect 2300 12830 2320 12870
rect 2240 12800 2320 12830
rect 2350 12870 2430 12900
rect 2350 12830 2370 12870
rect 2410 12830 2430 12870
rect 2350 12800 2430 12830
rect 2460 12870 2540 12900
rect 2460 12830 2480 12870
rect 2520 12830 2540 12870
rect 2460 12800 2540 12830
rect 2970 12870 3050 12900
rect 2970 12830 2990 12870
rect 3030 12830 3050 12870
rect 2970 12800 3050 12830
rect 3080 12870 3160 12900
rect 3080 12830 3100 12870
rect 3140 12830 3160 12870
rect 3080 12800 3160 12830
rect 3390 12870 3470 12900
rect 3390 12830 3410 12870
rect 3450 12830 3470 12870
rect 3390 12800 3470 12830
rect 3500 12870 3580 12900
rect 3500 12830 3520 12870
rect 3560 12830 3580 12870
rect 3500 12800 3580 12830
rect 3610 12870 3690 12900
rect 3610 12830 3630 12870
rect 3670 12830 3690 12870
rect 3610 12800 3690 12830
rect 3840 12870 3920 12900
rect 3840 12830 3860 12870
rect 3900 12830 3920 12870
rect 3840 12800 3920 12830
rect 3950 12870 4030 12900
rect 3950 12830 3970 12870
rect 4010 12830 4030 12870
rect 3950 12800 4030 12830
rect 4060 12870 4140 12900
rect 4060 12830 4080 12870
rect 4120 12830 4140 12870
rect 4060 12800 4140 12830
rect 4200 12870 4280 12900
rect 4200 12830 4220 12870
rect 4260 12830 4280 12870
rect 4200 12800 4280 12830
rect 4310 12870 4390 12900
rect 4310 12830 4330 12870
rect 4370 12830 4390 12870
rect 4310 12800 4390 12830
rect 4420 12870 4500 12900
rect 4420 12830 4440 12870
rect 4480 12830 4500 12870
rect 4420 12800 4500 12830
rect 4780 12870 4860 12900
rect 4780 12830 4800 12870
rect 4840 12830 4860 12870
rect 4780 12800 4860 12830
rect 4890 12870 4970 12900
rect 4890 12830 4910 12870
rect 4950 12830 4970 12870
rect 4890 12800 4970 12830
rect 5000 12870 5080 12900
rect 5000 12830 5020 12870
rect 5060 12830 5080 12870
rect 5000 12800 5080 12830
rect 5220 12870 5300 12900
rect 5220 12830 5240 12870
rect 5280 12830 5300 12870
rect 5220 12800 5300 12830
rect 5330 12870 5410 12900
rect 5330 12830 5350 12870
rect 5390 12830 5410 12870
rect 5330 12800 5410 12830
rect 5440 12870 5520 12900
rect 5440 12830 5460 12870
rect 5500 12830 5520 12870
rect 5440 12800 5520 12830
rect 5840 12870 5920 12900
rect 5840 12830 5860 12870
rect 5900 12830 5920 12870
rect 5840 12800 5920 12830
rect 5950 12870 6030 12900
rect 5950 12830 5970 12870
rect 6010 12830 6030 12870
rect 5950 12800 6030 12830
rect 6180 12870 6260 12900
rect 6180 12830 6200 12870
rect 6240 12830 6260 12870
rect 6180 12800 6260 12830
rect 6290 12870 6370 12900
rect 6290 12830 6310 12870
rect 6350 12830 6370 12870
rect 6290 12800 6370 12830
rect 6400 12870 6480 12900
rect 6400 12830 6420 12870
rect 6460 12830 6480 12870
rect 6400 12800 6480 12830
rect 6540 12870 6620 12900
rect 6540 12830 6560 12870
rect 6600 12830 6620 12870
rect 6540 12800 6620 12830
rect 6650 12870 6730 12900
rect 6650 12830 6670 12870
rect 6710 12830 6730 12870
rect 6650 12800 6730 12830
rect 6760 12870 6840 12900
rect 6760 12830 6780 12870
rect 6820 12830 6840 12870
rect 6760 12800 6840 12830
rect 7140 12870 7220 12900
rect 7140 12830 7160 12870
rect 7200 12830 7220 12870
rect 7140 12800 7220 12830
rect 7250 12870 7330 12900
rect 7250 12830 7270 12870
rect 7310 12830 7330 12870
rect 7250 12800 7330 12830
rect 7480 12870 7560 12900
rect 7480 12830 7500 12870
rect 7540 12830 7560 12870
rect 7480 12800 7560 12830
rect 7590 12870 7670 12900
rect 7590 12830 7610 12870
rect 7650 12830 7670 12870
rect 7590 12800 7670 12830
rect 7700 12870 7780 12900
rect 7700 12830 7720 12870
rect 7760 12830 7780 12870
rect 7700 12800 7780 12830
rect 7840 12870 7920 12900
rect 7840 12830 7860 12870
rect 7900 12830 7920 12870
rect 7840 12800 7920 12830
rect 7950 12870 8030 12900
rect 7950 12830 7970 12870
rect 8010 12830 8030 12870
rect 7950 12800 8030 12830
rect 8060 12870 8140 12900
rect 8060 12830 8080 12870
rect 8120 12830 8140 12870
rect 8060 12800 8140 12830
rect 8440 12870 8520 12900
rect 8440 12830 8460 12870
rect 8500 12830 8520 12870
rect 8440 12800 8520 12830
rect 8550 12870 8630 12900
rect 8550 12830 8570 12870
rect 8610 12830 8630 12870
rect 8550 12800 8630 12830
rect 8780 12870 8860 12900
rect 8780 12830 8800 12870
rect 8840 12830 8860 12870
rect 8780 12800 8860 12830
rect 8890 12870 8970 12900
rect 8890 12830 8910 12870
rect 8950 12830 8970 12870
rect 8890 12800 8970 12830
rect 9000 12870 9080 12900
rect 9000 12830 9020 12870
rect 9060 12830 9080 12870
rect 9000 12800 9080 12830
rect 9140 12870 9220 12900
rect 9140 12830 9160 12870
rect 9200 12830 9220 12870
rect 9140 12800 9220 12830
rect 9250 12870 9330 12900
rect 9250 12830 9270 12870
rect 9310 12830 9330 12870
rect 9250 12800 9330 12830
rect 9360 12870 9440 12900
rect 9360 12830 9380 12870
rect 9420 12830 9440 12870
rect 9360 12800 9440 12830
rect 9740 12870 9820 12900
rect 9740 12830 9760 12870
rect 9800 12830 9820 12870
rect 9740 12800 9820 12830
rect 9850 12870 9930 12900
rect 9850 12830 9870 12870
rect 9910 12830 9930 12870
rect 9850 12800 9930 12830
rect 10080 12870 10160 12900
rect 10080 12830 10100 12870
rect 10140 12830 10160 12870
rect 10080 12800 10160 12830
rect 10190 12870 10270 12900
rect 10190 12830 10210 12870
rect 10250 12830 10270 12870
rect 10190 12800 10270 12830
rect 10300 12870 10380 12900
rect 10300 12830 10320 12870
rect 10360 12830 10380 12870
rect 10300 12800 10380 12830
rect 10440 12870 10520 12900
rect 10440 12830 10460 12870
rect 10500 12830 10520 12870
rect 10440 12800 10520 12830
rect 10550 12870 10630 12900
rect 10550 12830 10570 12870
rect 10610 12830 10630 12870
rect 10550 12800 10630 12830
rect 10660 12870 10740 12900
rect 10660 12830 10680 12870
rect 10720 12830 10740 12870
rect 10660 12800 10740 12830
rect 11208 12740 11288 12770
rect 11208 12700 11228 12740
rect 11268 12700 11288 12740
rect 11208 12640 11288 12700
rect 11208 12600 11228 12640
rect 11268 12600 11288 12640
rect 11208 12540 11288 12600
rect 11208 12500 11228 12540
rect 11268 12500 11288 12540
rect 11208 12440 11288 12500
rect 11208 12400 11228 12440
rect 11268 12400 11288 12440
rect 11208 12370 11288 12400
rect 11320 12740 11400 12770
rect 11320 12700 11340 12740
rect 11380 12700 11400 12740
rect 11320 12640 11400 12700
rect 11320 12600 11340 12640
rect 11380 12600 11400 12640
rect 11320 12540 11400 12600
rect 11320 12500 11340 12540
rect 11380 12500 11400 12540
rect 11320 12440 11400 12500
rect 11320 12400 11340 12440
rect 11380 12400 11400 12440
rect 11320 12370 11400 12400
rect 11728 12740 11808 12770
rect 11728 12700 11748 12740
rect 11788 12700 11808 12740
rect 11728 12640 11808 12700
rect 11728 12600 11748 12640
rect 11788 12600 11808 12640
rect 11728 12540 11808 12600
rect 11728 12500 11748 12540
rect 11788 12500 11808 12540
rect 11728 12440 11808 12500
rect 11728 12400 11748 12440
rect 11788 12400 11808 12440
rect 11728 12370 11808 12400
rect 11840 12740 11920 12770
rect 11840 12700 11860 12740
rect 11900 12700 11920 12740
rect 11840 12640 11920 12700
rect 11840 12600 11860 12640
rect 11900 12600 11920 12640
rect 11840 12540 11920 12600
rect 11840 12500 11860 12540
rect 11900 12500 11920 12540
rect 11840 12440 11920 12500
rect 11840 12400 11860 12440
rect 11900 12400 11920 12440
rect 11840 12370 11920 12400
rect 12248 12740 12328 12770
rect 12248 12700 12268 12740
rect 12308 12700 12328 12740
rect 12248 12640 12328 12700
rect 12248 12600 12268 12640
rect 12308 12600 12328 12640
rect 12248 12540 12328 12600
rect 12248 12500 12268 12540
rect 12308 12500 12328 12540
rect 12248 12440 12328 12500
rect 12248 12400 12268 12440
rect 12308 12400 12328 12440
rect 12248 12370 12328 12400
rect 12360 12740 12440 12770
rect 12360 12700 12380 12740
rect 12420 12700 12440 12740
rect 12360 12640 12440 12700
rect 12360 12600 12380 12640
rect 12420 12600 12440 12640
rect 12360 12540 12440 12600
rect 12360 12500 12380 12540
rect 12420 12500 12440 12540
rect 12360 12440 12440 12500
rect 12360 12400 12380 12440
rect 12420 12400 12440 12440
rect 12360 12370 12440 12400
rect 11210 12160 11290 12190
rect 11210 12120 11230 12160
rect 11270 12120 11290 12160
rect 11210 12060 11290 12120
rect 11210 12020 11230 12060
rect 11270 12020 11290 12060
rect 11210 11960 11290 12020
rect 11210 11920 11230 11960
rect 11270 11920 11290 11960
rect 11210 11860 11290 11920
rect 11210 11820 11230 11860
rect 11270 11820 11290 11860
rect 11210 11760 11290 11820
rect 11210 11720 11230 11760
rect 11270 11720 11290 11760
rect 11210 11660 11290 11720
rect 11210 11620 11230 11660
rect 11270 11620 11290 11660
rect 11210 11590 11290 11620
rect 11320 12160 11400 12190
rect 11320 12120 11340 12160
rect 11380 12120 11400 12160
rect 11320 12060 11400 12120
rect 11320 12020 11340 12060
rect 11380 12020 11400 12060
rect 11320 11960 11400 12020
rect 11320 11920 11340 11960
rect 11380 11920 11400 11960
rect 11320 11860 11400 11920
rect 11320 11820 11340 11860
rect 11380 11820 11400 11860
rect 11320 11760 11400 11820
rect 11320 11720 11340 11760
rect 11380 11720 11400 11760
rect 11320 11660 11400 11720
rect 11320 11620 11340 11660
rect 11380 11620 11400 11660
rect 11320 11590 11400 11620
rect 11730 12160 11810 12190
rect 11730 12120 11750 12160
rect 11790 12120 11810 12160
rect 11730 12060 11810 12120
rect 11730 12020 11750 12060
rect 11790 12020 11810 12060
rect 11730 11960 11810 12020
rect 11730 11920 11750 11960
rect 11790 11920 11810 11960
rect 11730 11860 11810 11920
rect 11730 11820 11750 11860
rect 11790 11820 11810 11860
rect 11730 11760 11810 11820
rect 11730 11720 11750 11760
rect 11790 11720 11810 11760
rect 11730 11660 11810 11720
rect 11730 11620 11750 11660
rect 11790 11620 11810 11660
rect 11730 11590 11810 11620
rect 11840 12160 11920 12190
rect 11840 12120 11860 12160
rect 11900 12120 11920 12160
rect 11840 12060 11920 12120
rect 11840 12020 11860 12060
rect 11900 12020 11920 12060
rect 11840 11960 11920 12020
rect 11840 11920 11860 11960
rect 11900 11920 11920 11960
rect 11840 11860 11920 11920
rect 11840 11820 11860 11860
rect 11900 11820 11920 11860
rect 11840 11760 11920 11820
rect 11840 11720 11860 11760
rect 11900 11720 11920 11760
rect 11840 11660 11920 11720
rect 11840 11620 11860 11660
rect 11900 11620 11920 11660
rect 11840 11590 11920 11620
rect 12250 12160 12330 12190
rect 12250 12120 12270 12160
rect 12310 12120 12330 12160
rect 12250 12060 12330 12120
rect 12250 12020 12270 12060
rect 12310 12020 12330 12060
rect 12250 11960 12330 12020
rect 12250 11920 12270 11960
rect 12310 11920 12330 11960
rect 12250 11860 12330 11920
rect 12250 11820 12270 11860
rect 12310 11820 12330 11860
rect 12250 11760 12330 11820
rect 12250 11720 12270 11760
rect 12310 11720 12330 11760
rect 12250 11660 12330 11720
rect 12250 11620 12270 11660
rect 12310 11620 12330 11660
rect 12250 11590 12330 11620
rect 12360 12160 12440 12190
rect 12360 12120 12380 12160
rect 12420 12120 12440 12160
rect 12360 12060 12440 12120
rect 12360 12020 12380 12060
rect 12420 12020 12440 12060
rect 12360 11960 12440 12020
rect 12360 11920 12380 11960
rect 12420 11920 12440 11960
rect 12360 11860 12440 11920
rect 12360 11820 12380 11860
rect 12420 11820 12440 11860
rect 12360 11760 12440 11820
rect 12360 11720 12380 11760
rect 12420 11720 12440 11760
rect 12360 11660 12440 11720
rect 12360 11620 12380 11660
rect 12420 11620 12440 11660
rect 12360 11590 12440 11620
rect 11210 11270 11290 11300
rect 11210 11230 11230 11270
rect 11270 11230 11290 11270
rect 11210 11170 11290 11230
rect 11210 11130 11230 11170
rect 11270 11130 11290 11170
rect 11210 11070 11290 11130
rect 11210 11030 11230 11070
rect 11270 11030 11290 11070
rect 11210 10970 11290 11030
rect 11210 10930 11230 10970
rect 11270 10930 11290 10970
rect 11210 10900 11290 10930
rect 11590 11270 11670 11300
rect 11590 11230 11610 11270
rect 11650 11230 11670 11270
rect 11590 11170 11670 11230
rect 11590 11130 11610 11170
rect 11650 11130 11670 11170
rect 11590 11070 11670 11130
rect 11590 11030 11610 11070
rect 11650 11030 11670 11070
rect 11590 10970 11670 11030
rect 11590 10930 11610 10970
rect 11650 10930 11670 10970
rect 11590 10900 11670 10930
rect 11730 11270 11810 11300
rect 11730 11230 11750 11270
rect 11790 11230 11810 11270
rect 11730 11170 11810 11230
rect 11730 11130 11750 11170
rect 11790 11130 11810 11170
rect 11730 11070 11810 11130
rect 11730 11030 11750 11070
rect 11790 11030 11810 11070
rect 11730 10970 11810 11030
rect 11730 10930 11750 10970
rect 11790 10930 11810 10970
rect 11730 10900 11810 10930
rect 12110 11270 12190 11300
rect 12110 11230 12130 11270
rect 12170 11230 12190 11270
rect 12110 11170 12190 11230
rect 12110 11130 12130 11170
rect 12170 11130 12190 11170
rect 12110 11070 12190 11130
rect 12110 11030 12130 11070
rect 12170 11030 12190 11070
rect 12110 10970 12190 11030
rect 12110 10930 12130 10970
rect 12170 10930 12190 10970
rect 12110 10900 12190 10930
rect 12250 11270 12330 11300
rect 12250 11230 12270 11270
rect 12310 11230 12330 11270
rect 12250 11170 12330 11230
rect 12250 11130 12270 11170
rect 12310 11130 12330 11170
rect 12250 11070 12330 11130
rect 12250 11030 12270 11070
rect 12310 11030 12330 11070
rect 12250 10970 12330 11030
rect 12250 10930 12270 10970
rect 12310 10930 12330 10970
rect 12250 10900 12330 10930
rect 12630 11270 12710 11300
rect 12630 11230 12650 11270
rect 12690 11230 12710 11270
rect 12630 11170 12710 11230
rect 12630 11130 12650 11170
rect 12690 11130 12710 11170
rect 12630 11070 12710 11130
rect 12630 11030 12650 11070
rect 12690 11030 12710 11070
rect 12630 10970 12710 11030
rect 12630 10930 12650 10970
rect 12690 10930 12710 10970
rect 12630 10900 12710 10930
rect 12770 11270 12850 11300
rect 12770 11230 12790 11270
rect 12830 11230 12850 11270
rect 12770 11170 12850 11230
rect 12770 11130 12790 11170
rect 12830 11130 12850 11170
rect 12770 11070 12850 11130
rect 12770 11030 12790 11070
rect 12830 11030 12850 11070
rect 12770 10970 12850 11030
rect 12770 10930 12790 10970
rect 12830 10930 12850 10970
rect 12770 10900 12850 10930
rect 13150 11270 13230 11300
rect 13150 11230 13170 11270
rect 13210 11230 13230 11270
rect 13150 11170 13230 11230
rect 13150 11130 13170 11170
rect 13210 11130 13230 11170
rect 13150 11070 13230 11130
rect 13150 11030 13170 11070
rect 13210 11030 13230 11070
rect 13150 10970 13230 11030
rect 13150 10930 13170 10970
rect 13210 10930 13230 10970
rect 13150 10900 13230 10930
rect 1260 9790 1340 9820
rect 1260 9750 1280 9790
rect 1320 9750 1340 9790
rect 1260 9690 1340 9750
rect 1260 9650 1280 9690
rect 1320 9650 1340 9690
rect 1260 9590 1340 9650
rect 1260 9550 1280 9590
rect 1320 9550 1340 9590
rect 1260 9490 1340 9550
rect 1260 9450 1280 9490
rect 1320 9450 1340 9490
rect 1260 9420 1340 9450
rect 1370 9790 1450 9820
rect 1370 9750 1390 9790
rect 1430 9750 1450 9790
rect 1370 9690 1450 9750
rect 1370 9650 1390 9690
rect 1430 9650 1450 9690
rect 1370 9590 1450 9650
rect 1370 9550 1390 9590
rect 1430 9550 1450 9590
rect 1370 9490 1450 9550
rect 1370 9450 1390 9490
rect 1430 9450 1450 9490
rect 1370 9420 1450 9450
rect 1480 9790 1560 9820
rect 1480 9750 1500 9790
rect 1540 9750 1560 9790
rect 1480 9690 1560 9750
rect 1480 9650 1500 9690
rect 1540 9650 1560 9690
rect 1480 9590 1560 9650
rect 1480 9550 1500 9590
rect 1540 9550 1560 9590
rect 1480 9490 1560 9550
rect 1480 9450 1500 9490
rect 1540 9450 1560 9490
rect 1480 9420 1560 9450
rect 1780 9790 1860 9820
rect 1780 9750 1800 9790
rect 1840 9750 1860 9790
rect 1780 9690 1860 9750
rect 1780 9650 1800 9690
rect 1840 9650 1860 9690
rect 1780 9590 1860 9650
rect 1780 9550 1800 9590
rect 1840 9550 1860 9590
rect 1780 9490 1860 9550
rect 1780 9450 1800 9490
rect 1840 9450 1860 9490
rect 1780 9420 1860 9450
rect 1890 9790 1970 9820
rect 1890 9750 1910 9790
rect 1950 9750 1970 9790
rect 1890 9690 1970 9750
rect 1890 9650 1910 9690
rect 1950 9650 1970 9690
rect 1890 9590 1970 9650
rect 1890 9550 1910 9590
rect 1950 9550 1970 9590
rect 1890 9490 1970 9550
rect 1890 9450 1910 9490
rect 1950 9450 1970 9490
rect 1890 9420 1970 9450
rect 2000 9790 2080 9820
rect 2160 9790 2240 9820
rect 2000 9750 2020 9790
rect 2060 9750 2080 9790
rect 2160 9750 2180 9790
rect 2220 9750 2240 9790
rect 2000 9690 2080 9750
rect 2160 9690 2240 9750
rect 2000 9650 2020 9690
rect 2060 9650 2080 9690
rect 2160 9650 2180 9690
rect 2220 9650 2240 9690
rect 2000 9590 2080 9650
rect 2160 9590 2240 9650
rect 2000 9550 2020 9590
rect 2060 9550 2080 9590
rect 2160 9550 2180 9590
rect 2220 9550 2240 9590
rect 2000 9490 2080 9550
rect 2160 9490 2240 9550
rect 2000 9450 2020 9490
rect 2060 9450 2080 9490
rect 2160 9450 2180 9490
rect 2220 9450 2240 9490
rect 2000 9420 2080 9450
rect 2160 9420 2240 9450
rect 2270 9790 2350 9820
rect 2270 9750 2290 9790
rect 2330 9750 2350 9790
rect 2270 9690 2350 9750
rect 2270 9650 2290 9690
rect 2330 9650 2350 9690
rect 2270 9590 2350 9650
rect 2270 9550 2290 9590
rect 2330 9550 2350 9590
rect 2270 9490 2350 9550
rect 2270 9450 2290 9490
rect 2330 9450 2350 9490
rect 2270 9420 2350 9450
rect 2380 9790 2460 9820
rect 2380 9750 2400 9790
rect 2440 9750 2460 9790
rect 2380 9690 2460 9750
rect 2380 9650 2400 9690
rect 2440 9650 2460 9690
rect 2380 9590 2460 9650
rect 2380 9550 2400 9590
rect 2440 9550 2460 9590
rect 2380 9490 2460 9550
rect 2380 9450 2400 9490
rect 2440 9450 2460 9490
rect 2380 9420 2460 9450
rect 2680 9790 2760 9820
rect 2680 9750 2700 9790
rect 2740 9750 2760 9790
rect 2680 9690 2760 9750
rect 2680 9650 2700 9690
rect 2740 9650 2760 9690
rect 2680 9590 2760 9650
rect 2680 9550 2700 9590
rect 2740 9550 2760 9590
rect 2680 9490 2760 9550
rect 2680 9450 2700 9490
rect 2740 9450 2760 9490
rect 2680 9420 2760 9450
rect 2790 9790 2870 9820
rect 2790 9750 2810 9790
rect 2850 9750 2870 9790
rect 2790 9690 2870 9750
rect 2790 9650 2810 9690
rect 2850 9650 2870 9690
rect 2790 9590 2870 9650
rect 2790 9550 2810 9590
rect 2850 9550 2870 9590
rect 2790 9490 2870 9550
rect 2790 9450 2810 9490
rect 2850 9450 2870 9490
rect 2790 9420 2870 9450
rect 2900 9790 2980 9820
rect 2900 9750 2920 9790
rect 2960 9750 2980 9790
rect 2900 9690 2980 9750
rect 2900 9650 2920 9690
rect 2960 9650 2980 9690
rect 2900 9590 2980 9650
rect 2900 9550 2920 9590
rect 2960 9550 2980 9590
rect 2900 9490 2980 9550
rect 2900 9450 2920 9490
rect 2960 9450 2980 9490
rect 2900 9420 2980 9450
rect 3200 9790 3280 9820
rect 3200 9750 3220 9790
rect 3260 9750 3280 9790
rect 3200 9690 3280 9750
rect 3200 9650 3220 9690
rect 3260 9650 3280 9690
rect 3200 9590 3280 9650
rect 3200 9550 3220 9590
rect 3260 9550 3280 9590
rect 3200 9490 3280 9550
rect 3200 9450 3220 9490
rect 3260 9450 3280 9490
rect 3200 9430 3280 9450
rect 3180 9420 3280 9430
rect 3310 9790 3390 9820
rect 3310 9750 3330 9790
rect 3370 9750 3390 9790
rect 3310 9690 3390 9750
rect 3310 9650 3330 9690
rect 3370 9650 3390 9690
rect 3310 9590 3390 9650
rect 3310 9550 3330 9590
rect 3370 9550 3390 9590
rect 3310 9490 3390 9550
rect 3310 9450 3330 9490
rect 3370 9450 3390 9490
rect 3310 9420 3390 9450
rect 3420 9790 3500 9820
rect 3420 9750 3440 9790
rect 3480 9750 3500 9790
rect 3420 9690 3500 9750
rect 3420 9650 3440 9690
rect 3480 9650 3500 9690
rect 3420 9590 3500 9650
rect 3420 9550 3440 9590
rect 3480 9550 3500 9590
rect 3420 9490 3500 9550
rect 3420 9450 3440 9490
rect 3480 9450 3500 9490
rect 3420 9420 3500 9450
rect 3640 9790 3720 9820
rect 3640 9750 3660 9790
rect 3700 9750 3720 9790
rect 3640 9690 3720 9750
rect 3640 9650 3660 9690
rect 3700 9650 3720 9690
rect 3640 9590 3720 9650
rect 3640 9550 3660 9590
rect 3700 9550 3720 9590
rect 3640 9490 3720 9550
rect 3640 9450 3660 9490
rect 3700 9450 3720 9490
rect 3640 9420 3720 9450
rect 3750 9790 3830 9820
rect 3750 9750 3770 9790
rect 3810 9750 3830 9790
rect 3750 9690 3830 9750
rect 3750 9650 3770 9690
rect 3810 9650 3830 9690
rect 3750 9590 3830 9650
rect 3750 9550 3770 9590
rect 3810 9550 3830 9590
rect 3750 9490 3830 9550
rect 3750 9450 3770 9490
rect 3810 9450 3830 9490
rect 3750 9420 3830 9450
rect 3970 9790 4050 9820
rect 3970 9750 3990 9790
rect 4030 9750 4050 9790
rect 3970 9690 4050 9750
rect 3970 9650 3990 9690
rect 4030 9650 4050 9690
rect 3970 9590 4050 9650
rect 3970 9550 3990 9590
rect 4030 9550 4050 9590
rect 3970 9490 4050 9550
rect 3970 9450 3990 9490
rect 4030 9450 4050 9490
rect 3970 9420 4050 9450
rect 4080 9790 4160 9820
rect 4080 9750 4100 9790
rect 4140 9750 4160 9790
rect 4080 9690 4160 9750
rect 4080 9650 4100 9690
rect 4140 9650 4160 9690
rect 4080 9590 4160 9650
rect 4080 9550 4100 9590
rect 4140 9550 4160 9590
rect 4080 9490 4160 9550
rect 4080 9450 4100 9490
rect 4140 9450 4160 9490
rect 4080 9420 4160 9450
rect 4390 9790 4490 9820
rect 4390 9750 4420 9790
rect 4460 9750 4490 9790
rect 4390 9690 4490 9750
rect 4390 9650 4420 9690
rect 4460 9650 4490 9690
rect 4390 9590 4490 9650
rect 4390 9550 4420 9590
rect 4460 9550 4490 9590
rect 4390 9490 4490 9550
rect 4390 9450 4420 9490
rect 4460 9450 4490 9490
rect 4390 9420 4490 9450
rect 4520 9790 4620 9820
rect 4520 9750 4550 9790
rect 4590 9750 4620 9790
rect 4520 9690 4620 9750
rect 4520 9650 4550 9690
rect 4590 9650 4620 9690
rect 4520 9590 4620 9650
rect 4520 9550 4550 9590
rect 4590 9550 4620 9590
rect 4520 9490 4620 9550
rect 4520 9450 4550 9490
rect 4590 9450 4620 9490
rect 4520 9420 4620 9450
rect 4780 9790 4880 9820
rect 4780 9750 4810 9790
rect 4850 9750 4880 9790
rect 4780 9690 4880 9750
rect 4780 9650 4810 9690
rect 4850 9650 4880 9690
rect 4780 9590 4880 9650
rect 4780 9550 4810 9590
rect 4850 9550 4880 9590
rect 4780 9490 4880 9550
rect 4780 9450 4810 9490
rect 4850 9450 4880 9490
rect 4780 9420 4880 9450
rect 4910 9790 5010 9820
rect 4910 9750 4940 9790
rect 4980 9750 5010 9790
rect 4910 9690 5010 9750
rect 4910 9650 4940 9690
rect 4980 9650 5010 9690
rect 4910 9590 5010 9650
rect 4910 9550 4940 9590
rect 4980 9550 5010 9590
rect 4910 9490 5010 9550
rect 4910 9450 4940 9490
rect 4980 9450 5010 9490
rect 4910 9420 5010 9450
rect 5170 9790 5270 9820
rect 5170 9750 5200 9790
rect 5240 9750 5270 9790
rect 5170 9690 5270 9750
rect 5170 9650 5200 9690
rect 5240 9650 5270 9690
rect 5170 9590 5270 9650
rect 5170 9550 5200 9590
rect 5240 9550 5270 9590
rect 5170 9490 5270 9550
rect 5170 9450 5200 9490
rect 5240 9450 5270 9490
rect 5170 9420 5270 9450
rect 5300 9790 5400 9820
rect 5300 9750 5330 9790
rect 5370 9750 5400 9790
rect 5300 9690 5400 9750
rect 5300 9650 5330 9690
rect 5370 9650 5400 9690
rect 5300 9590 5400 9650
rect 5300 9550 5330 9590
rect 5370 9550 5400 9590
rect 5300 9490 5400 9550
rect 5300 9450 5330 9490
rect 5370 9450 5400 9490
rect 5300 9420 5400 9450
rect 5460 9790 5560 9820
rect 5460 9750 5490 9790
rect 5530 9750 5560 9790
rect 5460 9690 5560 9750
rect 5460 9650 5490 9690
rect 5530 9650 5560 9690
rect 5460 9590 5560 9650
rect 5460 9550 5490 9590
rect 5530 9550 5560 9590
rect 5460 9490 5560 9550
rect 5460 9450 5490 9490
rect 5530 9450 5560 9490
rect 5460 9420 5560 9450
rect 5590 9790 5690 9820
rect 5590 9750 5620 9790
rect 5660 9750 5690 9790
rect 5590 9690 5690 9750
rect 5590 9650 5620 9690
rect 5660 9650 5690 9690
rect 5590 9590 5690 9650
rect 5590 9550 5620 9590
rect 5660 9550 5690 9590
rect 5590 9490 5690 9550
rect 5590 9450 5620 9490
rect 5660 9450 5690 9490
rect 5590 9420 5690 9450
rect 5850 9790 5950 9820
rect 5850 9750 5880 9790
rect 5920 9750 5950 9790
rect 5850 9690 5950 9750
rect 5850 9650 5880 9690
rect 5920 9650 5950 9690
rect 5850 9590 5950 9650
rect 5850 9550 5880 9590
rect 5920 9550 5950 9590
rect 5850 9490 5950 9550
rect 5850 9450 5880 9490
rect 5920 9450 5950 9490
rect 5850 9420 5950 9450
rect 5980 9790 6080 9820
rect 5980 9750 6010 9790
rect 6050 9750 6080 9790
rect 5980 9690 6080 9750
rect 5980 9650 6010 9690
rect 6050 9650 6080 9690
rect 5980 9590 6080 9650
rect 5980 9550 6010 9590
rect 6050 9550 6080 9590
rect 5980 9490 6080 9550
rect 5980 9450 6010 9490
rect 6050 9450 6080 9490
rect 5980 9420 6080 9450
rect 7540 9760 7640 9790
rect 7540 9720 7570 9760
rect 7610 9720 7640 9760
rect 7540 9660 7640 9720
rect 7540 9620 7570 9660
rect 7610 9620 7640 9660
rect 7540 9560 7640 9620
rect 7540 9520 7570 9560
rect 7610 9520 7640 9560
rect 7540 9460 7640 9520
rect 7540 9420 7570 9460
rect 7610 9420 7640 9460
rect 7540 9390 7640 9420
rect 7760 9760 7860 9790
rect 7760 9720 7790 9760
rect 7830 9720 7860 9760
rect 7760 9660 7860 9720
rect 7760 9620 7790 9660
rect 7830 9620 7860 9660
rect 7760 9560 7860 9620
rect 7760 9520 7790 9560
rect 7830 9520 7860 9560
rect 7760 9460 7860 9520
rect 7760 9420 7790 9460
rect 7830 9420 7860 9460
rect 7760 9390 7860 9420
rect 7980 9760 8080 9790
rect 7980 9720 8010 9760
rect 8050 9720 8080 9760
rect 7980 9660 8080 9720
rect 7980 9620 8010 9660
rect 8050 9620 8080 9660
rect 7980 9560 8080 9620
rect 7980 9520 8010 9560
rect 8050 9520 8080 9560
rect 7980 9460 8080 9520
rect 7980 9420 8010 9460
rect 8050 9420 8080 9460
rect 7980 9390 8080 9420
rect 8200 9760 8300 9790
rect 8200 9720 8230 9760
rect 8270 9720 8300 9760
rect 8200 9660 8300 9720
rect 8200 9620 8230 9660
rect 8270 9620 8300 9660
rect 8200 9560 8300 9620
rect 8200 9520 8230 9560
rect 8270 9520 8300 9560
rect 8200 9460 8300 9520
rect 8200 9420 8230 9460
rect 8270 9420 8300 9460
rect 8200 9390 8300 9420
rect 8420 9760 8520 9790
rect 8420 9720 8450 9760
rect 8490 9720 8520 9760
rect 8420 9660 8520 9720
rect 8420 9620 8450 9660
rect 8490 9620 8520 9660
rect 8420 9560 8520 9620
rect 8420 9520 8450 9560
rect 8490 9520 8520 9560
rect 8420 9460 8520 9520
rect 8420 9420 8450 9460
rect 8490 9420 8520 9460
rect 8420 9390 8520 9420
rect 8640 9760 8740 9790
rect 8640 9720 8670 9760
rect 8710 9720 8740 9760
rect 8640 9660 8740 9720
rect 8640 9620 8670 9660
rect 8710 9620 8740 9660
rect 8640 9560 8740 9620
rect 8640 9520 8670 9560
rect 8710 9520 8740 9560
rect 8640 9460 8740 9520
rect 8640 9420 8670 9460
rect 8710 9420 8740 9460
rect 8640 9390 8740 9420
rect 8860 9760 8960 9790
rect 9060 9760 9160 9790
rect 8860 9720 8890 9760
rect 8930 9720 8960 9760
rect 9060 9720 9090 9760
rect 9130 9720 9160 9760
rect 8860 9660 8960 9720
rect 9060 9660 9160 9720
rect 8860 9620 8890 9660
rect 8930 9620 8960 9660
rect 9060 9620 9090 9660
rect 9130 9620 9160 9660
rect 8860 9560 8960 9620
rect 9060 9560 9160 9620
rect 8860 9520 8890 9560
rect 8930 9520 8960 9560
rect 9060 9520 9090 9560
rect 9130 9520 9160 9560
rect 8860 9460 8960 9520
rect 9060 9460 9160 9520
rect 8860 9420 8890 9460
rect 8930 9420 8960 9460
rect 9060 9420 9090 9460
rect 9130 9420 9160 9460
rect 8860 9390 8960 9420
rect 9060 9390 9160 9420
rect 9280 9760 9380 9790
rect 9280 9720 9310 9760
rect 9350 9720 9380 9760
rect 9280 9660 9380 9720
rect 9280 9620 9310 9660
rect 9350 9620 9380 9660
rect 9280 9560 9380 9620
rect 9280 9520 9310 9560
rect 9350 9520 9380 9560
rect 9280 9460 9380 9520
rect 9280 9420 9310 9460
rect 9350 9420 9380 9460
rect 9280 9390 9380 9420
rect 9500 9760 9600 9790
rect 9500 9720 9530 9760
rect 9570 9720 9600 9760
rect 9500 9660 9600 9720
rect 9500 9620 9530 9660
rect 9570 9620 9600 9660
rect 9500 9560 9600 9620
rect 9500 9520 9530 9560
rect 9570 9520 9600 9560
rect 9500 9460 9600 9520
rect 9500 9420 9530 9460
rect 9570 9420 9600 9460
rect 9500 9390 9600 9420
rect 9720 9760 9820 9790
rect 9720 9720 9750 9760
rect 9790 9720 9820 9760
rect 9720 9660 9820 9720
rect 9720 9620 9750 9660
rect 9790 9620 9820 9660
rect 9720 9560 9820 9620
rect 9720 9520 9750 9560
rect 9790 9520 9820 9560
rect 9720 9460 9820 9520
rect 9720 9420 9750 9460
rect 9790 9420 9820 9460
rect 9720 9390 9820 9420
rect 9940 9760 10040 9790
rect 9940 9720 9970 9760
rect 10010 9720 10040 9760
rect 9940 9660 10040 9720
rect 9940 9620 9970 9660
rect 10010 9620 10040 9660
rect 9940 9560 10040 9620
rect 9940 9520 9970 9560
rect 10010 9520 10040 9560
rect 9940 9460 10040 9520
rect 9940 9420 9970 9460
rect 10010 9420 10040 9460
rect 9940 9390 10040 9420
rect 10160 9760 10260 9790
rect 10160 9720 10190 9760
rect 10230 9720 10260 9760
rect 10160 9660 10260 9720
rect 10160 9620 10190 9660
rect 10230 9620 10260 9660
rect 10160 9560 10260 9620
rect 10160 9520 10190 9560
rect 10230 9520 10260 9560
rect 10160 9460 10260 9520
rect 10160 9420 10190 9460
rect 10230 9420 10260 9460
rect 10160 9390 10260 9420
rect 10380 9760 10480 9790
rect 10380 9720 10410 9760
rect 10450 9720 10480 9760
rect 10380 9660 10480 9720
rect 10380 9620 10410 9660
rect 10450 9620 10480 9660
rect 10380 9560 10480 9620
rect 10380 9520 10410 9560
rect 10450 9520 10480 9560
rect 10380 9460 10480 9520
rect 10380 9420 10410 9460
rect 10450 9420 10480 9460
rect 10380 9390 10480 9420
rect 1260 9030 1340 9060
rect 1260 8990 1280 9030
rect 1320 8990 1340 9030
rect 1260 8930 1340 8990
rect 1260 8890 1280 8930
rect 1320 8890 1340 8930
rect 1260 8830 1340 8890
rect 1260 8790 1280 8830
rect 1320 8790 1340 8830
rect 1260 8730 1340 8790
rect 1260 8690 1280 8730
rect 1320 8690 1340 8730
rect 1260 8660 1340 8690
rect 1370 9030 1450 9060
rect 1370 8990 1390 9030
rect 1430 8990 1450 9030
rect 1370 8930 1450 8990
rect 1370 8890 1390 8930
rect 1430 8890 1450 8930
rect 1370 8830 1450 8890
rect 1370 8790 1390 8830
rect 1430 8790 1450 8830
rect 1370 8730 1450 8790
rect 1370 8690 1390 8730
rect 1430 8690 1450 8730
rect 1370 8660 1450 8690
rect 1480 9030 1560 9060
rect 1480 8990 1500 9030
rect 1540 8990 1560 9030
rect 1480 8930 1560 8990
rect 1480 8890 1500 8930
rect 1540 8890 1560 8930
rect 1480 8830 1560 8890
rect 1480 8790 1500 8830
rect 1540 8790 1560 8830
rect 1480 8730 1560 8790
rect 1480 8690 1500 8730
rect 1540 8690 1560 8730
rect 1480 8660 1560 8690
rect 1780 9030 1860 9060
rect 1780 8990 1800 9030
rect 1840 8990 1860 9030
rect 1780 8930 1860 8990
rect 1780 8890 1800 8930
rect 1840 8890 1860 8930
rect 1780 8830 1860 8890
rect 1780 8790 1800 8830
rect 1840 8790 1860 8830
rect 1780 8730 1860 8790
rect 1780 8690 1800 8730
rect 1840 8690 1860 8730
rect 1780 8660 1860 8690
rect 1890 9030 1970 9060
rect 1890 8990 1910 9030
rect 1950 8990 1970 9030
rect 1890 8930 1970 8990
rect 1890 8890 1910 8930
rect 1950 8890 1970 8930
rect 1890 8830 1970 8890
rect 1890 8790 1910 8830
rect 1950 8790 1970 8830
rect 1890 8730 1970 8790
rect 1890 8690 1910 8730
rect 1950 8690 1970 8730
rect 1890 8660 1970 8690
rect 2000 9030 2080 9060
rect 2160 9030 2240 9060
rect 2000 8990 2020 9030
rect 2060 8990 2080 9030
rect 2160 8990 2180 9030
rect 2220 8990 2240 9030
rect 2000 8930 2080 8990
rect 2160 8930 2240 8990
rect 2000 8890 2020 8930
rect 2060 8890 2080 8930
rect 2160 8890 2180 8930
rect 2220 8890 2240 8930
rect 2000 8830 2080 8890
rect 2160 8830 2240 8890
rect 2000 8790 2020 8830
rect 2060 8790 2080 8830
rect 2160 8790 2180 8830
rect 2220 8790 2240 8830
rect 2000 8730 2080 8790
rect 2160 8730 2240 8790
rect 2000 8690 2020 8730
rect 2060 8690 2080 8730
rect 2160 8690 2180 8730
rect 2220 8690 2240 8730
rect 2000 8660 2080 8690
rect 2160 8660 2240 8690
rect 2270 9030 2350 9060
rect 2270 8990 2290 9030
rect 2330 8990 2350 9030
rect 2270 8930 2350 8990
rect 2270 8890 2290 8930
rect 2330 8890 2350 8930
rect 2270 8830 2350 8890
rect 2270 8790 2290 8830
rect 2330 8790 2350 8830
rect 2270 8730 2350 8790
rect 2270 8690 2290 8730
rect 2330 8690 2350 8730
rect 2270 8660 2350 8690
rect 2380 9030 2460 9060
rect 2380 8990 2400 9030
rect 2440 8990 2460 9030
rect 2380 8930 2460 8990
rect 2380 8890 2400 8930
rect 2440 8890 2460 8930
rect 2380 8830 2460 8890
rect 2380 8790 2400 8830
rect 2440 8790 2460 8830
rect 2380 8730 2460 8790
rect 2380 8690 2400 8730
rect 2440 8690 2460 8730
rect 2380 8660 2460 8690
rect 2680 9030 2760 9060
rect 2680 8990 2700 9030
rect 2740 8990 2760 9030
rect 2680 8930 2760 8990
rect 2680 8890 2700 8930
rect 2740 8890 2760 8930
rect 2680 8830 2760 8890
rect 2680 8790 2700 8830
rect 2740 8790 2760 8830
rect 2680 8730 2760 8790
rect 2680 8690 2700 8730
rect 2740 8690 2760 8730
rect 2680 8660 2760 8690
rect 2790 9030 2870 9060
rect 2790 8990 2810 9030
rect 2850 8990 2870 9030
rect 2790 8930 2870 8990
rect 2790 8890 2810 8930
rect 2850 8890 2870 8930
rect 2790 8830 2870 8890
rect 2790 8790 2810 8830
rect 2850 8790 2870 8830
rect 2790 8730 2870 8790
rect 2790 8690 2810 8730
rect 2850 8690 2870 8730
rect 2790 8660 2870 8690
rect 2900 9030 2980 9060
rect 2900 8990 2920 9030
rect 2960 8990 2980 9030
rect 2900 8930 2980 8990
rect 2900 8890 2920 8930
rect 2960 8890 2980 8930
rect 2900 8830 2980 8890
rect 2900 8790 2920 8830
rect 2960 8790 2980 8830
rect 2900 8730 2980 8790
rect 2900 8690 2920 8730
rect 2960 8690 2980 8730
rect 2900 8660 2980 8690
rect 3190 9030 3270 9060
rect 3190 8990 3210 9030
rect 3250 8990 3270 9030
rect 3190 8930 3270 8990
rect 3190 8890 3210 8930
rect 3250 8890 3270 8930
rect 3190 8830 3270 8890
rect 3190 8790 3210 8830
rect 3250 8790 3270 8830
rect 3190 8730 3270 8790
rect 3190 8690 3210 8730
rect 3250 8690 3270 8730
rect 3190 8660 3270 8690
rect 3300 9030 3380 9060
rect 3300 8990 3320 9030
rect 3360 8990 3380 9030
rect 3300 8930 3380 8990
rect 3300 8890 3320 8930
rect 3360 8890 3380 8930
rect 3300 8830 3380 8890
rect 3300 8790 3320 8830
rect 3360 8790 3380 8830
rect 3300 8730 3380 8790
rect 3300 8690 3320 8730
rect 3360 8690 3380 8730
rect 3300 8660 3380 8690
rect 3520 9030 3600 9060
rect 3520 8990 3540 9030
rect 3580 8990 3600 9030
rect 3520 8930 3600 8990
rect 3520 8890 3540 8930
rect 3580 8890 3600 8930
rect 3520 8830 3600 8890
rect 3520 8790 3540 8830
rect 3580 8790 3600 8830
rect 3520 8730 3600 8790
rect 3520 8690 3540 8730
rect 3580 8690 3600 8730
rect 3520 8660 3600 8690
rect 3630 9030 3710 9060
rect 3630 8990 3650 9030
rect 3690 8990 3710 9030
rect 3630 8930 3710 8990
rect 3630 8890 3650 8930
rect 3690 8890 3710 8930
rect 3630 8830 3710 8890
rect 3630 8790 3650 8830
rect 3690 8790 3710 8830
rect 3630 8730 3710 8790
rect 3630 8690 3650 8730
rect 3690 8690 3710 8730
rect 3630 8660 3710 8690
rect 3850 9030 3930 9060
rect 3850 8990 3870 9030
rect 3910 8990 3930 9030
rect 3850 8930 3930 8990
rect 3850 8890 3870 8930
rect 3910 8890 3930 8930
rect 3850 8830 3930 8890
rect 3850 8790 3870 8830
rect 3910 8790 3930 8830
rect 3850 8730 3930 8790
rect 3850 8690 3870 8730
rect 3910 8690 3930 8730
rect 3850 8660 3930 8690
rect 3960 9030 4040 9060
rect 3960 8990 3980 9030
rect 4020 8990 4040 9030
rect 3960 8930 4040 8990
rect 3960 8890 3980 8930
rect 4020 8890 4040 8930
rect 3960 8830 4040 8890
rect 3960 8790 3980 8830
rect 4020 8790 4040 8830
rect 3960 8730 4040 8790
rect 3960 8690 3980 8730
rect 4020 8690 4040 8730
rect 3960 8660 4040 8690
rect 4390 9030 4490 9060
rect 4390 8990 4420 9030
rect 4460 8990 4490 9030
rect 4390 8930 4490 8990
rect 4390 8890 4420 8930
rect 4460 8890 4490 8930
rect 4390 8830 4490 8890
rect 4390 8790 4420 8830
rect 4460 8790 4490 8830
rect 4390 8730 4490 8790
rect 4390 8690 4420 8730
rect 4460 8690 4490 8730
rect 4390 8660 4490 8690
rect 4520 9030 4620 9060
rect 4520 8990 4550 9030
rect 4590 8990 4620 9030
rect 4520 8930 4620 8990
rect 4520 8890 4550 8930
rect 4590 8890 4620 8930
rect 4520 8830 4620 8890
rect 4520 8790 4550 8830
rect 4590 8790 4620 8830
rect 4520 8730 4620 8790
rect 4520 8690 4550 8730
rect 4590 8690 4620 8730
rect 4520 8660 4620 8690
rect 4780 9030 4880 9060
rect 4780 8990 4810 9030
rect 4850 8990 4880 9030
rect 4780 8930 4880 8990
rect 4780 8890 4810 8930
rect 4850 8890 4880 8930
rect 4780 8830 4880 8890
rect 4780 8790 4810 8830
rect 4850 8790 4880 8830
rect 4780 8730 4880 8790
rect 4780 8690 4810 8730
rect 4850 8690 4880 8730
rect 4780 8660 4880 8690
rect 4910 9030 5010 9060
rect 4910 8990 4940 9030
rect 4980 8990 5010 9030
rect 4910 8930 5010 8990
rect 4910 8890 4940 8930
rect 4980 8890 5010 8930
rect 4910 8830 5010 8890
rect 4910 8790 4940 8830
rect 4980 8790 5010 8830
rect 4910 8730 5010 8790
rect 4910 8690 4940 8730
rect 4980 8690 5010 8730
rect 4910 8660 5010 8690
rect 5170 9030 5270 9060
rect 5170 8990 5200 9030
rect 5240 8990 5270 9030
rect 5170 8930 5270 8990
rect 5170 8890 5200 8930
rect 5240 8890 5270 8930
rect 5170 8830 5270 8890
rect 5170 8790 5200 8830
rect 5240 8790 5270 8830
rect 5170 8730 5270 8790
rect 5170 8690 5200 8730
rect 5240 8690 5270 8730
rect 5170 8660 5270 8690
rect 5300 9030 5400 9060
rect 5300 8990 5330 9030
rect 5370 8990 5400 9030
rect 5300 8930 5400 8990
rect 5300 8890 5330 8930
rect 5370 8890 5400 8930
rect 5300 8830 5400 8890
rect 5300 8790 5330 8830
rect 5370 8790 5400 8830
rect 5300 8730 5400 8790
rect 5300 8690 5330 8730
rect 5370 8690 5400 8730
rect 5300 8660 5400 8690
rect 5460 9030 5560 9060
rect 5460 8990 5490 9030
rect 5530 8990 5560 9030
rect 5460 8930 5560 8990
rect 5460 8890 5490 8930
rect 5530 8890 5560 8930
rect 5460 8830 5560 8890
rect 5460 8790 5490 8830
rect 5530 8790 5560 8830
rect 5460 8730 5560 8790
rect 5460 8690 5490 8730
rect 5530 8690 5560 8730
rect 5460 8660 5560 8690
rect 5590 9030 5690 9060
rect 5590 8990 5620 9030
rect 5660 8990 5690 9030
rect 5590 8930 5690 8990
rect 5590 8890 5620 8930
rect 5660 8890 5690 8930
rect 5590 8830 5690 8890
rect 5590 8790 5620 8830
rect 5660 8790 5690 8830
rect 5590 8730 5690 8790
rect 5590 8690 5620 8730
rect 5660 8690 5690 8730
rect 5590 8660 5690 8690
rect -360 6840 -280 6870
rect -360 6800 -340 6840
rect -300 6800 -280 6840
rect -360 6740 -280 6800
rect -360 6700 -340 6740
rect -300 6700 -280 6740
rect -360 6670 -280 6700
rect -250 6840 -170 6870
rect -250 6800 -230 6840
rect -190 6800 -170 6840
rect -250 6740 -170 6800
rect -250 6700 -230 6740
rect -190 6700 -170 6740
rect -250 6670 -170 6700
rect -140 6840 -60 6870
rect -140 6800 -120 6840
rect -80 6800 -60 6840
rect -140 6740 -60 6800
rect -140 6700 -120 6740
rect -80 6700 -60 6740
rect -140 6670 -60 6700
rect -30 6840 50 6870
rect -30 6800 -10 6840
rect 30 6800 50 6840
rect -30 6740 50 6800
rect -30 6700 -10 6740
rect 30 6700 50 6740
rect -30 6670 50 6700
rect 80 6840 160 6870
rect 80 6800 100 6840
rect 140 6800 160 6840
rect 80 6740 160 6800
rect 80 6700 100 6740
rect 140 6700 160 6740
rect 80 6670 160 6700
rect 190 6840 270 6870
rect 190 6800 210 6840
rect 250 6800 270 6840
rect 190 6740 270 6800
rect 190 6700 210 6740
rect 250 6700 270 6740
rect 190 6670 270 6700
rect 300 6840 380 6870
rect 300 6800 320 6840
rect 360 6800 380 6840
rect 300 6740 380 6800
rect 300 6700 320 6740
rect 360 6700 380 6740
rect 300 6670 380 6700
rect 410 6840 490 6870
rect 410 6800 430 6840
rect 470 6800 490 6840
rect 410 6740 490 6800
rect 410 6700 430 6740
rect 470 6700 490 6740
rect 410 6670 490 6700
rect 520 6840 600 6870
rect 520 6800 540 6840
rect 580 6800 600 6840
rect 520 6740 600 6800
rect 520 6700 540 6740
rect 580 6700 600 6740
rect 520 6670 600 6700
rect 630 6840 710 6870
rect 630 6800 650 6840
rect 690 6800 710 6840
rect 630 6740 710 6800
rect 630 6700 650 6740
rect 690 6700 710 6740
rect 630 6670 710 6700
rect 740 6840 820 6870
rect 740 6800 760 6840
rect 800 6800 820 6840
rect 740 6740 820 6800
rect 740 6700 760 6740
rect 800 6700 820 6740
rect 740 6670 820 6700
rect 850 6840 930 6870
rect 850 6800 870 6840
rect 910 6800 930 6840
rect 850 6740 930 6800
rect 850 6700 870 6740
rect 910 6700 930 6740
rect 850 6670 930 6700
rect 960 6840 1040 6870
rect 960 6800 980 6840
rect 1020 6800 1040 6840
rect 960 6740 1040 6800
rect 960 6700 980 6740
rect 1020 6700 1040 6740
rect 960 6670 1040 6700
rect 1540 6840 1620 6870
rect 1540 6800 1560 6840
rect 1600 6800 1620 6840
rect 1540 6740 1620 6800
rect 1540 6700 1560 6740
rect 1600 6700 1620 6740
rect 1540 6670 1620 6700
rect 1650 6840 1730 6870
rect 1650 6800 1670 6840
rect 1710 6800 1730 6840
rect 1650 6740 1730 6800
rect 1650 6700 1670 6740
rect 1710 6700 1730 6740
rect 1650 6670 1730 6700
rect 1760 6840 1840 6870
rect 1760 6800 1780 6840
rect 1820 6800 1840 6840
rect 1760 6740 1840 6800
rect 1760 6700 1780 6740
rect 1820 6700 1840 6740
rect 1760 6670 1840 6700
rect 1870 6840 1950 6870
rect 1870 6800 1890 6840
rect 1930 6800 1950 6840
rect 1870 6740 1950 6800
rect 1870 6700 1890 6740
rect 1930 6700 1950 6740
rect 1870 6670 1950 6700
rect 1980 6840 2060 6870
rect 1980 6800 2000 6840
rect 2040 6800 2060 6840
rect 1980 6740 2060 6800
rect 1980 6700 2000 6740
rect 2040 6700 2060 6740
rect 1980 6670 2060 6700
rect 2090 6840 2170 6870
rect 2090 6800 2110 6840
rect 2150 6800 2170 6840
rect 2090 6740 2170 6800
rect 2090 6700 2110 6740
rect 2150 6700 2170 6740
rect 2090 6670 2170 6700
rect 2200 6840 2280 6870
rect 2200 6800 2220 6840
rect 2260 6800 2280 6840
rect 2200 6740 2280 6800
rect 2200 6700 2220 6740
rect 2260 6700 2280 6740
rect 2200 6670 2280 6700
rect 2310 6840 2390 6870
rect 2310 6800 2330 6840
rect 2370 6800 2390 6840
rect 2310 6740 2390 6800
rect 2310 6700 2330 6740
rect 2370 6700 2390 6740
rect 2310 6670 2390 6700
rect 2420 6840 2500 6870
rect 2420 6800 2440 6840
rect 2480 6800 2500 6840
rect 2420 6740 2500 6800
rect 2420 6700 2440 6740
rect 2480 6700 2500 6740
rect 2420 6670 2500 6700
rect 2530 6840 2610 6870
rect 2530 6800 2550 6840
rect 2590 6800 2610 6840
rect 2530 6740 2610 6800
rect 2530 6700 2550 6740
rect 2590 6700 2610 6740
rect 2530 6670 2610 6700
rect 2640 6840 2720 6870
rect 2640 6800 2660 6840
rect 2700 6800 2720 6840
rect 2640 6740 2720 6800
rect 2640 6700 2660 6740
rect 2700 6700 2720 6740
rect 2640 6670 2720 6700
rect 2750 6840 2830 6870
rect 2750 6800 2770 6840
rect 2810 6800 2830 6840
rect 2750 6740 2830 6800
rect 2750 6700 2770 6740
rect 2810 6700 2830 6740
rect 2750 6670 2830 6700
rect 2860 6840 2940 6870
rect 2860 6800 2880 6840
rect 2920 6800 2940 6840
rect 2860 6740 2940 6800
rect 2860 6700 2880 6740
rect 2920 6700 2940 6740
rect 2860 6670 2940 6700
rect -370 6240 -290 6270
rect -370 6200 -350 6240
rect -310 6200 -290 6240
rect -370 6140 -290 6200
rect -370 6100 -350 6140
rect -310 6100 -290 6140
rect -370 6040 -290 6100
rect -370 6000 -350 6040
rect -310 6000 -290 6040
rect -370 5940 -290 6000
rect -370 5900 -350 5940
rect -310 5900 -290 5940
rect -370 5840 -290 5900
rect -370 5800 -350 5840
rect -310 5800 -290 5840
rect -370 5740 -290 5800
rect -370 5700 -350 5740
rect -310 5700 -290 5740
rect -370 5670 -290 5700
rect -190 6240 -110 6270
rect -190 6200 -170 6240
rect -130 6200 -110 6240
rect -190 6140 -110 6200
rect -190 6100 -170 6140
rect -130 6100 -110 6140
rect -190 6040 -110 6100
rect -190 6000 -170 6040
rect -130 6000 -110 6040
rect -190 5940 -110 6000
rect -190 5900 -170 5940
rect -130 5900 -110 5940
rect -190 5840 -110 5900
rect -190 5800 -170 5840
rect -130 5800 -110 5840
rect -190 5740 -110 5800
rect -190 5700 -170 5740
rect -130 5700 -110 5740
rect -190 5670 -110 5700
rect -10 6240 70 6270
rect -10 6200 10 6240
rect 50 6200 70 6240
rect -10 6140 70 6200
rect -10 6100 10 6140
rect 50 6100 70 6140
rect -10 6040 70 6100
rect -10 6000 10 6040
rect 50 6000 70 6040
rect -10 5940 70 6000
rect -10 5900 10 5940
rect 50 5900 70 5940
rect -10 5840 70 5900
rect -10 5800 10 5840
rect 50 5800 70 5840
rect -10 5740 70 5800
rect -10 5700 10 5740
rect 50 5700 70 5740
rect -10 5670 70 5700
rect 170 6240 250 6270
rect 170 6200 190 6240
rect 230 6200 250 6240
rect 170 6140 250 6200
rect 170 6100 190 6140
rect 230 6100 250 6140
rect 170 6040 250 6100
rect 170 6000 190 6040
rect 230 6000 250 6040
rect 170 5940 250 6000
rect 170 5900 190 5940
rect 230 5900 250 5940
rect 170 5840 250 5900
rect 170 5800 190 5840
rect 230 5800 250 5840
rect 170 5740 250 5800
rect 170 5700 190 5740
rect 230 5700 250 5740
rect 170 5670 250 5700
rect 350 6240 430 6270
rect 350 6200 370 6240
rect 410 6200 430 6240
rect 350 6140 430 6200
rect 350 6100 370 6140
rect 410 6100 430 6140
rect 350 6040 430 6100
rect 350 6000 370 6040
rect 410 6000 430 6040
rect 350 5940 430 6000
rect 350 5900 370 5940
rect 410 5900 430 5940
rect 350 5840 430 5900
rect 350 5800 370 5840
rect 410 5800 430 5840
rect 350 5740 430 5800
rect 350 5700 370 5740
rect 410 5700 430 5740
rect 350 5670 430 5700
rect 530 6240 610 6270
rect 530 6200 550 6240
rect 590 6200 610 6240
rect 530 6140 610 6200
rect 530 6100 550 6140
rect 590 6100 610 6140
rect 530 6040 610 6100
rect 530 6000 550 6040
rect 590 6000 610 6040
rect 530 5940 610 6000
rect 530 5900 550 5940
rect 590 5900 610 5940
rect 530 5840 610 5900
rect 530 5800 550 5840
rect 590 5800 610 5840
rect 530 5740 610 5800
rect 530 5700 550 5740
rect 590 5700 610 5740
rect 530 5670 610 5700
rect 710 6240 790 6270
rect 710 6200 730 6240
rect 770 6200 790 6240
rect 710 6140 790 6200
rect 710 6100 730 6140
rect 770 6100 790 6140
rect 710 6040 790 6100
rect 710 6000 730 6040
rect 770 6000 790 6040
rect 710 5940 790 6000
rect 710 5900 730 5940
rect 770 5900 790 5940
rect 710 5840 790 5900
rect 710 5800 730 5840
rect 770 5800 790 5840
rect 710 5740 790 5800
rect 710 5700 730 5740
rect 770 5700 790 5740
rect 710 5670 790 5700
rect 890 6240 970 6270
rect 890 6200 910 6240
rect 950 6200 970 6240
rect 890 6140 970 6200
rect 890 6100 910 6140
rect 950 6100 970 6140
rect 890 6040 970 6100
rect 890 6000 910 6040
rect 950 6000 970 6040
rect 890 5940 970 6000
rect 890 5900 910 5940
rect 950 5900 970 5940
rect 890 5840 970 5900
rect 890 5800 910 5840
rect 950 5800 970 5840
rect 890 5740 970 5800
rect 890 5700 910 5740
rect 950 5700 970 5740
rect 890 5670 970 5700
rect 1070 6240 1150 6270
rect 1070 6200 1090 6240
rect 1130 6200 1150 6240
rect 1070 6140 1150 6200
rect 1070 6100 1090 6140
rect 1130 6100 1150 6140
rect 1070 6040 1150 6100
rect 1070 6000 1090 6040
rect 1130 6000 1150 6040
rect 1070 5940 1150 6000
rect 1070 5900 1090 5940
rect 1130 5900 1150 5940
rect 1070 5840 1150 5900
rect 1070 5800 1090 5840
rect 1130 5800 1150 5840
rect 1070 5740 1150 5800
rect 1070 5700 1090 5740
rect 1130 5700 1150 5740
rect 1070 5670 1150 5700
rect 1250 6240 1330 6270
rect 1250 6200 1270 6240
rect 1310 6200 1330 6240
rect 1250 6140 1330 6200
rect 1250 6100 1270 6140
rect 1310 6100 1330 6140
rect 1250 6040 1330 6100
rect 1250 6000 1270 6040
rect 1310 6000 1330 6040
rect 1250 5940 1330 6000
rect 1250 5900 1270 5940
rect 1310 5900 1330 5940
rect 1250 5840 1330 5900
rect 1250 5800 1270 5840
rect 1310 5800 1330 5840
rect 1250 5740 1330 5800
rect 1250 5700 1270 5740
rect 1310 5700 1330 5740
rect 1250 5670 1330 5700
rect 1430 6240 1510 6270
rect 1430 6200 1450 6240
rect 1490 6200 1510 6240
rect 1430 6140 1510 6200
rect 1430 6100 1450 6140
rect 1490 6100 1510 6140
rect 1430 6040 1510 6100
rect 1430 6000 1450 6040
rect 1490 6000 1510 6040
rect 1430 5940 1510 6000
rect 1430 5900 1450 5940
rect 1490 5900 1510 5940
rect 1430 5840 1510 5900
rect 1430 5800 1450 5840
rect 1490 5800 1510 5840
rect 1430 5740 1510 5800
rect 1430 5700 1450 5740
rect 1490 5700 1510 5740
rect 1430 5670 1510 5700
rect 1610 6240 1690 6270
rect 1610 6200 1630 6240
rect 1670 6200 1690 6240
rect 1610 6140 1690 6200
rect 1610 6100 1630 6140
rect 1670 6100 1690 6140
rect 1610 6040 1690 6100
rect 1610 6000 1630 6040
rect 1670 6000 1690 6040
rect 1610 5940 1690 6000
rect 1610 5900 1630 5940
rect 1670 5900 1690 5940
rect 1610 5840 1690 5900
rect 1610 5800 1630 5840
rect 1670 5800 1690 5840
rect 1610 5740 1690 5800
rect 1610 5700 1630 5740
rect 1670 5700 1690 5740
rect 1610 5670 1690 5700
rect 1790 6240 1870 6270
rect 1790 6200 1810 6240
rect 1850 6200 1870 6240
rect 1790 6140 1870 6200
rect 1790 6100 1810 6140
rect 1850 6100 1870 6140
rect 1790 6040 1870 6100
rect 1790 6000 1810 6040
rect 1850 6000 1870 6040
rect 1790 5940 1870 6000
rect 1790 5900 1810 5940
rect 1850 5900 1870 5940
rect 1790 5840 1870 5900
rect 1790 5800 1810 5840
rect 1850 5800 1870 5840
rect 1790 5740 1870 5800
rect 1790 5700 1810 5740
rect 1850 5700 1870 5740
rect 1790 5670 1870 5700
rect 1970 6240 2050 6270
rect 1970 6200 1990 6240
rect 2030 6200 2050 6240
rect 1970 6140 2050 6200
rect 1970 6100 1990 6140
rect 2030 6100 2050 6140
rect 1970 6040 2050 6100
rect 1970 6000 1990 6040
rect 2030 6000 2050 6040
rect 1970 5940 2050 6000
rect 1970 5900 1990 5940
rect 2030 5900 2050 5940
rect 1970 5840 2050 5900
rect 1970 5800 1990 5840
rect 2030 5800 2050 5840
rect 1970 5740 2050 5800
rect 1970 5700 1990 5740
rect 2030 5700 2050 5740
rect 1970 5670 2050 5700
rect 2150 6240 2230 6270
rect 2150 6200 2170 6240
rect 2210 6200 2230 6240
rect 2150 6140 2230 6200
rect 2150 6100 2170 6140
rect 2210 6100 2230 6140
rect 2150 6040 2230 6100
rect 2150 6000 2170 6040
rect 2210 6000 2230 6040
rect 2150 5940 2230 6000
rect 2150 5900 2170 5940
rect 2210 5900 2230 5940
rect 2150 5840 2230 5900
rect 2150 5800 2170 5840
rect 2210 5800 2230 5840
rect 2150 5740 2230 5800
rect 2150 5700 2170 5740
rect 2210 5700 2230 5740
rect 2150 5670 2230 5700
rect 2330 6240 2410 6270
rect 2330 6200 2350 6240
rect 2390 6200 2410 6240
rect 2330 6140 2410 6200
rect 2330 6100 2350 6140
rect 2390 6100 2410 6140
rect 2330 6040 2410 6100
rect 2330 6000 2350 6040
rect 2390 6000 2410 6040
rect 2330 5940 2410 6000
rect 2330 5900 2350 5940
rect 2390 5900 2410 5940
rect 2330 5840 2410 5900
rect 2330 5800 2350 5840
rect 2390 5800 2410 5840
rect 2330 5740 2410 5800
rect 2330 5700 2350 5740
rect 2390 5700 2410 5740
rect 2330 5670 2410 5700
rect 2510 6240 2590 6270
rect 2510 6200 2530 6240
rect 2570 6200 2590 6240
rect 2510 6140 2590 6200
rect 2510 6100 2530 6140
rect 2570 6100 2590 6140
rect 2510 6040 2590 6100
rect 2510 6000 2530 6040
rect 2570 6000 2590 6040
rect 2510 5940 2590 6000
rect 2510 5900 2530 5940
rect 2570 5900 2590 5940
rect 2510 5840 2590 5900
rect 2510 5800 2530 5840
rect 2570 5800 2590 5840
rect 2510 5740 2590 5800
rect 2510 5700 2530 5740
rect 2570 5700 2590 5740
rect 2510 5670 2590 5700
rect 2690 6240 2770 6270
rect 2690 6200 2710 6240
rect 2750 6200 2770 6240
rect 2690 6140 2770 6200
rect 2690 6100 2710 6140
rect 2750 6100 2770 6140
rect 2690 6040 2770 6100
rect 2690 6000 2710 6040
rect 2750 6000 2770 6040
rect 2690 5940 2770 6000
rect 2690 5900 2710 5940
rect 2750 5900 2770 5940
rect 2690 5840 2770 5900
rect 2690 5800 2710 5840
rect 2750 5800 2770 5840
rect 2690 5740 2770 5800
rect 2690 5700 2710 5740
rect 2750 5700 2770 5740
rect 2690 5670 2770 5700
rect 2870 6240 2950 6270
rect 2870 6200 2890 6240
rect 2930 6200 2950 6240
rect 2870 6140 2950 6200
rect 2870 6100 2890 6140
rect 2930 6100 2950 6140
rect 2870 6040 2950 6100
rect 2870 6000 2890 6040
rect 2930 6000 2950 6040
rect 2870 5940 2950 6000
rect 2870 5900 2890 5940
rect 2930 5900 2950 5940
rect 2870 5840 2950 5900
rect 3490 6040 3580 6070
rect 3490 6000 3520 6040
rect 3560 6000 3580 6040
rect 3490 5940 3580 6000
rect 3490 5900 3520 5940
rect 3560 5900 3580 5940
rect 3490 5870 3580 5900
rect 3610 6040 3690 6070
rect 3610 6000 3630 6040
rect 3670 6000 3690 6040
rect 3610 5940 3690 6000
rect 3610 5900 3630 5940
rect 3670 5900 3690 5940
rect 3610 5870 3690 5900
rect 3720 6040 3800 6070
rect 3720 6000 3740 6040
rect 3780 6000 3800 6040
rect 3720 5940 3800 6000
rect 3720 5900 3740 5940
rect 3780 5900 3800 5940
rect 3720 5870 3800 5900
rect 3830 6040 3910 6070
rect 3830 6000 3850 6040
rect 3890 6000 3910 6040
rect 3830 5940 3910 6000
rect 3830 5900 3850 5940
rect 3890 5900 3910 5940
rect 3830 5870 3910 5900
rect 3940 6040 4020 6070
rect 3940 6000 3960 6040
rect 4000 6000 4020 6040
rect 3940 5940 4020 6000
rect 3940 5900 3960 5940
rect 4000 5900 4020 5940
rect 3940 5870 4020 5900
rect 2870 5800 2890 5840
rect 2930 5800 2950 5840
rect 2870 5740 2950 5800
rect 2870 5700 2890 5740
rect 2930 5700 2950 5740
rect 2870 5670 2950 5700
rect 7450 4760 7550 4790
rect 7450 4720 7480 4760
rect 7520 4720 7550 4760
rect -1470 4680 -1390 4710
rect -1470 4640 -1450 4680
rect -1410 4640 -1390 4680
rect -1470 4580 -1390 4640
rect -1470 4540 -1450 4580
rect -1410 4540 -1390 4580
rect -1470 4510 -1390 4540
rect -1350 4680 -1270 4710
rect -1350 4640 -1330 4680
rect -1290 4640 -1270 4680
rect -1350 4580 -1270 4640
rect -1350 4540 -1330 4580
rect -1290 4540 -1270 4580
rect -1350 4510 -1270 4540
rect -1230 4680 -1150 4710
rect -1230 4640 -1210 4680
rect -1170 4640 -1150 4680
rect -1230 4580 -1150 4640
rect -1230 4540 -1210 4580
rect -1170 4540 -1150 4580
rect -1230 4510 -1150 4540
rect -1110 4680 -1030 4710
rect -1110 4640 -1090 4680
rect -1050 4640 -1030 4680
rect -1110 4580 -1030 4640
rect -1110 4540 -1090 4580
rect -1050 4540 -1030 4580
rect -1110 4510 -1030 4540
rect -990 4680 -910 4710
rect -990 4640 -970 4680
rect -930 4640 -910 4680
rect -990 4580 -910 4640
rect -990 4540 -970 4580
rect -930 4540 -910 4580
rect -990 4510 -910 4540
rect -870 4680 -790 4710
rect -870 4640 -850 4680
rect -810 4640 -790 4680
rect -870 4580 -790 4640
rect -870 4540 -850 4580
rect -810 4540 -790 4580
rect -870 4510 -790 4540
rect -750 4680 -670 4710
rect -750 4640 -730 4680
rect -690 4640 -670 4680
rect -750 4580 -670 4640
rect -750 4540 -730 4580
rect -690 4540 -670 4580
rect -750 4510 -670 4540
rect -630 4680 -550 4710
rect -630 4640 -610 4680
rect -570 4640 -550 4680
rect -630 4580 -550 4640
rect -630 4540 -610 4580
rect -570 4540 -550 4580
rect -630 4510 -550 4540
rect -510 4680 -430 4710
rect -510 4640 -490 4680
rect -450 4640 -430 4680
rect -510 4580 -430 4640
rect -510 4540 -490 4580
rect -450 4540 -430 4580
rect -510 4510 -430 4540
rect -390 4680 -310 4710
rect -390 4640 -370 4680
rect -330 4640 -310 4680
rect -390 4580 -310 4640
rect -390 4540 -370 4580
rect -330 4540 -310 4580
rect -390 4510 -310 4540
rect -270 4680 -190 4710
rect -270 4640 -250 4680
rect -210 4640 -190 4680
rect -270 4580 -190 4640
rect -270 4540 -250 4580
rect -210 4540 -190 4580
rect -270 4510 -190 4540
rect -150 4680 -70 4710
rect -150 4640 -130 4680
rect -90 4640 -70 4680
rect -150 4580 -70 4640
rect -150 4540 -130 4580
rect -90 4540 -70 4580
rect -150 4510 -70 4540
rect -30 4680 50 4710
rect -30 4640 -10 4680
rect 30 4640 50 4680
rect -30 4580 50 4640
rect -30 4540 -10 4580
rect 30 4540 50 4580
rect -30 4510 50 4540
rect 90 4680 170 4710
rect 90 4640 110 4680
rect 150 4640 170 4680
rect 90 4580 170 4640
rect 90 4540 110 4580
rect 150 4540 170 4580
rect 90 4510 170 4540
rect 210 4680 290 4710
rect 210 4640 230 4680
rect 270 4640 290 4680
rect 210 4580 290 4640
rect 210 4540 230 4580
rect 270 4540 290 4580
rect 210 4510 290 4540
rect 330 4680 410 4710
rect 330 4640 350 4680
rect 390 4640 410 4680
rect 330 4580 410 4640
rect 330 4540 350 4580
rect 390 4540 410 4580
rect 330 4510 410 4540
rect 450 4680 530 4710
rect 450 4640 470 4680
rect 510 4640 530 4680
rect 450 4580 530 4640
rect 450 4540 470 4580
rect 510 4540 530 4580
rect 450 4510 530 4540
rect 570 4680 650 4710
rect 570 4640 590 4680
rect 630 4640 650 4680
rect 570 4580 650 4640
rect 570 4540 590 4580
rect 630 4540 650 4580
rect 570 4510 650 4540
rect 690 4680 770 4710
rect 690 4640 710 4680
rect 750 4640 770 4680
rect 690 4580 770 4640
rect 690 4540 710 4580
rect 750 4540 770 4580
rect 690 4510 770 4540
rect 810 4680 890 4710
rect 810 4640 830 4680
rect 870 4640 890 4680
rect 810 4580 890 4640
rect 810 4540 830 4580
rect 870 4540 890 4580
rect 810 4510 890 4540
rect 930 4680 1010 4710
rect 930 4640 950 4680
rect 990 4640 1010 4680
rect 930 4580 1010 4640
rect 930 4540 950 4580
rect 990 4540 1010 4580
rect 930 4510 1010 4540
rect 1570 4680 1650 4710
rect 1570 4640 1590 4680
rect 1630 4640 1650 4680
rect 1570 4580 1650 4640
rect 1570 4540 1590 4580
rect 1630 4540 1650 4580
rect 1570 4510 1650 4540
rect 1690 4680 1770 4710
rect 1690 4640 1710 4680
rect 1750 4640 1770 4680
rect 1690 4580 1770 4640
rect 1690 4540 1710 4580
rect 1750 4540 1770 4580
rect 1690 4510 1770 4540
rect 1810 4680 1890 4710
rect 1810 4640 1830 4680
rect 1870 4640 1890 4680
rect 1810 4580 1890 4640
rect 1810 4540 1830 4580
rect 1870 4540 1890 4580
rect 1810 4510 1890 4540
rect 1930 4680 2010 4710
rect 1930 4640 1950 4680
rect 1990 4640 2010 4680
rect 1930 4580 2010 4640
rect 1930 4540 1950 4580
rect 1990 4540 2010 4580
rect 1930 4510 2010 4540
rect 2050 4680 2130 4710
rect 2050 4640 2070 4680
rect 2110 4640 2130 4680
rect 2050 4580 2130 4640
rect 2050 4540 2070 4580
rect 2110 4540 2130 4580
rect 2050 4510 2130 4540
rect 2170 4680 2250 4710
rect 2170 4640 2190 4680
rect 2230 4640 2250 4680
rect 2170 4580 2250 4640
rect 2170 4540 2190 4580
rect 2230 4540 2250 4580
rect 2170 4510 2250 4540
rect 2290 4680 2370 4710
rect 2290 4640 2310 4680
rect 2350 4640 2370 4680
rect 2290 4580 2370 4640
rect 2290 4540 2310 4580
rect 2350 4540 2370 4580
rect 2290 4510 2370 4540
rect 2410 4680 2490 4710
rect 2410 4640 2430 4680
rect 2470 4640 2490 4680
rect 2410 4580 2490 4640
rect 2410 4540 2430 4580
rect 2470 4540 2490 4580
rect 2410 4510 2490 4540
rect 2530 4680 2610 4710
rect 2530 4640 2550 4680
rect 2590 4640 2610 4680
rect 2530 4580 2610 4640
rect 2530 4540 2550 4580
rect 2590 4540 2610 4580
rect 2530 4510 2610 4540
rect 2650 4680 2730 4710
rect 2650 4640 2670 4680
rect 2710 4640 2730 4680
rect 2650 4580 2730 4640
rect 2650 4540 2670 4580
rect 2710 4540 2730 4580
rect 2650 4510 2730 4540
rect 2770 4680 2850 4710
rect 2770 4640 2790 4680
rect 2830 4640 2850 4680
rect 2770 4580 2850 4640
rect 2770 4540 2790 4580
rect 2830 4540 2850 4580
rect 2770 4510 2850 4540
rect 2890 4680 2970 4710
rect 2890 4640 2910 4680
rect 2950 4640 2970 4680
rect 2890 4580 2970 4640
rect 2890 4540 2910 4580
rect 2950 4540 2970 4580
rect 2890 4510 2970 4540
rect 3010 4680 3090 4710
rect 3010 4640 3030 4680
rect 3070 4640 3090 4680
rect 3010 4580 3090 4640
rect 3010 4540 3030 4580
rect 3070 4540 3090 4580
rect 3010 4510 3090 4540
rect 3130 4680 3210 4710
rect 3130 4640 3150 4680
rect 3190 4640 3210 4680
rect 3130 4580 3210 4640
rect 3130 4540 3150 4580
rect 3190 4540 3210 4580
rect 3130 4510 3210 4540
rect 3250 4680 3330 4710
rect 3250 4640 3270 4680
rect 3310 4640 3330 4680
rect 3250 4580 3330 4640
rect 3250 4540 3270 4580
rect 3310 4540 3330 4580
rect 3250 4510 3330 4540
rect 3370 4680 3450 4710
rect 3370 4640 3390 4680
rect 3430 4640 3450 4680
rect 3370 4580 3450 4640
rect 3370 4540 3390 4580
rect 3430 4540 3450 4580
rect 3370 4510 3450 4540
rect 3490 4680 3570 4710
rect 3490 4640 3510 4680
rect 3550 4640 3570 4680
rect 3490 4580 3570 4640
rect 3490 4540 3510 4580
rect 3550 4540 3570 4580
rect 3490 4510 3570 4540
rect 3610 4680 3690 4710
rect 3610 4640 3630 4680
rect 3670 4640 3690 4680
rect 3610 4580 3690 4640
rect 3610 4540 3630 4580
rect 3670 4540 3690 4580
rect 3610 4510 3690 4540
rect 3730 4680 3810 4710
rect 3730 4640 3750 4680
rect 3790 4640 3810 4680
rect 3730 4580 3810 4640
rect 3730 4540 3750 4580
rect 3790 4540 3810 4580
rect 3730 4510 3810 4540
rect 3850 4680 3930 4710
rect 3850 4640 3870 4680
rect 3910 4640 3930 4680
rect 3850 4580 3930 4640
rect 3850 4540 3870 4580
rect 3910 4540 3930 4580
rect 3850 4510 3930 4540
rect 3970 4680 4050 4710
rect 3970 4640 3990 4680
rect 4030 4640 4050 4680
rect 3970 4580 4050 4640
rect 7450 4660 7550 4720
rect 7450 4620 7480 4660
rect 7520 4620 7550 4660
rect 7450 4590 7550 4620
rect 7580 4760 7680 4790
rect 7580 4720 7610 4760
rect 7650 4720 7680 4760
rect 7580 4660 7680 4720
rect 7580 4620 7610 4660
rect 7650 4620 7680 4660
rect 7580 4590 7680 4620
rect 7710 4760 7810 4790
rect 7710 4720 7740 4760
rect 7780 4720 7810 4760
rect 7710 4660 7810 4720
rect 7710 4620 7740 4660
rect 7780 4620 7810 4660
rect 7710 4590 7810 4620
rect 7840 4760 7940 4790
rect 7840 4720 7870 4760
rect 7910 4720 7940 4760
rect 7840 4660 7940 4720
rect 7840 4620 7870 4660
rect 7910 4620 7940 4660
rect 7840 4590 7940 4620
rect 7970 4760 8070 4790
rect 7970 4720 8000 4760
rect 8040 4720 8070 4760
rect 7970 4660 8070 4720
rect 7970 4620 8000 4660
rect 8040 4620 8070 4660
rect 7970 4590 8070 4620
rect 8100 4760 8200 4790
rect 8100 4720 8130 4760
rect 8170 4720 8200 4760
rect 8100 4660 8200 4720
rect 8100 4620 8130 4660
rect 8170 4620 8200 4660
rect 8100 4590 8200 4620
rect 8230 4760 8330 4790
rect 8230 4720 8260 4760
rect 8300 4720 8330 4760
rect 8230 4660 8330 4720
rect 8230 4620 8260 4660
rect 8300 4620 8330 4660
rect 8230 4590 8330 4620
rect 8590 4760 8690 4790
rect 8590 4720 8620 4760
rect 8660 4720 8690 4760
rect 8590 4660 8690 4720
rect 8590 4620 8620 4660
rect 8660 4620 8690 4660
rect 8590 4590 8690 4620
rect 8720 4760 8820 4790
rect 8720 4720 8750 4760
rect 8790 4720 8820 4760
rect 8720 4660 8820 4720
rect 8720 4620 8750 4660
rect 8790 4620 8820 4660
rect 8720 4590 8820 4620
rect 8850 4760 8950 4790
rect 8850 4720 8880 4760
rect 8920 4720 8950 4760
rect 8850 4660 8950 4720
rect 8850 4620 8880 4660
rect 8920 4620 8950 4660
rect 8850 4590 8950 4620
rect 8980 4760 9080 4790
rect 8980 4720 9010 4760
rect 9050 4720 9080 4760
rect 8980 4660 9080 4720
rect 8980 4620 9010 4660
rect 9050 4620 9080 4660
rect 8980 4590 9080 4620
rect 9110 4760 9210 4790
rect 9110 4720 9140 4760
rect 9180 4720 9210 4760
rect 9110 4660 9210 4720
rect 9110 4620 9140 4660
rect 9180 4620 9210 4660
rect 9110 4590 9210 4620
rect 9240 4760 9340 4790
rect 9240 4720 9270 4760
rect 9310 4720 9340 4760
rect 9240 4660 9340 4720
rect 9240 4620 9270 4660
rect 9310 4620 9340 4660
rect 9240 4590 9340 4620
rect 9370 4760 9470 4790
rect 9370 4720 9400 4760
rect 9440 4720 9470 4760
rect 9370 4660 9470 4720
rect 9370 4620 9400 4660
rect 9440 4620 9470 4660
rect 9370 4590 9470 4620
rect 9730 4760 9830 4790
rect 9730 4720 9760 4760
rect 9800 4720 9830 4760
rect 9730 4660 9830 4720
rect 9730 4620 9760 4660
rect 9800 4620 9830 4660
rect 9730 4590 9830 4620
rect 9860 4760 9960 4790
rect 9860 4720 9890 4760
rect 9930 4720 9960 4760
rect 9860 4660 9960 4720
rect 9860 4620 9890 4660
rect 9930 4620 9960 4660
rect 9860 4590 9960 4620
rect 9990 4760 10090 4790
rect 9990 4720 10020 4760
rect 10060 4720 10090 4760
rect 9990 4660 10090 4720
rect 9990 4620 10020 4660
rect 10060 4620 10090 4660
rect 9990 4590 10090 4620
rect 10120 4760 10220 4790
rect 10120 4720 10150 4760
rect 10190 4720 10220 4760
rect 10120 4660 10220 4720
rect 10120 4620 10150 4660
rect 10190 4620 10220 4660
rect 10120 4590 10220 4620
rect 10250 4760 10350 4790
rect 10250 4720 10280 4760
rect 10320 4720 10350 4760
rect 10250 4660 10350 4720
rect 10250 4620 10280 4660
rect 10320 4620 10350 4660
rect 10250 4590 10350 4620
rect 10380 4760 10480 4790
rect 10380 4720 10410 4760
rect 10450 4720 10480 4760
rect 10380 4660 10480 4720
rect 10380 4620 10410 4660
rect 10450 4620 10480 4660
rect 10380 4590 10480 4620
rect 10510 4760 10610 4790
rect 10510 4720 10540 4760
rect 10580 4720 10610 4760
rect 10510 4660 10610 4720
rect 10510 4620 10540 4660
rect 10580 4620 10610 4660
rect 10510 4590 10610 4620
rect 3970 4540 3990 4580
rect 4030 4540 4050 4580
rect 3970 4510 4050 4540
rect 7520 4110 7620 4140
rect 7520 4070 7550 4110
rect 7590 4070 7620 4110
rect 7520 4010 7620 4070
rect 7520 3970 7550 4010
rect 7590 3970 7620 4010
rect 7520 3910 7620 3970
rect 7520 3870 7550 3910
rect 7590 3870 7620 3910
rect 7520 3810 7620 3870
rect 7520 3770 7550 3810
rect 7590 3770 7620 3810
rect 7520 3710 7620 3770
rect 7520 3670 7550 3710
rect 7590 3670 7620 3710
rect 7520 3640 7620 3670
rect 7720 4110 7820 4140
rect 7720 4070 7750 4110
rect 7790 4070 7820 4110
rect 7720 4010 7820 4070
rect 7720 3970 7750 4010
rect 7790 3970 7820 4010
rect 7720 3910 7820 3970
rect 7720 3870 7750 3910
rect 7790 3870 7820 3910
rect 7720 3810 7820 3870
rect 7720 3770 7750 3810
rect 7790 3770 7820 3810
rect 7720 3710 7820 3770
rect 7720 3670 7750 3710
rect 7790 3670 7820 3710
rect 7720 3640 7820 3670
rect 7920 4110 8020 4140
rect 7920 4070 7950 4110
rect 7990 4070 8020 4110
rect 7920 4010 8020 4070
rect 7920 3970 7950 4010
rect 7990 3970 8020 4010
rect 7920 3910 8020 3970
rect 7920 3870 7950 3910
rect 7990 3870 8020 3910
rect 7920 3810 8020 3870
rect 7920 3770 7950 3810
rect 7990 3770 8020 3810
rect 7920 3710 8020 3770
rect 7920 3670 7950 3710
rect 7990 3670 8020 3710
rect 7920 3640 8020 3670
rect 8120 4110 8220 4140
rect 8120 4070 8150 4110
rect 8190 4070 8220 4110
rect 8120 4010 8220 4070
rect 8120 3970 8150 4010
rect 8190 3970 8220 4010
rect 8120 3910 8220 3970
rect 8120 3870 8150 3910
rect 8190 3870 8220 3910
rect 8120 3810 8220 3870
rect 8120 3770 8150 3810
rect 8190 3770 8220 3810
rect 8120 3710 8220 3770
rect 8120 3670 8150 3710
rect 8190 3670 8220 3710
rect 8120 3640 8220 3670
rect 8320 4110 8420 4140
rect 8320 4070 8350 4110
rect 8390 4070 8420 4110
rect 8320 4010 8420 4070
rect 8320 3970 8350 4010
rect 8390 3970 8420 4010
rect 8320 3910 8420 3970
rect 8320 3870 8350 3910
rect 8390 3870 8420 3910
rect 8320 3810 8420 3870
rect 8320 3770 8350 3810
rect 8390 3770 8420 3810
rect 8320 3710 8420 3770
rect 8320 3670 8350 3710
rect 8390 3670 8420 3710
rect 8320 3640 8420 3670
rect 8520 4110 8620 4140
rect 8520 4070 8550 4110
rect 8590 4070 8620 4110
rect 8520 4010 8620 4070
rect 8520 3970 8550 4010
rect 8590 3970 8620 4010
rect 8520 3910 8620 3970
rect 8520 3870 8550 3910
rect 8590 3870 8620 3910
rect 8520 3810 8620 3870
rect 8520 3770 8550 3810
rect 8590 3770 8620 3810
rect 8520 3710 8620 3770
rect 8520 3670 8550 3710
rect 8590 3670 8620 3710
rect 8520 3640 8620 3670
rect 8720 4110 8820 4140
rect 8720 4070 8750 4110
rect 8790 4070 8820 4110
rect 8720 4010 8820 4070
rect 8720 3970 8750 4010
rect 8790 3970 8820 4010
rect 8720 3910 8820 3970
rect 8720 3870 8750 3910
rect 8790 3870 8820 3910
rect 8720 3810 8820 3870
rect 8720 3770 8750 3810
rect 8790 3770 8820 3810
rect 8720 3710 8820 3770
rect 8720 3670 8750 3710
rect 8790 3670 8820 3710
rect 8720 3640 8820 3670
rect 8920 4110 9020 4140
rect 8920 4070 8950 4110
rect 8990 4070 9020 4110
rect 8920 4010 9020 4070
rect 8920 3970 8950 4010
rect 8990 3970 9020 4010
rect 8920 3910 9020 3970
rect 8920 3870 8950 3910
rect 8990 3870 9020 3910
rect 8920 3810 9020 3870
rect 8920 3770 8950 3810
rect 8990 3770 9020 3810
rect 8920 3710 9020 3770
rect 8920 3670 8950 3710
rect 8990 3670 9020 3710
rect 8920 3640 9020 3670
rect 9120 4110 9220 4140
rect 9120 4070 9150 4110
rect 9190 4070 9220 4110
rect 9120 4010 9220 4070
rect 9120 3970 9150 4010
rect 9190 3970 9220 4010
rect 9120 3910 9220 3970
rect 9120 3870 9150 3910
rect 9190 3870 9220 3910
rect 9120 3810 9220 3870
rect 9120 3770 9150 3810
rect 9190 3770 9220 3810
rect 9120 3710 9220 3770
rect 9120 3670 9150 3710
rect 9190 3670 9220 3710
rect 9120 3640 9220 3670
rect 9320 4110 9420 4140
rect 9320 4070 9350 4110
rect 9390 4070 9420 4110
rect 9320 4010 9420 4070
rect 9320 3970 9350 4010
rect 9390 3970 9420 4010
rect 9320 3910 9420 3970
rect 9320 3870 9350 3910
rect 9390 3870 9420 3910
rect 9320 3810 9420 3870
rect 9320 3770 9350 3810
rect 9390 3770 9420 3810
rect 9320 3710 9420 3770
rect 9320 3670 9350 3710
rect 9390 3670 9420 3710
rect 9320 3640 9420 3670
rect 9520 4110 9620 4140
rect 9520 4070 9550 4110
rect 9590 4070 9620 4110
rect 9520 4010 9620 4070
rect 9520 3970 9550 4010
rect 9590 3970 9620 4010
rect 9520 3910 9620 3970
rect 9520 3870 9550 3910
rect 9590 3870 9620 3910
rect 9520 3810 9620 3870
rect 9520 3770 9550 3810
rect 9590 3770 9620 3810
rect 9520 3710 9620 3770
rect 9520 3670 9550 3710
rect 9590 3670 9620 3710
rect 9520 3640 9620 3670
rect -410 1198 270 1250
rect -410 1164 -358 1198
rect -324 1164 -268 1198
rect -234 1164 -178 1198
rect -144 1164 -88 1198
rect -54 1164 2 1198
rect 36 1164 92 1198
rect 126 1164 182 1198
rect 216 1164 270 1198
rect -410 1108 270 1164
rect -410 1074 -358 1108
rect -324 1074 -268 1108
rect -234 1074 -178 1108
rect -144 1074 -88 1108
rect -54 1074 2 1108
rect 36 1074 92 1108
rect 126 1074 182 1108
rect 216 1074 270 1108
rect -410 1018 270 1074
rect -410 984 -358 1018
rect -324 984 -268 1018
rect -234 984 -178 1018
rect -144 984 -88 1018
rect -54 984 2 1018
rect 36 984 92 1018
rect 126 984 182 1018
rect 216 984 270 1018
rect -410 928 270 984
rect -410 894 -358 928
rect -324 894 -268 928
rect -234 894 -178 928
rect -144 894 -88 928
rect -54 894 2 928
rect 36 894 92 928
rect 126 894 182 928
rect 216 894 270 928
rect -410 838 270 894
rect -410 804 -358 838
rect -324 804 -268 838
rect -234 804 -178 838
rect -144 804 -88 838
rect -54 804 2 838
rect 36 804 92 838
rect 126 804 182 838
rect 216 804 270 838
rect -410 748 270 804
rect -410 714 -358 748
rect -324 714 -268 748
rect -234 714 -178 748
rect -144 714 -88 748
rect -54 714 2 748
rect 36 714 92 748
rect 126 714 182 748
rect 216 714 270 748
rect -410 658 270 714
rect -410 624 -358 658
rect -324 624 -268 658
rect -234 624 -178 658
rect -144 624 -88 658
rect -54 624 2 658
rect 36 624 92 658
rect 126 624 182 658
rect 216 624 270 658
rect -410 570 270 624
rect 950 1198 1630 1250
rect 950 1164 1002 1198
rect 1036 1164 1092 1198
rect 1126 1164 1182 1198
rect 1216 1164 1272 1198
rect 1306 1164 1362 1198
rect 1396 1164 1452 1198
rect 1486 1164 1542 1198
rect 1576 1164 1630 1198
rect 950 1108 1630 1164
rect 950 1074 1002 1108
rect 1036 1074 1092 1108
rect 1126 1074 1182 1108
rect 1216 1074 1272 1108
rect 1306 1074 1362 1108
rect 1396 1074 1452 1108
rect 1486 1074 1542 1108
rect 1576 1074 1630 1108
rect 950 1018 1630 1074
rect 950 984 1002 1018
rect 1036 984 1092 1018
rect 1126 984 1182 1018
rect 1216 984 1272 1018
rect 1306 984 1362 1018
rect 1396 984 1452 1018
rect 1486 984 1542 1018
rect 1576 984 1630 1018
rect 950 928 1630 984
rect 950 894 1002 928
rect 1036 894 1092 928
rect 1126 894 1182 928
rect 1216 894 1272 928
rect 1306 894 1362 928
rect 1396 894 1452 928
rect 1486 894 1542 928
rect 1576 894 1630 928
rect 950 838 1630 894
rect 950 804 1002 838
rect 1036 804 1092 838
rect 1126 804 1182 838
rect 1216 804 1272 838
rect 1306 804 1362 838
rect 1396 804 1452 838
rect 1486 804 1542 838
rect 1576 804 1630 838
rect 950 748 1630 804
rect 950 714 1002 748
rect 1036 714 1092 748
rect 1126 714 1182 748
rect 1216 714 1272 748
rect 1306 714 1362 748
rect 1396 714 1452 748
rect 1486 714 1542 748
rect 1576 714 1630 748
rect 950 658 1630 714
rect 950 624 1002 658
rect 1036 624 1092 658
rect 1126 624 1182 658
rect 1216 624 1272 658
rect 1306 624 1362 658
rect 1396 624 1452 658
rect 1486 624 1542 658
rect 1576 624 1630 658
rect 950 570 1630 624
rect 2310 1198 2990 1250
rect 2310 1164 2362 1198
rect 2396 1164 2452 1198
rect 2486 1164 2542 1198
rect 2576 1164 2632 1198
rect 2666 1164 2722 1198
rect 2756 1164 2812 1198
rect 2846 1164 2902 1198
rect 2936 1164 2990 1198
rect 2310 1108 2990 1164
rect 2310 1074 2362 1108
rect 2396 1074 2452 1108
rect 2486 1074 2542 1108
rect 2576 1074 2632 1108
rect 2666 1074 2722 1108
rect 2756 1074 2812 1108
rect 2846 1074 2902 1108
rect 2936 1074 2990 1108
rect 2310 1018 2990 1074
rect 2310 984 2362 1018
rect 2396 984 2452 1018
rect 2486 984 2542 1018
rect 2576 984 2632 1018
rect 2666 984 2722 1018
rect 2756 984 2812 1018
rect 2846 984 2902 1018
rect 2936 984 2990 1018
rect 2310 928 2990 984
rect 2310 894 2362 928
rect 2396 894 2452 928
rect 2486 894 2542 928
rect 2576 894 2632 928
rect 2666 894 2722 928
rect 2756 894 2812 928
rect 2846 894 2902 928
rect 2936 894 2990 928
rect 2310 838 2990 894
rect 2310 804 2362 838
rect 2396 804 2452 838
rect 2486 804 2542 838
rect 2576 804 2632 838
rect 2666 804 2722 838
rect 2756 804 2812 838
rect 2846 804 2902 838
rect 2936 804 2990 838
rect 2310 748 2990 804
rect 2310 714 2362 748
rect 2396 714 2452 748
rect 2486 714 2542 748
rect 2576 714 2632 748
rect 2666 714 2722 748
rect 2756 714 2812 748
rect 2846 714 2902 748
rect 2936 714 2990 748
rect 2310 658 2990 714
rect 2310 624 2362 658
rect 2396 624 2452 658
rect 2486 624 2542 658
rect 2576 624 2632 658
rect 2666 624 2722 658
rect 2756 624 2812 658
rect 2846 624 2902 658
rect 2936 624 2990 658
rect 2310 570 2990 624
rect -410 -162 270 -110
rect -410 -196 -358 -162
rect -324 -196 -268 -162
rect -234 -196 -178 -162
rect -144 -196 -88 -162
rect -54 -196 2 -162
rect 36 -196 92 -162
rect 126 -196 182 -162
rect 216 -196 270 -162
rect -410 -252 270 -196
rect -410 -286 -358 -252
rect -324 -286 -268 -252
rect -234 -286 -178 -252
rect -144 -286 -88 -252
rect -54 -286 2 -252
rect 36 -286 92 -252
rect 126 -286 182 -252
rect 216 -286 270 -252
rect -410 -342 270 -286
rect -410 -376 -358 -342
rect -324 -376 -268 -342
rect -234 -376 -178 -342
rect -144 -376 -88 -342
rect -54 -376 2 -342
rect 36 -376 92 -342
rect 126 -376 182 -342
rect 216 -376 270 -342
rect -410 -432 270 -376
rect -410 -466 -358 -432
rect -324 -466 -268 -432
rect -234 -466 -178 -432
rect -144 -466 -88 -432
rect -54 -466 2 -432
rect 36 -466 92 -432
rect 126 -466 182 -432
rect 216 -466 270 -432
rect -410 -522 270 -466
rect -410 -556 -358 -522
rect -324 -556 -268 -522
rect -234 -556 -178 -522
rect -144 -556 -88 -522
rect -54 -556 2 -522
rect 36 -556 92 -522
rect 126 -556 182 -522
rect 216 -556 270 -522
rect -410 -612 270 -556
rect -410 -646 -358 -612
rect -324 -646 -268 -612
rect -234 -646 -178 -612
rect -144 -646 -88 -612
rect -54 -646 2 -612
rect 36 -646 92 -612
rect 126 -646 182 -612
rect 216 -646 270 -612
rect -410 -702 270 -646
rect -410 -736 -358 -702
rect -324 -736 -268 -702
rect -234 -736 -178 -702
rect -144 -736 -88 -702
rect -54 -736 2 -702
rect 36 -736 92 -702
rect 126 -736 182 -702
rect 216 -736 270 -702
rect -410 -790 270 -736
rect 950 -162 1630 -110
rect 950 -196 1002 -162
rect 1036 -196 1092 -162
rect 1126 -196 1182 -162
rect 1216 -196 1272 -162
rect 1306 -196 1362 -162
rect 1396 -196 1452 -162
rect 1486 -196 1542 -162
rect 1576 -196 1630 -162
rect 950 -252 1630 -196
rect 950 -286 1002 -252
rect 1036 -286 1092 -252
rect 1126 -286 1182 -252
rect 1216 -286 1272 -252
rect 1306 -286 1362 -252
rect 1396 -286 1452 -252
rect 1486 -286 1542 -252
rect 1576 -286 1630 -252
rect 950 -342 1630 -286
rect 950 -376 1002 -342
rect 1036 -376 1092 -342
rect 1126 -376 1182 -342
rect 1216 -376 1272 -342
rect 1306 -376 1362 -342
rect 1396 -376 1452 -342
rect 1486 -376 1542 -342
rect 1576 -376 1630 -342
rect 950 -432 1630 -376
rect 950 -466 1002 -432
rect 1036 -466 1092 -432
rect 1126 -466 1182 -432
rect 1216 -466 1272 -432
rect 1306 -466 1362 -432
rect 1396 -466 1452 -432
rect 1486 -466 1542 -432
rect 1576 -466 1630 -432
rect 950 -522 1630 -466
rect 950 -556 1002 -522
rect 1036 -556 1092 -522
rect 1126 -556 1182 -522
rect 1216 -556 1272 -522
rect 1306 -556 1362 -522
rect 1396 -556 1452 -522
rect 1486 -556 1542 -522
rect 1576 -556 1630 -522
rect 950 -612 1630 -556
rect 950 -646 1002 -612
rect 1036 -646 1092 -612
rect 1126 -646 1182 -612
rect 1216 -646 1272 -612
rect 1306 -646 1362 -612
rect 1396 -646 1452 -612
rect 1486 -646 1542 -612
rect 1576 -646 1630 -612
rect 950 -702 1630 -646
rect 950 -736 1002 -702
rect 1036 -736 1092 -702
rect 1126 -736 1182 -702
rect 1216 -736 1272 -702
rect 1306 -736 1362 -702
rect 1396 -736 1452 -702
rect 1486 -736 1542 -702
rect 1576 -736 1630 -702
rect 950 -790 1630 -736
rect 2310 -162 2990 -110
rect 2310 -196 2362 -162
rect 2396 -196 2452 -162
rect 2486 -196 2542 -162
rect 2576 -196 2632 -162
rect 2666 -196 2722 -162
rect 2756 -196 2812 -162
rect 2846 -196 2902 -162
rect 2936 -196 2990 -162
rect 2310 -252 2990 -196
rect 2310 -286 2362 -252
rect 2396 -286 2452 -252
rect 2486 -286 2542 -252
rect 2576 -286 2632 -252
rect 2666 -286 2722 -252
rect 2756 -286 2812 -252
rect 2846 -286 2902 -252
rect 2936 -286 2990 -252
rect 2310 -342 2990 -286
rect 2310 -376 2362 -342
rect 2396 -376 2452 -342
rect 2486 -376 2542 -342
rect 2576 -376 2632 -342
rect 2666 -376 2722 -342
rect 2756 -376 2812 -342
rect 2846 -376 2902 -342
rect 2936 -376 2990 -342
rect 2310 -432 2990 -376
rect 2310 -466 2362 -432
rect 2396 -466 2452 -432
rect 2486 -466 2542 -432
rect 2576 -466 2632 -432
rect 2666 -466 2722 -432
rect 2756 -466 2812 -432
rect 2846 -466 2902 -432
rect 2936 -466 2990 -432
rect 2310 -522 2990 -466
rect 2310 -556 2362 -522
rect 2396 -556 2452 -522
rect 2486 -556 2542 -522
rect 2576 -556 2632 -522
rect 2666 -556 2722 -522
rect 2756 -556 2812 -522
rect 2846 -556 2902 -522
rect 2936 -556 2990 -522
rect 2310 -612 2990 -556
rect 2310 -646 2362 -612
rect 2396 -646 2452 -612
rect 2486 -646 2542 -612
rect 2576 -646 2632 -612
rect 2666 -646 2722 -612
rect 2756 -646 2812 -612
rect 2846 -646 2902 -612
rect 2936 -646 2990 -612
rect 2310 -702 2990 -646
rect 2310 -736 2362 -702
rect 2396 -736 2452 -702
rect 2486 -736 2542 -702
rect 2576 -736 2632 -702
rect 2666 -736 2722 -702
rect 2756 -736 2812 -702
rect 2846 -736 2902 -702
rect 2936 -736 2990 -702
rect 2310 -790 2990 -736
rect -410 -1522 270 -1470
rect -410 -1556 -358 -1522
rect -324 -1556 -268 -1522
rect -234 -1556 -178 -1522
rect -144 -1556 -88 -1522
rect -54 -1556 2 -1522
rect 36 -1556 92 -1522
rect 126 -1556 182 -1522
rect 216 -1556 270 -1522
rect -410 -1612 270 -1556
rect -410 -1646 -358 -1612
rect -324 -1646 -268 -1612
rect -234 -1646 -178 -1612
rect -144 -1646 -88 -1612
rect -54 -1646 2 -1612
rect 36 -1646 92 -1612
rect 126 -1646 182 -1612
rect 216 -1646 270 -1612
rect -410 -1702 270 -1646
rect -410 -1736 -358 -1702
rect -324 -1736 -268 -1702
rect -234 -1736 -178 -1702
rect -144 -1736 -88 -1702
rect -54 -1736 2 -1702
rect 36 -1736 92 -1702
rect 126 -1736 182 -1702
rect 216 -1736 270 -1702
rect -410 -1792 270 -1736
rect -410 -1826 -358 -1792
rect -324 -1826 -268 -1792
rect -234 -1826 -178 -1792
rect -144 -1826 -88 -1792
rect -54 -1826 2 -1792
rect 36 -1826 92 -1792
rect 126 -1826 182 -1792
rect 216 -1826 270 -1792
rect -410 -1882 270 -1826
rect -410 -1916 -358 -1882
rect -324 -1916 -268 -1882
rect -234 -1916 -178 -1882
rect -144 -1916 -88 -1882
rect -54 -1916 2 -1882
rect 36 -1916 92 -1882
rect 126 -1916 182 -1882
rect 216 -1916 270 -1882
rect -410 -1972 270 -1916
rect -410 -2006 -358 -1972
rect -324 -2006 -268 -1972
rect -234 -2006 -178 -1972
rect -144 -2006 -88 -1972
rect -54 -2006 2 -1972
rect 36 -2006 92 -1972
rect 126 -2006 182 -1972
rect 216 -2006 270 -1972
rect -410 -2062 270 -2006
rect -410 -2096 -358 -2062
rect -324 -2096 -268 -2062
rect -234 -2096 -178 -2062
rect -144 -2096 -88 -2062
rect -54 -2096 2 -2062
rect 36 -2096 92 -2062
rect 126 -2096 182 -2062
rect 216 -2096 270 -2062
rect -410 -2150 270 -2096
rect 950 -1522 1630 -1470
rect 950 -1556 1002 -1522
rect 1036 -1556 1092 -1522
rect 1126 -1556 1182 -1522
rect 1216 -1556 1272 -1522
rect 1306 -1556 1362 -1522
rect 1396 -1556 1452 -1522
rect 1486 -1556 1542 -1522
rect 1576 -1556 1630 -1522
rect 950 -1612 1630 -1556
rect 950 -1646 1002 -1612
rect 1036 -1646 1092 -1612
rect 1126 -1646 1182 -1612
rect 1216 -1646 1272 -1612
rect 1306 -1646 1362 -1612
rect 1396 -1646 1452 -1612
rect 1486 -1646 1542 -1612
rect 1576 -1646 1630 -1612
rect 950 -1702 1630 -1646
rect 950 -1736 1002 -1702
rect 1036 -1736 1092 -1702
rect 1126 -1736 1182 -1702
rect 1216 -1736 1272 -1702
rect 1306 -1736 1362 -1702
rect 1396 -1736 1452 -1702
rect 1486 -1736 1542 -1702
rect 1576 -1736 1630 -1702
rect 950 -1792 1630 -1736
rect 950 -1826 1002 -1792
rect 1036 -1826 1092 -1792
rect 1126 -1826 1182 -1792
rect 1216 -1826 1272 -1792
rect 1306 -1826 1362 -1792
rect 1396 -1826 1452 -1792
rect 1486 -1826 1542 -1792
rect 1576 -1826 1630 -1792
rect 950 -1882 1630 -1826
rect 950 -1916 1002 -1882
rect 1036 -1916 1092 -1882
rect 1126 -1916 1182 -1882
rect 1216 -1916 1272 -1882
rect 1306 -1916 1362 -1882
rect 1396 -1916 1452 -1882
rect 1486 -1916 1542 -1882
rect 1576 -1916 1630 -1882
rect 950 -1972 1630 -1916
rect 950 -2006 1002 -1972
rect 1036 -2006 1092 -1972
rect 1126 -2006 1182 -1972
rect 1216 -2006 1272 -1972
rect 1306 -2006 1362 -1972
rect 1396 -2006 1452 -1972
rect 1486 -2006 1542 -1972
rect 1576 -2006 1630 -1972
rect 950 -2062 1630 -2006
rect 950 -2096 1002 -2062
rect 1036 -2096 1092 -2062
rect 1126 -2096 1182 -2062
rect 1216 -2096 1272 -2062
rect 1306 -2096 1362 -2062
rect 1396 -2096 1452 -2062
rect 1486 -2096 1542 -2062
rect 1576 -2096 1630 -2062
rect 950 -2150 1630 -2096
rect 2310 -1522 2990 -1470
rect 2310 -1556 2362 -1522
rect 2396 -1556 2452 -1522
rect 2486 -1556 2542 -1522
rect 2576 -1556 2632 -1522
rect 2666 -1556 2722 -1522
rect 2756 -1556 2812 -1522
rect 2846 -1556 2902 -1522
rect 2936 -1556 2990 -1522
rect 2310 -1612 2990 -1556
rect 2310 -1646 2362 -1612
rect 2396 -1646 2452 -1612
rect 2486 -1646 2542 -1612
rect 2576 -1646 2632 -1612
rect 2666 -1646 2722 -1612
rect 2756 -1646 2812 -1612
rect 2846 -1646 2902 -1612
rect 2936 -1646 2990 -1612
rect 2310 -1702 2990 -1646
rect 2310 -1736 2362 -1702
rect 2396 -1736 2452 -1702
rect 2486 -1736 2542 -1702
rect 2576 -1736 2632 -1702
rect 2666 -1736 2722 -1702
rect 2756 -1736 2812 -1702
rect 2846 -1736 2902 -1702
rect 2936 -1736 2990 -1702
rect 2310 -1792 2990 -1736
rect 2310 -1826 2362 -1792
rect 2396 -1826 2452 -1792
rect 2486 -1826 2542 -1792
rect 2576 -1826 2632 -1792
rect 2666 -1826 2722 -1792
rect 2756 -1826 2812 -1792
rect 2846 -1826 2902 -1792
rect 2936 -1826 2990 -1792
rect 2310 -1882 2990 -1826
rect 2310 -1916 2362 -1882
rect 2396 -1916 2452 -1882
rect 2486 -1916 2542 -1882
rect 2576 -1916 2632 -1882
rect 2666 -1916 2722 -1882
rect 2756 -1916 2812 -1882
rect 2846 -1916 2902 -1882
rect 2936 -1916 2990 -1882
rect 2310 -1972 2990 -1916
rect 2310 -2006 2362 -1972
rect 2396 -2006 2452 -1972
rect 2486 -2006 2542 -1972
rect 2576 -2006 2632 -1972
rect 2666 -2006 2722 -1972
rect 2756 -2006 2812 -1972
rect 2846 -2006 2902 -1972
rect 2936 -2006 2990 -1972
rect 2310 -2062 2990 -2006
rect 2310 -2096 2362 -2062
rect 2396 -2096 2452 -2062
rect 2486 -2096 2542 -2062
rect 2576 -2096 2632 -2062
rect 2666 -2096 2722 -2062
rect 2756 -2096 2812 -2062
rect 2846 -2096 2902 -2062
rect 2936 -2096 2990 -2062
rect 2310 -2150 2990 -2096
<< ndiffc >>
rect 11230 14280 11270 14320
rect 11230 14180 11270 14220
rect 11340 14280 11380 14320
rect 11340 14180 11380 14220
rect 11750 14280 11790 14320
rect 11750 14180 11790 14220
rect 11860 14280 11900 14320
rect 11860 14180 11900 14220
rect 12270 14280 12310 14320
rect 12270 14180 12310 14220
rect 12380 14280 12420 14320
rect 12380 14180 12420 14220
rect 12870 14280 12910 14320
rect 12870 14180 12910 14220
rect 12980 14280 13020 14320
rect 12980 14180 13020 14220
rect 11230 13900 11270 13940
rect 11230 13800 11270 13840
rect 11230 13700 11270 13740
rect 11340 13900 11380 13940
rect 11340 13800 11380 13840
rect 11340 13700 11380 13740
rect 11750 13900 11790 13940
rect 11750 13800 11790 13840
rect 11750 13700 11790 13740
rect 11860 13900 11900 13940
rect 11860 13800 11900 13840
rect 11860 13700 11900 13740
rect 12270 13900 12310 13940
rect 12270 13800 12310 13840
rect 12270 13700 12310 13740
rect 12380 13900 12420 13940
rect 12380 13800 12420 13840
rect 12380 13700 12420 13740
rect 460 13150 500 13190
rect 570 13150 610 13190
rect 680 13150 720 13190
rect 790 13150 830 13190
rect 900 13150 940 13190
rect 1040 13150 1080 13190
rect 1150 13150 1190 13190
rect 1260 13150 1300 13190
rect 1490 13150 1530 13190
rect 1600 13150 1640 13190
rect 1710 13150 1750 13190
rect 1820 13150 1860 13190
rect 1930 13150 1970 13190
rect 2150 13150 2190 13190
rect 2260 13150 2300 13190
rect 2370 13150 2410 13190
rect 2480 13150 2520 13190
rect 2590 13150 2630 13190
rect 2830 13150 2870 13190
rect 2940 13150 2980 13190
rect 3050 13150 3090 13190
rect 3160 13150 3200 13190
rect 3270 13150 3310 13190
rect 3410 13150 3450 13190
rect 3520 13150 3560 13190
rect 3630 13150 3670 13190
rect 3970 13150 4010 13190
rect 4080 13150 4120 13190
rect 4330 13150 4370 13190
rect 4440 13150 4480 13190
rect 4580 13150 4620 13190
rect 4690 13150 4730 13190
rect 4800 13150 4840 13190
rect 4910 13150 4950 13190
rect 5020 13150 5060 13190
rect 5240 13150 5280 13190
rect 5350 13150 5390 13190
rect 5460 13150 5500 13190
rect 5570 13150 5610 13190
rect 5790 13150 5830 13190
rect 5900 13150 5940 13190
rect 6010 13150 6050 13190
rect 6120 13150 6160 13190
rect 6230 13150 6270 13190
rect 6450 13150 6490 13190
rect 6560 13150 6600 13190
rect 6670 13150 6710 13190
rect 7090 13240 7130 13280
rect 7200 13240 7240 13280
rect 7310 13240 7350 13280
rect 7420 13240 7460 13280
rect 7530 13240 7570 13280
rect 7750 13240 7790 13280
rect 7860 13240 7900 13280
rect 7970 13240 8010 13280
rect 8080 13240 8120 13280
rect 8390 13240 8430 13280
rect 8500 13240 8540 13280
rect 8610 13240 8650 13280
rect 8720 13240 8760 13280
rect 8830 13240 8870 13280
rect 9050 13240 9090 13280
rect 9160 13240 9200 13280
rect 9270 13240 9310 13280
rect 9380 13240 9420 13280
rect 9690 13240 9730 13280
rect 9800 13240 9840 13280
rect 9910 13240 9950 13280
rect 10020 13240 10060 13280
rect 10130 13240 10170 13280
rect 10350 13240 10390 13280
rect 10460 13240 10500 13280
rect 10570 13240 10610 13280
rect 10680 13240 10720 13280
rect 6780 13150 6820 13190
rect 11228 13420 11268 13460
rect 11228 13320 11268 13360
rect 11340 13420 11380 13460
rect 11340 13320 11380 13360
rect 11748 13420 11788 13460
rect 11748 13320 11788 13360
rect 11860 13420 11900 13460
rect 11860 13320 11900 13360
rect 12268 13420 12308 13460
rect 12268 13320 12308 13360
rect 12380 13420 12420 13460
rect 12380 13320 12420 13360
rect 1280 10170 1320 10210
rect 1280 10070 1320 10110
rect 1390 10170 1430 10210
rect 1390 10070 1430 10110
rect 1500 10170 1540 10210
rect 1500 10070 1540 10110
rect 1800 10170 1840 10210
rect 1800 10070 1840 10110
rect 1910 10170 1950 10210
rect 1910 10070 1950 10110
rect 2020 10170 2060 10210
rect 2180 10170 2220 10210
rect 2020 10070 2060 10110
rect 2180 10070 2220 10110
rect 2290 10170 2330 10210
rect 2290 10070 2330 10110
rect 2400 10170 2440 10210
rect 2400 10070 2440 10110
rect 2700 10170 2740 10210
rect 2700 10070 2740 10110
rect 2810 10170 2850 10210
rect 2810 10070 2850 10110
rect 2920 10170 2960 10210
rect 2920 10070 2960 10110
rect 3220 10170 3260 10210
rect 3220 10070 3260 10110
rect 3330 10170 3370 10210
rect 3330 10070 3370 10110
rect 3440 10170 3480 10210
rect 3440 10070 3480 10110
rect 3660 10170 3700 10210
rect 3660 10070 3700 10110
rect 3770 10170 3810 10210
rect 3770 10070 3810 10110
rect 3990 10170 4030 10210
rect 3990 10070 4030 10110
rect 4100 10170 4140 10210
rect 4100 10070 4140 10110
rect 4420 10170 4460 10210
rect 4420 10070 4460 10110
rect 4550 10170 4590 10210
rect 4550 10070 4590 10110
rect 4810 10170 4850 10210
rect 4810 10070 4850 10110
rect 4940 10170 4980 10210
rect 4940 10070 4980 10110
rect 5200 10170 5240 10210
rect 5200 10070 5240 10110
rect 5330 10170 5370 10210
rect 5330 10070 5370 10110
rect 5490 10170 5530 10210
rect 5490 10070 5530 10110
rect 5620 10170 5660 10210
rect 5620 10070 5660 10110
rect 7370 8620 7410 8660
rect 7370 8520 7410 8560
rect 1280 8370 1320 8410
rect 1280 8270 1320 8310
rect 1390 8370 1430 8410
rect 1390 8270 1430 8310
rect 1500 8370 1540 8410
rect 1500 8270 1540 8310
rect 1800 8370 1840 8410
rect 1800 8270 1840 8310
rect 1910 8370 1950 8410
rect 1910 8270 1950 8310
rect 2020 8370 2060 8410
rect 2180 8370 2220 8410
rect 2020 8270 2060 8310
rect 2180 8270 2220 8310
rect 2290 8370 2330 8410
rect 2290 8270 2330 8310
rect 2400 8370 2440 8410
rect 2400 8270 2440 8310
rect 2700 8370 2740 8410
rect 2700 8270 2740 8310
rect 2810 8370 2850 8410
rect 2810 8270 2850 8310
rect 2920 8370 2960 8410
rect 2920 8270 2960 8310
rect 3210 8370 3250 8410
rect 3210 8270 3250 8310
rect 3320 8370 3360 8410
rect 3320 8270 3360 8310
rect 3540 8370 3580 8410
rect 3540 8270 3580 8310
rect 3650 8370 3690 8410
rect 3650 8270 3690 8310
rect 3870 8370 3910 8410
rect 3870 8270 3910 8310
rect 3980 8370 4020 8410
rect 3980 8270 4020 8310
rect 4420 8370 4460 8410
rect 4420 8270 4460 8310
rect 4550 8370 4590 8410
rect 4550 8270 4590 8310
rect 4810 8370 4850 8410
rect 4810 8270 4850 8310
rect 4940 8370 4980 8410
rect 4940 8270 4980 8310
rect 5200 8370 5240 8410
rect 5200 8270 5240 8310
rect 5330 8370 5370 8410
rect 5330 8270 5370 8310
rect 5490 8370 5530 8410
rect 5490 8270 5530 8310
rect 5620 8370 5660 8410
rect 5620 8270 5660 8310
rect 5880 8370 5920 8410
rect 5880 8270 5920 8310
rect 6010 8370 6050 8410
rect 6010 8270 6050 8310
rect 7370 8420 7410 8460
rect 7370 8320 7410 8360
rect 7590 8620 7630 8660
rect 7590 8520 7630 8560
rect 7590 8420 7630 8460
rect 7590 8320 7630 8360
rect 7810 8620 7850 8660
rect 7810 8520 7850 8560
rect 7810 8420 7850 8460
rect 7810 8320 7850 8360
rect 8030 8620 8070 8660
rect 8030 8520 8070 8560
rect 8030 8420 8070 8460
rect 8030 8320 8070 8360
rect 8250 8620 8290 8660
rect 8450 8620 8490 8660
rect 8250 8520 8290 8560
rect 8450 8520 8490 8560
rect 8250 8420 8290 8460
rect 8450 8420 8490 8460
rect 8250 8320 8290 8360
rect 8450 8320 8490 8360
rect 8670 8620 8710 8660
rect 8670 8520 8710 8560
rect 8670 8420 8710 8460
rect 8670 8320 8710 8360
rect 8890 8620 8930 8660
rect 8890 8520 8930 8560
rect 8890 8420 8930 8460
rect 8890 8320 8930 8360
rect 9110 8620 9150 8660
rect 9110 8520 9150 8560
rect 9110 8420 9150 8460
rect 9110 8320 9150 8360
rect 9330 8620 9370 8660
rect 9530 8620 9570 8660
rect 9330 8520 9370 8560
rect 9530 8520 9570 8560
rect 9330 8420 9370 8460
rect 9530 8420 9570 8460
rect 9330 8320 9370 8360
rect 9530 8320 9570 8360
rect 9750 8620 9790 8660
rect 9750 8520 9790 8560
rect 9750 8420 9790 8460
rect 9750 8320 9790 8360
rect 9970 8620 10010 8660
rect 9970 8520 10010 8560
rect 9970 8420 10010 8460
rect 9970 8320 10010 8360
rect 10190 8620 10230 8660
rect 10190 8520 10230 8560
rect 10190 8420 10230 8460
rect 10190 8320 10230 8360
rect 10410 8620 10450 8660
rect 10410 8520 10450 8560
rect 10410 8420 10450 8460
rect 10410 8320 10450 8360
rect 7430 5980 7470 6030
rect 7430 5840 7470 5890
rect 7630 5980 7670 6030
rect 7630 5840 7670 5890
rect 7830 5980 7870 6030
rect 7830 5840 7870 5890
rect 8030 5980 8070 6030
rect 8030 5840 8070 5890
rect 8230 5980 8270 6030
rect 8230 5840 8270 5890
rect 8430 5980 8470 6030
rect 8430 5840 8470 5890
rect 8630 5980 8670 6030
rect 8630 5840 8670 5890
rect 8830 5980 8870 6030
rect 8830 5840 8870 5890
rect 9030 5980 9070 6030
rect 9030 5840 9070 5890
rect 9230 5980 9270 6030
rect 9230 5840 9270 5890
rect 9430 5980 9470 6030
rect 9430 5840 9470 5890
rect 7480 5300 7520 5340
rect 7610 5300 7650 5340
rect 7740 5300 7780 5340
rect 7870 5300 7910 5340
rect 8000 5300 8040 5340
rect 8130 5300 8170 5340
rect 8260 5300 8300 5340
rect 8620 5300 8660 5340
rect 8750 5300 8790 5340
rect 8880 5300 8920 5340
rect 9010 5300 9050 5340
rect 9140 5300 9180 5340
rect 9270 5300 9310 5340
rect 9400 5300 9440 5340
rect 9760 5300 9800 5340
rect 9890 5300 9930 5340
rect 10020 5300 10060 5340
rect 10150 5300 10190 5340
rect 10280 5300 10320 5340
rect 10410 5300 10450 5340
rect 10540 5300 10580 5340
rect -610 3700 -570 3740
rect -490 3700 -450 3740
rect -370 3700 -330 3740
rect -250 3700 -210 3740
rect -130 3700 -90 3740
rect -10 3700 30 3740
rect 110 3700 150 3740
rect 230 3700 270 3740
rect 350 3700 390 3740
rect 470 3700 510 3740
rect 590 3700 630 3740
rect 1950 3700 1990 3740
rect 2070 3700 2110 3740
rect 2190 3700 2230 3740
rect 2310 3700 2350 3740
rect 2430 3700 2470 3740
rect 2550 3700 2590 3740
rect 2670 3700 2710 3740
rect 2790 3700 2830 3740
rect 2910 3700 2950 3740
rect 3030 3700 3070 3740
rect 3150 3700 3190 3740
rect -1230 3090 -1190 3130
rect -1230 2990 -1190 3030
rect -1230 2890 -1190 2930
rect -1230 2790 -1190 2830
rect -1230 2690 -1190 2730
rect -150 3090 -110 3130
rect 10 3090 50 3130
rect -150 2990 -110 3030
rect 10 2990 50 3030
rect -150 2890 -110 2930
rect 10 2890 50 2930
rect -150 2790 -110 2830
rect 10 2790 50 2830
rect -150 2690 -110 2730
rect 10 2690 50 2730
rect 1090 3090 1130 3130
rect 1090 2990 1130 3030
rect 1090 2890 1130 2930
rect 1090 2790 1130 2830
rect 1090 2690 1130 2730
rect 1450 3090 1490 3130
rect 1450 2990 1490 3030
rect 1450 2890 1490 2930
rect 1450 2790 1490 2830
rect 1450 2690 1490 2730
rect 2530 3090 2570 3130
rect 2690 3090 2730 3130
rect 2530 2990 2570 3030
rect 2690 2990 2730 3030
rect 2530 2890 2570 2930
rect 2690 2890 2730 2930
rect 2530 2790 2570 2830
rect 2690 2790 2730 2830
rect 2530 2690 2570 2730
rect 2690 2690 2730 2730
rect 3770 3090 3810 3130
rect 3770 2990 3810 3030
rect 3770 2890 3810 2930
rect 3770 2790 3810 2830
rect 3770 2690 3810 2730
rect -810 2180 -770 2220
rect -810 2080 -770 2120
rect 1270 2180 1310 2220
rect 1270 2080 1310 2120
rect 3350 2180 3390 2220
rect 3350 2080 3390 2120
<< pdiffc >>
rect 620 12830 660 12870
rect 730 12830 770 12870
rect 1040 12830 1080 12870
rect 1150 12830 1190 12870
rect 1260 12830 1300 12870
rect 1710 12830 1750 12870
rect 1820 12830 1860 12870
rect 1930 12830 1970 12870
rect 2150 12830 2190 12870
rect 2260 12830 2300 12870
rect 2370 12830 2410 12870
rect 2480 12830 2520 12870
rect 2990 12830 3030 12870
rect 3100 12830 3140 12870
rect 3410 12830 3450 12870
rect 3520 12830 3560 12870
rect 3630 12830 3670 12870
rect 3860 12830 3900 12870
rect 3970 12830 4010 12870
rect 4080 12830 4120 12870
rect 4220 12830 4260 12870
rect 4330 12830 4370 12870
rect 4440 12830 4480 12870
rect 4800 12830 4840 12870
rect 4910 12830 4950 12870
rect 5020 12830 5060 12870
rect 5240 12830 5280 12870
rect 5350 12830 5390 12870
rect 5460 12830 5500 12870
rect 5860 12830 5900 12870
rect 5970 12830 6010 12870
rect 6200 12830 6240 12870
rect 6310 12830 6350 12870
rect 6420 12830 6460 12870
rect 6560 12830 6600 12870
rect 6670 12830 6710 12870
rect 6780 12830 6820 12870
rect 7160 12830 7200 12870
rect 7270 12830 7310 12870
rect 7500 12830 7540 12870
rect 7610 12830 7650 12870
rect 7720 12830 7760 12870
rect 7860 12830 7900 12870
rect 7970 12830 8010 12870
rect 8080 12830 8120 12870
rect 8460 12830 8500 12870
rect 8570 12830 8610 12870
rect 8800 12830 8840 12870
rect 8910 12830 8950 12870
rect 9020 12830 9060 12870
rect 9160 12830 9200 12870
rect 9270 12830 9310 12870
rect 9380 12830 9420 12870
rect 9760 12830 9800 12870
rect 9870 12830 9910 12870
rect 10100 12830 10140 12870
rect 10210 12830 10250 12870
rect 10320 12830 10360 12870
rect 10460 12830 10500 12870
rect 10570 12830 10610 12870
rect 10680 12830 10720 12870
rect 11228 12700 11268 12740
rect 11228 12600 11268 12640
rect 11228 12500 11268 12540
rect 11228 12400 11268 12440
rect 11340 12700 11380 12740
rect 11340 12600 11380 12640
rect 11340 12500 11380 12540
rect 11340 12400 11380 12440
rect 11748 12700 11788 12740
rect 11748 12600 11788 12640
rect 11748 12500 11788 12540
rect 11748 12400 11788 12440
rect 11860 12700 11900 12740
rect 11860 12600 11900 12640
rect 11860 12500 11900 12540
rect 11860 12400 11900 12440
rect 12268 12700 12308 12740
rect 12268 12600 12308 12640
rect 12268 12500 12308 12540
rect 12268 12400 12308 12440
rect 12380 12700 12420 12740
rect 12380 12600 12420 12640
rect 12380 12500 12420 12540
rect 12380 12400 12420 12440
rect 11230 12120 11270 12160
rect 11230 12020 11270 12060
rect 11230 11920 11270 11960
rect 11230 11820 11270 11860
rect 11230 11720 11270 11760
rect 11230 11620 11270 11660
rect 11340 12120 11380 12160
rect 11340 12020 11380 12060
rect 11340 11920 11380 11960
rect 11340 11820 11380 11860
rect 11340 11720 11380 11760
rect 11340 11620 11380 11660
rect 11750 12120 11790 12160
rect 11750 12020 11790 12060
rect 11750 11920 11790 11960
rect 11750 11820 11790 11860
rect 11750 11720 11790 11760
rect 11750 11620 11790 11660
rect 11860 12120 11900 12160
rect 11860 12020 11900 12060
rect 11860 11920 11900 11960
rect 11860 11820 11900 11860
rect 11860 11720 11900 11760
rect 11860 11620 11900 11660
rect 12270 12120 12310 12160
rect 12270 12020 12310 12060
rect 12270 11920 12310 11960
rect 12270 11820 12310 11860
rect 12270 11720 12310 11760
rect 12270 11620 12310 11660
rect 12380 12120 12420 12160
rect 12380 12020 12420 12060
rect 12380 11920 12420 11960
rect 12380 11820 12420 11860
rect 12380 11720 12420 11760
rect 12380 11620 12420 11660
rect 11230 11230 11270 11270
rect 11230 11130 11270 11170
rect 11230 11030 11270 11070
rect 11230 10930 11270 10970
rect 11610 11230 11650 11270
rect 11610 11130 11650 11170
rect 11610 11030 11650 11070
rect 11610 10930 11650 10970
rect 11750 11230 11790 11270
rect 11750 11130 11790 11170
rect 11750 11030 11790 11070
rect 11750 10930 11790 10970
rect 12130 11230 12170 11270
rect 12130 11130 12170 11170
rect 12130 11030 12170 11070
rect 12130 10930 12170 10970
rect 12270 11230 12310 11270
rect 12270 11130 12310 11170
rect 12270 11030 12310 11070
rect 12270 10930 12310 10970
rect 12650 11230 12690 11270
rect 12650 11130 12690 11170
rect 12650 11030 12690 11070
rect 12650 10930 12690 10970
rect 12790 11230 12830 11270
rect 12790 11130 12830 11170
rect 12790 11030 12830 11070
rect 12790 10930 12830 10970
rect 13170 11230 13210 11270
rect 13170 11130 13210 11170
rect 13170 11030 13210 11070
rect 13170 10930 13210 10970
rect 1280 9750 1320 9790
rect 1280 9650 1320 9690
rect 1280 9550 1320 9590
rect 1280 9450 1320 9490
rect 1390 9750 1430 9790
rect 1390 9650 1430 9690
rect 1390 9550 1430 9590
rect 1390 9450 1430 9490
rect 1500 9750 1540 9790
rect 1500 9650 1540 9690
rect 1500 9550 1540 9590
rect 1500 9450 1540 9490
rect 1800 9750 1840 9790
rect 1800 9650 1840 9690
rect 1800 9550 1840 9590
rect 1800 9450 1840 9490
rect 1910 9750 1950 9790
rect 1910 9650 1950 9690
rect 1910 9550 1950 9590
rect 1910 9450 1950 9490
rect 2020 9750 2060 9790
rect 2180 9750 2220 9790
rect 2020 9650 2060 9690
rect 2180 9650 2220 9690
rect 2020 9550 2060 9590
rect 2180 9550 2220 9590
rect 2020 9450 2060 9490
rect 2180 9450 2220 9490
rect 2290 9750 2330 9790
rect 2290 9650 2330 9690
rect 2290 9550 2330 9590
rect 2290 9450 2330 9490
rect 2400 9750 2440 9790
rect 2400 9650 2440 9690
rect 2400 9550 2440 9590
rect 2400 9450 2440 9490
rect 2700 9750 2740 9790
rect 2700 9650 2740 9690
rect 2700 9550 2740 9590
rect 2700 9450 2740 9490
rect 2810 9750 2850 9790
rect 2810 9650 2850 9690
rect 2810 9550 2850 9590
rect 2810 9450 2850 9490
rect 2920 9750 2960 9790
rect 2920 9650 2960 9690
rect 2920 9550 2960 9590
rect 2920 9450 2960 9490
rect 3220 9750 3260 9790
rect 3220 9650 3260 9690
rect 3220 9550 3260 9590
rect 3220 9450 3260 9490
rect 3330 9750 3370 9790
rect 3330 9650 3370 9690
rect 3330 9550 3370 9590
rect 3330 9450 3370 9490
rect 3440 9750 3480 9790
rect 3440 9650 3480 9690
rect 3440 9550 3480 9590
rect 3440 9450 3480 9490
rect 3660 9750 3700 9790
rect 3660 9650 3700 9690
rect 3660 9550 3700 9590
rect 3660 9450 3700 9490
rect 3770 9750 3810 9790
rect 3770 9650 3810 9690
rect 3770 9550 3810 9590
rect 3770 9450 3810 9490
rect 3990 9750 4030 9790
rect 3990 9650 4030 9690
rect 3990 9550 4030 9590
rect 3990 9450 4030 9490
rect 4100 9750 4140 9790
rect 4100 9650 4140 9690
rect 4100 9550 4140 9590
rect 4100 9450 4140 9490
rect 4420 9750 4460 9790
rect 4420 9650 4460 9690
rect 4420 9550 4460 9590
rect 4420 9450 4460 9490
rect 4550 9750 4590 9790
rect 4550 9650 4590 9690
rect 4550 9550 4590 9590
rect 4550 9450 4590 9490
rect 4810 9750 4850 9790
rect 4810 9650 4850 9690
rect 4810 9550 4850 9590
rect 4810 9450 4850 9490
rect 4940 9750 4980 9790
rect 4940 9650 4980 9690
rect 4940 9550 4980 9590
rect 4940 9450 4980 9490
rect 5200 9750 5240 9790
rect 5200 9650 5240 9690
rect 5200 9550 5240 9590
rect 5200 9450 5240 9490
rect 5330 9750 5370 9790
rect 5330 9650 5370 9690
rect 5330 9550 5370 9590
rect 5330 9450 5370 9490
rect 5490 9750 5530 9790
rect 5490 9650 5530 9690
rect 5490 9550 5530 9590
rect 5490 9450 5530 9490
rect 5620 9750 5660 9790
rect 5620 9650 5660 9690
rect 5620 9550 5660 9590
rect 5620 9450 5660 9490
rect 5880 9750 5920 9790
rect 5880 9650 5920 9690
rect 5880 9550 5920 9590
rect 5880 9450 5920 9490
rect 6010 9750 6050 9790
rect 6010 9650 6050 9690
rect 6010 9550 6050 9590
rect 6010 9450 6050 9490
rect 7570 9720 7610 9760
rect 7570 9620 7610 9660
rect 7570 9520 7610 9560
rect 7570 9420 7610 9460
rect 7790 9720 7830 9760
rect 7790 9620 7830 9660
rect 7790 9520 7830 9560
rect 7790 9420 7830 9460
rect 8010 9720 8050 9760
rect 8010 9620 8050 9660
rect 8010 9520 8050 9560
rect 8010 9420 8050 9460
rect 8230 9720 8270 9760
rect 8230 9620 8270 9660
rect 8230 9520 8270 9560
rect 8230 9420 8270 9460
rect 8450 9720 8490 9760
rect 8450 9620 8490 9660
rect 8450 9520 8490 9560
rect 8450 9420 8490 9460
rect 8670 9720 8710 9760
rect 8670 9620 8710 9660
rect 8670 9520 8710 9560
rect 8670 9420 8710 9460
rect 8890 9720 8930 9760
rect 9090 9720 9130 9760
rect 8890 9620 8930 9660
rect 9090 9620 9130 9660
rect 8890 9520 8930 9560
rect 9090 9520 9130 9560
rect 8890 9420 8930 9460
rect 9090 9420 9130 9460
rect 9310 9720 9350 9760
rect 9310 9620 9350 9660
rect 9310 9520 9350 9560
rect 9310 9420 9350 9460
rect 9530 9720 9570 9760
rect 9530 9620 9570 9660
rect 9530 9520 9570 9560
rect 9530 9420 9570 9460
rect 9750 9720 9790 9760
rect 9750 9620 9790 9660
rect 9750 9520 9790 9560
rect 9750 9420 9790 9460
rect 9970 9720 10010 9760
rect 9970 9620 10010 9660
rect 9970 9520 10010 9560
rect 9970 9420 10010 9460
rect 10190 9720 10230 9760
rect 10190 9620 10230 9660
rect 10190 9520 10230 9560
rect 10190 9420 10230 9460
rect 10410 9720 10450 9760
rect 10410 9620 10450 9660
rect 10410 9520 10450 9560
rect 10410 9420 10450 9460
rect 1280 8990 1320 9030
rect 1280 8890 1320 8930
rect 1280 8790 1320 8830
rect 1280 8690 1320 8730
rect 1390 8990 1430 9030
rect 1390 8890 1430 8930
rect 1390 8790 1430 8830
rect 1390 8690 1430 8730
rect 1500 8990 1540 9030
rect 1500 8890 1540 8930
rect 1500 8790 1540 8830
rect 1500 8690 1540 8730
rect 1800 8990 1840 9030
rect 1800 8890 1840 8930
rect 1800 8790 1840 8830
rect 1800 8690 1840 8730
rect 1910 8990 1950 9030
rect 1910 8890 1950 8930
rect 1910 8790 1950 8830
rect 1910 8690 1950 8730
rect 2020 8990 2060 9030
rect 2180 8990 2220 9030
rect 2020 8890 2060 8930
rect 2180 8890 2220 8930
rect 2020 8790 2060 8830
rect 2180 8790 2220 8830
rect 2020 8690 2060 8730
rect 2180 8690 2220 8730
rect 2290 8990 2330 9030
rect 2290 8890 2330 8930
rect 2290 8790 2330 8830
rect 2290 8690 2330 8730
rect 2400 8990 2440 9030
rect 2400 8890 2440 8930
rect 2400 8790 2440 8830
rect 2400 8690 2440 8730
rect 2700 8990 2740 9030
rect 2700 8890 2740 8930
rect 2700 8790 2740 8830
rect 2700 8690 2740 8730
rect 2810 8990 2850 9030
rect 2810 8890 2850 8930
rect 2810 8790 2850 8830
rect 2810 8690 2850 8730
rect 2920 8990 2960 9030
rect 2920 8890 2960 8930
rect 2920 8790 2960 8830
rect 2920 8690 2960 8730
rect 3210 8990 3250 9030
rect 3210 8890 3250 8930
rect 3210 8790 3250 8830
rect 3210 8690 3250 8730
rect 3320 8990 3360 9030
rect 3320 8890 3360 8930
rect 3320 8790 3360 8830
rect 3320 8690 3360 8730
rect 3540 8990 3580 9030
rect 3540 8890 3580 8930
rect 3540 8790 3580 8830
rect 3540 8690 3580 8730
rect 3650 8990 3690 9030
rect 3650 8890 3690 8930
rect 3650 8790 3690 8830
rect 3650 8690 3690 8730
rect 3870 8990 3910 9030
rect 3870 8890 3910 8930
rect 3870 8790 3910 8830
rect 3870 8690 3910 8730
rect 3980 8990 4020 9030
rect 3980 8890 4020 8930
rect 3980 8790 4020 8830
rect 3980 8690 4020 8730
rect 4420 8990 4460 9030
rect 4420 8890 4460 8930
rect 4420 8790 4460 8830
rect 4420 8690 4460 8730
rect 4550 8990 4590 9030
rect 4550 8890 4590 8930
rect 4550 8790 4590 8830
rect 4550 8690 4590 8730
rect 4810 8990 4850 9030
rect 4810 8890 4850 8930
rect 4810 8790 4850 8830
rect 4810 8690 4850 8730
rect 4940 8990 4980 9030
rect 4940 8890 4980 8930
rect 4940 8790 4980 8830
rect 4940 8690 4980 8730
rect 5200 8990 5240 9030
rect 5200 8890 5240 8930
rect 5200 8790 5240 8830
rect 5200 8690 5240 8730
rect 5330 8990 5370 9030
rect 5330 8890 5370 8930
rect 5330 8790 5370 8830
rect 5330 8690 5370 8730
rect 5490 8990 5530 9030
rect 5490 8890 5530 8930
rect 5490 8790 5530 8830
rect 5490 8690 5530 8730
rect 5620 8990 5660 9030
rect 5620 8890 5660 8930
rect 5620 8790 5660 8830
rect 5620 8690 5660 8730
rect -340 6800 -300 6840
rect -340 6700 -300 6740
rect -230 6800 -190 6840
rect -230 6700 -190 6740
rect -120 6800 -80 6840
rect -120 6700 -80 6740
rect -10 6800 30 6840
rect -10 6700 30 6740
rect 100 6800 140 6840
rect 100 6700 140 6740
rect 210 6800 250 6840
rect 210 6700 250 6740
rect 320 6800 360 6840
rect 320 6700 360 6740
rect 430 6800 470 6840
rect 430 6700 470 6740
rect 540 6800 580 6840
rect 540 6700 580 6740
rect 650 6800 690 6840
rect 650 6700 690 6740
rect 760 6800 800 6840
rect 760 6700 800 6740
rect 870 6800 910 6840
rect 870 6700 910 6740
rect 980 6800 1020 6840
rect 980 6700 1020 6740
rect 1560 6800 1600 6840
rect 1560 6700 1600 6740
rect 1670 6800 1710 6840
rect 1670 6700 1710 6740
rect 1780 6800 1820 6840
rect 1780 6700 1820 6740
rect 1890 6800 1930 6840
rect 1890 6700 1930 6740
rect 2000 6800 2040 6840
rect 2000 6700 2040 6740
rect 2110 6800 2150 6840
rect 2110 6700 2150 6740
rect 2220 6800 2260 6840
rect 2220 6700 2260 6740
rect 2330 6800 2370 6840
rect 2330 6700 2370 6740
rect 2440 6800 2480 6840
rect 2440 6700 2480 6740
rect 2550 6800 2590 6840
rect 2550 6700 2590 6740
rect 2660 6800 2700 6840
rect 2660 6700 2700 6740
rect 2770 6800 2810 6840
rect 2770 6700 2810 6740
rect 2880 6800 2920 6840
rect 2880 6700 2920 6740
rect -350 6200 -310 6240
rect -350 6100 -310 6140
rect -350 6000 -310 6040
rect -350 5900 -310 5940
rect -350 5800 -310 5840
rect -350 5700 -310 5740
rect -170 6200 -130 6240
rect -170 6100 -130 6140
rect -170 6000 -130 6040
rect -170 5900 -130 5940
rect -170 5800 -130 5840
rect -170 5700 -130 5740
rect 10 6200 50 6240
rect 10 6100 50 6140
rect 10 6000 50 6040
rect 10 5900 50 5940
rect 10 5800 50 5840
rect 10 5700 50 5740
rect 190 6200 230 6240
rect 190 6100 230 6140
rect 190 6000 230 6040
rect 190 5900 230 5940
rect 190 5800 230 5840
rect 190 5700 230 5740
rect 370 6200 410 6240
rect 370 6100 410 6140
rect 370 6000 410 6040
rect 370 5900 410 5940
rect 370 5800 410 5840
rect 370 5700 410 5740
rect 550 6200 590 6240
rect 550 6100 590 6140
rect 550 6000 590 6040
rect 550 5900 590 5940
rect 550 5800 590 5840
rect 550 5700 590 5740
rect 730 6200 770 6240
rect 730 6100 770 6140
rect 730 6000 770 6040
rect 730 5900 770 5940
rect 730 5800 770 5840
rect 730 5700 770 5740
rect 910 6200 950 6240
rect 910 6100 950 6140
rect 910 6000 950 6040
rect 910 5900 950 5940
rect 910 5800 950 5840
rect 910 5700 950 5740
rect 1090 6200 1130 6240
rect 1090 6100 1130 6140
rect 1090 6000 1130 6040
rect 1090 5900 1130 5940
rect 1090 5800 1130 5840
rect 1090 5700 1130 5740
rect 1270 6200 1310 6240
rect 1270 6100 1310 6140
rect 1270 6000 1310 6040
rect 1270 5900 1310 5940
rect 1270 5800 1310 5840
rect 1270 5700 1310 5740
rect 1450 6200 1490 6240
rect 1450 6100 1490 6140
rect 1450 6000 1490 6040
rect 1450 5900 1490 5940
rect 1450 5800 1490 5840
rect 1450 5700 1490 5740
rect 1630 6200 1670 6240
rect 1630 6100 1670 6140
rect 1630 6000 1670 6040
rect 1630 5900 1670 5940
rect 1630 5800 1670 5840
rect 1630 5700 1670 5740
rect 1810 6200 1850 6240
rect 1810 6100 1850 6140
rect 1810 6000 1850 6040
rect 1810 5900 1850 5940
rect 1810 5800 1850 5840
rect 1810 5700 1850 5740
rect 1990 6200 2030 6240
rect 1990 6100 2030 6140
rect 1990 6000 2030 6040
rect 1990 5900 2030 5940
rect 1990 5800 2030 5840
rect 1990 5700 2030 5740
rect 2170 6200 2210 6240
rect 2170 6100 2210 6140
rect 2170 6000 2210 6040
rect 2170 5900 2210 5940
rect 2170 5800 2210 5840
rect 2170 5700 2210 5740
rect 2350 6200 2390 6240
rect 2350 6100 2390 6140
rect 2350 6000 2390 6040
rect 2350 5900 2390 5940
rect 2350 5800 2390 5840
rect 2350 5700 2390 5740
rect 2530 6200 2570 6240
rect 2530 6100 2570 6140
rect 2530 6000 2570 6040
rect 2530 5900 2570 5940
rect 2530 5800 2570 5840
rect 2530 5700 2570 5740
rect 2710 6200 2750 6240
rect 2710 6100 2750 6140
rect 2710 6000 2750 6040
rect 2710 5900 2750 5940
rect 2710 5800 2750 5840
rect 2710 5700 2750 5740
rect 2890 6200 2930 6240
rect 2890 6100 2930 6140
rect 2890 6000 2930 6040
rect 2890 5900 2930 5940
rect 3520 6000 3560 6040
rect 3520 5900 3560 5940
rect 3630 6000 3670 6040
rect 3630 5900 3670 5940
rect 3740 6000 3780 6040
rect 3740 5900 3780 5940
rect 3850 6000 3890 6040
rect 3850 5900 3890 5940
rect 3960 6000 4000 6040
rect 3960 5900 4000 5940
rect 2890 5800 2930 5840
rect 2890 5700 2930 5740
rect 7480 4720 7520 4760
rect -1450 4640 -1410 4680
rect -1450 4540 -1410 4580
rect -1330 4640 -1290 4680
rect -1330 4540 -1290 4580
rect -1210 4640 -1170 4680
rect -1210 4540 -1170 4580
rect -1090 4640 -1050 4680
rect -1090 4540 -1050 4580
rect -970 4640 -930 4680
rect -970 4540 -930 4580
rect -850 4640 -810 4680
rect -850 4540 -810 4580
rect -730 4640 -690 4680
rect -730 4540 -690 4580
rect -610 4640 -570 4680
rect -610 4540 -570 4580
rect -490 4640 -450 4680
rect -490 4540 -450 4580
rect -370 4640 -330 4680
rect -370 4540 -330 4580
rect -250 4640 -210 4680
rect -250 4540 -210 4580
rect -130 4640 -90 4680
rect -130 4540 -90 4580
rect -10 4640 30 4680
rect -10 4540 30 4580
rect 110 4640 150 4680
rect 110 4540 150 4580
rect 230 4640 270 4680
rect 230 4540 270 4580
rect 350 4640 390 4680
rect 350 4540 390 4580
rect 470 4640 510 4680
rect 470 4540 510 4580
rect 590 4640 630 4680
rect 590 4540 630 4580
rect 710 4640 750 4680
rect 710 4540 750 4580
rect 830 4640 870 4680
rect 830 4540 870 4580
rect 950 4640 990 4680
rect 950 4540 990 4580
rect 1590 4640 1630 4680
rect 1590 4540 1630 4580
rect 1710 4640 1750 4680
rect 1710 4540 1750 4580
rect 1830 4640 1870 4680
rect 1830 4540 1870 4580
rect 1950 4640 1990 4680
rect 1950 4540 1990 4580
rect 2070 4640 2110 4680
rect 2070 4540 2110 4580
rect 2190 4640 2230 4680
rect 2190 4540 2230 4580
rect 2310 4640 2350 4680
rect 2310 4540 2350 4580
rect 2430 4640 2470 4680
rect 2430 4540 2470 4580
rect 2550 4640 2590 4680
rect 2550 4540 2590 4580
rect 2670 4640 2710 4680
rect 2670 4540 2710 4580
rect 2790 4640 2830 4680
rect 2790 4540 2830 4580
rect 2910 4640 2950 4680
rect 2910 4540 2950 4580
rect 3030 4640 3070 4680
rect 3030 4540 3070 4580
rect 3150 4640 3190 4680
rect 3150 4540 3190 4580
rect 3270 4640 3310 4680
rect 3270 4540 3310 4580
rect 3390 4640 3430 4680
rect 3390 4540 3430 4580
rect 3510 4640 3550 4680
rect 3510 4540 3550 4580
rect 3630 4640 3670 4680
rect 3630 4540 3670 4580
rect 3750 4640 3790 4680
rect 3750 4540 3790 4580
rect 3870 4640 3910 4680
rect 3870 4540 3910 4580
rect 3990 4640 4030 4680
rect 7480 4620 7520 4660
rect 7610 4720 7650 4760
rect 7610 4620 7650 4660
rect 7740 4720 7780 4760
rect 7740 4620 7780 4660
rect 7870 4720 7910 4760
rect 7870 4620 7910 4660
rect 8000 4720 8040 4760
rect 8000 4620 8040 4660
rect 8130 4720 8170 4760
rect 8130 4620 8170 4660
rect 8260 4720 8300 4760
rect 8260 4620 8300 4660
rect 8620 4720 8660 4760
rect 8620 4620 8660 4660
rect 8750 4720 8790 4760
rect 8750 4620 8790 4660
rect 8880 4720 8920 4760
rect 8880 4620 8920 4660
rect 9010 4720 9050 4760
rect 9010 4620 9050 4660
rect 9140 4720 9180 4760
rect 9140 4620 9180 4660
rect 9270 4720 9310 4760
rect 9270 4620 9310 4660
rect 9400 4720 9440 4760
rect 9400 4620 9440 4660
rect 9760 4720 9800 4760
rect 9760 4620 9800 4660
rect 9890 4720 9930 4760
rect 9890 4620 9930 4660
rect 10020 4720 10060 4760
rect 10020 4620 10060 4660
rect 10150 4720 10190 4760
rect 10150 4620 10190 4660
rect 10280 4720 10320 4760
rect 10280 4620 10320 4660
rect 10410 4720 10450 4760
rect 10410 4620 10450 4660
rect 10540 4720 10580 4760
rect 10540 4620 10580 4660
rect 3990 4540 4030 4580
rect 7550 4070 7590 4110
rect 7550 3970 7590 4010
rect 7550 3870 7590 3910
rect 7550 3770 7590 3810
rect 7550 3670 7590 3710
rect 7750 4070 7790 4110
rect 7750 3970 7790 4010
rect 7750 3870 7790 3910
rect 7750 3770 7790 3810
rect 7750 3670 7790 3710
rect 7950 4070 7990 4110
rect 7950 3970 7990 4010
rect 7950 3870 7990 3910
rect 7950 3770 7990 3810
rect 7950 3670 7990 3710
rect 8150 4070 8190 4110
rect 8150 3970 8190 4010
rect 8150 3870 8190 3910
rect 8150 3770 8190 3810
rect 8150 3670 8190 3710
rect 8350 4070 8390 4110
rect 8350 3970 8390 4010
rect 8350 3870 8390 3910
rect 8350 3770 8390 3810
rect 8350 3670 8390 3710
rect 8550 4070 8590 4110
rect 8550 3970 8590 4010
rect 8550 3870 8590 3910
rect 8550 3770 8590 3810
rect 8550 3670 8590 3710
rect 8750 4070 8790 4110
rect 8750 3970 8790 4010
rect 8750 3870 8790 3910
rect 8750 3770 8790 3810
rect 8750 3670 8790 3710
rect 8950 4070 8990 4110
rect 8950 3970 8990 4010
rect 8950 3870 8990 3910
rect 8950 3770 8990 3810
rect 8950 3670 8990 3710
rect 9150 4070 9190 4110
rect 9150 3970 9190 4010
rect 9150 3870 9190 3910
rect 9150 3770 9190 3810
rect 9150 3670 9190 3710
rect 9350 4070 9390 4110
rect 9350 3970 9390 4010
rect 9350 3870 9390 3910
rect 9350 3770 9390 3810
rect 9350 3670 9390 3710
rect 9550 4070 9590 4110
rect 9550 3970 9590 4010
rect 9550 3870 9590 3910
rect 9550 3770 9590 3810
rect 9550 3670 9590 3710
rect -358 1164 -324 1198
rect -268 1164 -234 1198
rect -178 1164 -144 1198
rect -88 1164 -54 1198
rect 2 1164 36 1198
rect 92 1164 126 1198
rect 182 1164 216 1198
rect -358 1074 -324 1108
rect -268 1074 -234 1108
rect -178 1074 -144 1108
rect -88 1074 -54 1108
rect 2 1074 36 1108
rect 92 1074 126 1108
rect 182 1074 216 1108
rect -358 984 -324 1018
rect -268 984 -234 1018
rect -178 984 -144 1018
rect -88 984 -54 1018
rect 2 984 36 1018
rect 92 984 126 1018
rect 182 984 216 1018
rect -358 894 -324 928
rect -268 894 -234 928
rect -178 894 -144 928
rect -88 894 -54 928
rect 2 894 36 928
rect 92 894 126 928
rect 182 894 216 928
rect -358 804 -324 838
rect -268 804 -234 838
rect -178 804 -144 838
rect -88 804 -54 838
rect 2 804 36 838
rect 92 804 126 838
rect 182 804 216 838
rect -358 714 -324 748
rect -268 714 -234 748
rect -178 714 -144 748
rect -88 714 -54 748
rect 2 714 36 748
rect 92 714 126 748
rect 182 714 216 748
rect -358 624 -324 658
rect -268 624 -234 658
rect -178 624 -144 658
rect -88 624 -54 658
rect 2 624 36 658
rect 92 624 126 658
rect 182 624 216 658
rect 1002 1164 1036 1198
rect 1092 1164 1126 1198
rect 1182 1164 1216 1198
rect 1272 1164 1306 1198
rect 1362 1164 1396 1198
rect 1452 1164 1486 1198
rect 1542 1164 1576 1198
rect 1002 1074 1036 1108
rect 1092 1074 1126 1108
rect 1182 1074 1216 1108
rect 1272 1074 1306 1108
rect 1362 1074 1396 1108
rect 1452 1074 1486 1108
rect 1542 1074 1576 1108
rect 1002 984 1036 1018
rect 1092 984 1126 1018
rect 1182 984 1216 1018
rect 1272 984 1306 1018
rect 1362 984 1396 1018
rect 1452 984 1486 1018
rect 1542 984 1576 1018
rect 1002 894 1036 928
rect 1092 894 1126 928
rect 1182 894 1216 928
rect 1272 894 1306 928
rect 1362 894 1396 928
rect 1452 894 1486 928
rect 1542 894 1576 928
rect 1002 804 1036 838
rect 1092 804 1126 838
rect 1182 804 1216 838
rect 1272 804 1306 838
rect 1362 804 1396 838
rect 1452 804 1486 838
rect 1542 804 1576 838
rect 1002 714 1036 748
rect 1092 714 1126 748
rect 1182 714 1216 748
rect 1272 714 1306 748
rect 1362 714 1396 748
rect 1452 714 1486 748
rect 1542 714 1576 748
rect 1002 624 1036 658
rect 1092 624 1126 658
rect 1182 624 1216 658
rect 1272 624 1306 658
rect 1362 624 1396 658
rect 1452 624 1486 658
rect 1542 624 1576 658
rect 2362 1164 2396 1198
rect 2452 1164 2486 1198
rect 2542 1164 2576 1198
rect 2632 1164 2666 1198
rect 2722 1164 2756 1198
rect 2812 1164 2846 1198
rect 2902 1164 2936 1198
rect 2362 1074 2396 1108
rect 2452 1074 2486 1108
rect 2542 1074 2576 1108
rect 2632 1074 2666 1108
rect 2722 1074 2756 1108
rect 2812 1074 2846 1108
rect 2902 1074 2936 1108
rect 2362 984 2396 1018
rect 2452 984 2486 1018
rect 2542 984 2576 1018
rect 2632 984 2666 1018
rect 2722 984 2756 1018
rect 2812 984 2846 1018
rect 2902 984 2936 1018
rect 2362 894 2396 928
rect 2452 894 2486 928
rect 2542 894 2576 928
rect 2632 894 2666 928
rect 2722 894 2756 928
rect 2812 894 2846 928
rect 2902 894 2936 928
rect 2362 804 2396 838
rect 2452 804 2486 838
rect 2542 804 2576 838
rect 2632 804 2666 838
rect 2722 804 2756 838
rect 2812 804 2846 838
rect 2902 804 2936 838
rect 2362 714 2396 748
rect 2452 714 2486 748
rect 2542 714 2576 748
rect 2632 714 2666 748
rect 2722 714 2756 748
rect 2812 714 2846 748
rect 2902 714 2936 748
rect 2362 624 2396 658
rect 2452 624 2486 658
rect 2542 624 2576 658
rect 2632 624 2666 658
rect 2722 624 2756 658
rect 2812 624 2846 658
rect 2902 624 2936 658
rect -358 -196 -324 -162
rect -268 -196 -234 -162
rect -178 -196 -144 -162
rect -88 -196 -54 -162
rect 2 -196 36 -162
rect 92 -196 126 -162
rect 182 -196 216 -162
rect -358 -286 -324 -252
rect -268 -286 -234 -252
rect -178 -286 -144 -252
rect -88 -286 -54 -252
rect 2 -286 36 -252
rect 92 -286 126 -252
rect 182 -286 216 -252
rect -358 -376 -324 -342
rect -268 -376 -234 -342
rect -178 -376 -144 -342
rect -88 -376 -54 -342
rect 2 -376 36 -342
rect 92 -376 126 -342
rect 182 -376 216 -342
rect -358 -466 -324 -432
rect -268 -466 -234 -432
rect -178 -466 -144 -432
rect -88 -466 -54 -432
rect 2 -466 36 -432
rect 92 -466 126 -432
rect 182 -466 216 -432
rect -358 -556 -324 -522
rect -268 -556 -234 -522
rect -178 -556 -144 -522
rect -88 -556 -54 -522
rect 2 -556 36 -522
rect 92 -556 126 -522
rect 182 -556 216 -522
rect -358 -646 -324 -612
rect -268 -646 -234 -612
rect -178 -646 -144 -612
rect -88 -646 -54 -612
rect 2 -646 36 -612
rect 92 -646 126 -612
rect 182 -646 216 -612
rect -358 -736 -324 -702
rect -268 -736 -234 -702
rect -178 -736 -144 -702
rect -88 -736 -54 -702
rect 2 -736 36 -702
rect 92 -736 126 -702
rect 182 -736 216 -702
rect 1002 -196 1036 -162
rect 1092 -196 1126 -162
rect 1182 -196 1216 -162
rect 1272 -196 1306 -162
rect 1362 -196 1396 -162
rect 1452 -196 1486 -162
rect 1542 -196 1576 -162
rect 1002 -286 1036 -252
rect 1092 -286 1126 -252
rect 1182 -286 1216 -252
rect 1272 -286 1306 -252
rect 1362 -286 1396 -252
rect 1452 -286 1486 -252
rect 1542 -286 1576 -252
rect 1002 -376 1036 -342
rect 1092 -376 1126 -342
rect 1182 -376 1216 -342
rect 1272 -376 1306 -342
rect 1362 -376 1396 -342
rect 1452 -376 1486 -342
rect 1542 -376 1576 -342
rect 1002 -466 1036 -432
rect 1092 -466 1126 -432
rect 1182 -466 1216 -432
rect 1272 -466 1306 -432
rect 1362 -466 1396 -432
rect 1452 -466 1486 -432
rect 1542 -466 1576 -432
rect 1002 -556 1036 -522
rect 1092 -556 1126 -522
rect 1182 -556 1216 -522
rect 1272 -556 1306 -522
rect 1362 -556 1396 -522
rect 1452 -556 1486 -522
rect 1542 -556 1576 -522
rect 1002 -646 1036 -612
rect 1092 -646 1126 -612
rect 1182 -646 1216 -612
rect 1272 -646 1306 -612
rect 1362 -646 1396 -612
rect 1452 -646 1486 -612
rect 1542 -646 1576 -612
rect 1002 -736 1036 -702
rect 1092 -736 1126 -702
rect 1182 -736 1216 -702
rect 1272 -736 1306 -702
rect 1362 -736 1396 -702
rect 1452 -736 1486 -702
rect 1542 -736 1576 -702
rect 2362 -196 2396 -162
rect 2452 -196 2486 -162
rect 2542 -196 2576 -162
rect 2632 -196 2666 -162
rect 2722 -196 2756 -162
rect 2812 -196 2846 -162
rect 2902 -196 2936 -162
rect 2362 -286 2396 -252
rect 2452 -286 2486 -252
rect 2542 -286 2576 -252
rect 2632 -286 2666 -252
rect 2722 -286 2756 -252
rect 2812 -286 2846 -252
rect 2902 -286 2936 -252
rect 2362 -376 2396 -342
rect 2452 -376 2486 -342
rect 2542 -376 2576 -342
rect 2632 -376 2666 -342
rect 2722 -376 2756 -342
rect 2812 -376 2846 -342
rect 2902 -376 2936 -342
rect 2362 -466 2396 -432
rect 2452 -466 2486 -432
rect 2542 -466 2576 -432
rect 2632 -466 2666 -432
rect 2722 -466 2756 -432
rect 2812 -466 2846 -432
rect 2902 -466 2936 -432
rect 2362 -556 2396 -522
rect 2452 -556 2486 -522
rect 2542 -556 2576 -522
rect 2632 -556 2666 -522
rect 2722 -556 2756 -522
rect 2812 -556 2846 -522
rect 2902 -556 2936 -522
rect 2362 -646 2396 -612
rect 2452 -646 2486 -612
rect 2542 -646 2576 -612
rect 2632 -646 2666 -612
rect 2722 -646 2756 -612
rect 2812 -646 2846 -612
rect 2902 -646 2936 -612
rect 2362 -736 2396 -702
rect 2452 -736 2486 -702
rect 2542 -736 2576 -702
rect 2632 -736 2666 -702
rect 2722 -736 2756 -702
rect 2812 -736 2846 -702
rect 2902 -736 2936 -702
rect -358 -1556 -324 -1522
rect -268 -1556 -234 -1522
rect -178 -1556 -144 -1522
rect -88 -1556 -54 -1522
rect 2 -1556 36 -1522
rect 92 -1556 126 -1522
rect 182 -1556 216 -1522
rect -358 -1646 -324 -1612
rect -268 -1646 -234 -1612
rect -178 -1646 -144 -1612
rect -88 -1646 -54 -1612
rect 2 -1646 36 -1612
rect 92 -1646 126 -1612
rect 182 -1646 216 -1612
rect -358 -1736 -324 -1702
rect -268 -1736 -234 -1702
rect -178 -1736 -144 -1702
rect -88 -1736 -54 -1702
rect 2 -1736 36 -1702
rect 92 -1736 126 -1702
rect 182 -1736 216 -1702
rect -358 -1826 -324 -1792
rect -268 -1826 -234 -1792
rect -178 -1826 -144 -1792
rect -88 -1826 -54 -1792
rect 2 -1826 36 -1792
rect 92 -1826 126 -1792
rect 182 -1826 216 -1792
rect -358 -1916 -324 -1882
rect -268 -1916 -234 -1882
rect -178 -1916 -144 -1882
rect -88 -1916 -54 -1882
rect 2 -1916 36 -1882
rect 92 -1916 126 -1882
rect 182 -1916 216 -1882
rect -358 -2006 -324 -1972
rect -268 -2006 -234 -1972
rect -178 -2006 -144 -1972
rect -88 -2006 -54 -1972
rect 2 -2006 36 -1972
rect 92 -2006 126 -1972
rect 182 -2006 216 -1972
rect -358 -2096 -324 -2062
rect -268 -2096 -234 -2062
rect -178 -2096 -144 -2062
rect -88 -2096 -54 -2062
rect 2 -2096 36 -2062
rect 92 -2096 126 -2062
rect 182 -2096 216 -2062
rect 1002 -1556 1036 -1522
rect 1092 -1556 1126 -1522
rect 1182 -1556 1216 -1522
rect 1272 -1556 1306 -1522
rect 1362 -1556 1396 -1522
rect 1452 -1556 1486 -1522
rect 1542 -1556 1576 -1522
rect 1002 -1646 1036 -1612
rect 1092 -1646 1126 -1612
rect 1182 -1646 1216 -1612
rect 1272 -1646 1306 -1612
rect 1362 -1646 1396 -1612
rect 1452 -1646 1486 -1612
rect 1542 -1646 1576 -1612
rect 1002 -1736 1036 -1702
rect 1092 -1736 1126 -1702
rect 1182 -1736 1216 -1702
rect 1272 -1736 1306 -1702
rect 1362 -1736 1396 -1702
rect 1452 -1736 1486 -1702
rect 1542 -1736 1576 -1702
rect 1002 -1826 1036 -1792
rect 1092 -1826 1126 -1792
rect 1182 -1826 1216 -1792
rect 1272 -1826 1306 -1792
rect 1362 -1826 1396 -1792
rect 1452 -1826 1486 -1792
rect 1542 -1826 1576 -1792
rect 1002 -1916 1036 -1882
rect 1092 -1916 1126 -1882
rect 1182 -1916 1216 -1882
rect 1272 -1916 1306 -1882
rect 1362 -1916 1396 -1882
rect 1452 -1916 1486 -1882
rect 1542 -1916 1576 -1882
rect 1002 -2006 1036 -1972
rect 1092 -2006 1126 -1972
rect 1182 -2006 1216 -1972
rect 1272 -2006 1306 -1972
rect 1362 -2006 1396 -1972
rect 1452 -2006 1486 -1972
rect 1542 -2006 1576 -1972
rect 1002 -2096 1036 -2062
rect 1092 -2096 1126 -2062
rect 1182 -2096 1216 -2062
rect 1272 -2096 1306 -2062
rect 1362 -2096 1396 -2062
rect 1452 -2096 1486 -2062
rect 1542 -2096 1576 -2062
rect 2362 -1556 2396 -1522
rect 2452 -1556 2486 -1522
rect 2542 -1556 2576 -1522
rect 2632 -1556 2666 -1522
rect 2722 -1556 2756 -1522
rect 2812 -1556 2846 -1522
rect 2902 -1556 2936 -1522
rect 2362 -1646 2396 -1612
rect 2452 -1646 2486 -1612
rect 2542 -1646 2576 -1612
rect 2632 -1646 2666 -1612
rect 2722 -1646 2756 -1612
rect 2812 -1646 2846 -1612
rect 2902 -1646 2936 -1612
rect 2362 -1736 2396 -1702
rect 2452 -1736 2486 -1702
rect 2542 -1736 2576 -1702
rect 2632 -1736 2666 -1702
rect 2722 -1736 2756 -1702
rect 2812 -1736 2846 -1702
rect 2902 -1736 2936 -1702
rect 2362 -1826 2396 -1792
rect 2452 -1826 2486 -1792
rect 2542 -1826 2576 -1792
rect 2632 -1826 2666 -1792
rect 2722 -1826 2756 -1792
rect 2812 -1826 2846 -1792
rect 2902 -1826 2936 -1792
rect 2362 -1916 2396 -1882
rect 2452 -1916 2486 -1882
rect 2542 -1916 2576 -1882
rect 2632 -1916 2666 -1882
rect 2722 -1916 2756 -1882
rect 2812 -1916 2846 -1882
rect 2902 -1916 2936 -1882
rect 2362 -2006 2396 -1972
rect 2452 -2006 2486 -1972
rect 2542 -2006 2576 -1972
rect 2632 -2006 2666 -1972
rect 2722 -2006 2756 -1972
rect 2812 -2006 2846 -1972
rect 2902 -2006 2936 -1972
rect 2362 -2096 2396 -2062
rect 2452 -2096 2486 -2062
rect 2542 -2096 2576 -2062
rect 2632 -2096 2666 -2062
rect 2722 -2096 2756 -2062
rect 2812 -2096 2846 -2062
rect 2902 -2096 2936 -2062
<< psubdiff >>
rect 11100 14410 12240 14450
rect 12380 14410 13140 14450
rect 11100 13880 11140 14410
rect 13100 13880 13140 14410
rect 6930 13280 7010 13310
rect 6930 13240 6950 13280
rect 6990 13240 7010 13280
rect 3690 13190 3770 13220
rect 3690 13150 3710 13190
rect 3750 13150 3770 13190
rect 3690 13120 3770 13150
rect 5140 13190 5220 13220
rect 5140 13150 5160 13190
rect 5200 13150 5220 13190
rect 5140 13120 5220 13150
rect 6930 13210 7010 13240
rect 8230 13280 8310 13310
rect 8230 13240 8250 13280
rect 8290 13240 8310 13280
rect 8230 13210 8310 13240
rect 9530 13280 9610 13310
rect 9530 13240 9550 13280
rect 9590 13240 9610 13280
rect 9530 13210 9610 13240
rect 11100 13150 11140 13670
rect 13100 13150 13140 13670
rect 11100 13110 12240 13150
rect 12380 13110 13140 13150
rect 1180 10210 1260 10240
rect 1180 10170 1200 10210
rect 1240 10170 1260 10210
rect 1180 10110 1260 10170
rect 1180 10070 1200 10110
rect 1240 10070 1260 10110
rect 1180 10040 1260 10070
rect 2080 10210 2160 10240
rect 2080 10170 2100 10210
rect 2140 10170 2160 10210
rect 2080 10110 2160 10170
rect 2080 10070 2100 10110
rect 2140 10070 2160 10110
rect 2080 10040 2160 10070
rect 2980 10210 3060 10240
rect 2980 10170 3000 10210
rect 3040 10170 3060 10210
rect 2980 10110 3060 10170
rect 2980 10070 3000 10110
rect 3040 10070 3060 10110
rect 2980 10040 3060 10070
rect 3120 10210 3200 10240
rect 3120 10170 3140 10210
rect 3180 10170 3200 10210
rect 3120 10110 3200 10170
rect 3120 10070 3140 10110
rect 3180 10070 3200 10110
rect 3120 10040 3200 10070
rect 3560 10210 3640 10240
rect 3560 10170 3580 10210
rect 3620 10170 3640 10210
rect 3560 10110 3640 10170
rect 3560 10070 3580 10110
rect 3620 10070 3640 10110
rect 3560 10040 3640 10070
rect 3890 10210 3970 10240
rect 3890 10170 3910 10210
rect 3950 10170 3970 10210
rect 3890 10110 3970 10170
rect 3890 10070 3910 10110
rect 3950 10070 3970 10110
rect 3890 10040 3970 10070
rect 4310 10210 4390 10240
rect 4310 10170 4330 10210
rect 4370 10170 4390 10210
rect 4310 10110 4390 10170
rect 4310 10070 4330 10110
rect 4370 10070 4390 10110
rect 4310 10040 4390 10070
rect 4700 10210 4780 10240
rect 4700 10170 4720 10210
rect 4760 10170 4780 10210
rect 4700 10110 4780 10170
rect 4700 10070 4720 10110
rect 4760 10070 4780 10110
rect 4700 10040 4780 10070
rect 5090 10210 5170 10240
rect 5090 10170 5110 10210
rect 5150 10170 5170 10210
rect 5090 10110 5170 10170
rect 5090 10070 5110 10110
rect 5150 10070 5170 10110
rect 5090 10040 5170 10070
rect 7240 8660 7340 8690
rect 7240 8620 7270 8660
rect 7310 8620 7340 8660
rect 7240 8560 7340 8620
rect 7240 8520 7270 8560
rect 7310 8520 7340 8560
rect 7240 8460 7340 8520
rect 1180 8410 1260 8440
rect 1180 8370 1200 8410
rect 1240 8370 1260 8410
rect 1180 8310 1260 8370
rect 1180 8270 1200 8310
rect 1240 8270 1260 8310
rect 1180 8240 1260 8270
rect 2080 8410 2160 8440
rect 2080 8370 2100 8410
rect 2140 8370 2160 8410
rect 2080 8310 2160 8370
rect 2080 8270 2100 8310
rect 2140 8270 2160 8310
rect 2080 8240 2160 8270
rect 2980 8410 3060 8440
rect 2980 8370 3000 8410
rect 3040 8370 3060 8410
rect 2980 8310 3060 8370
rect 2980 8270 3000 8310
rect 3040 8270 3060 8310
rect 2980 8240 3060 8270
rect 3380 8410 3460 8440
rect 3380 8370 3400 8410
rect 3440 8370 3460 8410
rect 3380 8310 3460 8370
rect 3380 8270 3400 8310
rect 3440 8270 3460 8310
rect 3380 8240 3460 8270
rect 3710 8410 3790 8440
rect 3710 8370 3730 8410
rect 3770 8370 3790 8410
rect 3710 8310 3790 8370
rect 3710 8270 3730 8310
rect 3770 8270 3790 8310
rect 3710 8240 3790 8270
rect 4040 8410 4120 8440
rect 4040 8370 4060 8410
rect 4100 8370 4120 8410
rect 4040 8310 4120 8370
rect 4040 8270 4060 8310
rect 4100 8270 4120 8310
rect 4040 8240 4120 8270
rect 4290 8410 4390 8440
rect 4290 8370 4320 8410
rect 4360 8370 4390 8410
rect 4290 8310 4390 8370
rect 4290 8270 4320 8310
rect 4360 8270 4390 8310
rect 4290 8240 4390 8270
rect 5070 8410 5170 8440
rect 5070 8370 5100 8410
rect 5140 8370 5170 8410
rect 5070 8310 5170 8370
rect 5070 8270 5100 8310
rect 5140 8270 5170 8310
rect 5070 8240 5170 8270
rect 5750 8410 5850 8440
rect 5750 8370 5780 8410
rect 5820 8370 5850 8410
rect 5750 8310 5850 8370
rect 5750 8270 5780 8310
rect 5820 8270 5850 8310
rect 5750 8240 5850 8270
rect 7240 8420 7270 8460
rect 7310 8420 7340 8460
rect 7240 8360 7340 8420
rect 7240 8320 7270 8360
rect 7310 8320 7340 8360
rect 7240 8290 7340 8320
rect 8320 8660 8420 8690
rect 8320 8620 8350 8660
rect 8390 8620 8420 8660
rect 8320 8560 8420 8620
rect 8320 8520 8350 8560
rect 8390 8520 8420 8560
rect 8320 8460 8420 8520
rect 8320 8420 8350 8460
rect 8390 8420 8420 8460
rect 8320 8360 8420 8420
rect 8320 8320 8350 8360
rect 8390 8320 8420 8360
rect 8320 8290 8420 8320
rect 9400 8660 9500 8690
rect 9400 8620 9430 8660
rect 9470 8620 9500 8660
rect 9400 8560 9500 8620
rect 9400 8520 9430 8560
rect 9470 8520 9500 8560
rect 9400 8460 9500 8520
rect 9400 8420 9430 8460
rect 9470 8420 9500 8460
rect 9400 8360 9500 8420
rect 9400 8320 9430 8360
rect 9470 8320 9500 8360
rect 9400 8290 9500 8320
rect 10480 8660 10580 8690
rect 10480 8620 10510 8660
rect 10550 8620 10580 8660
rect 10480 8560 10580 8620
rect 10480 8520 10510 8560
rect 10550 8520 10580 8560
rect 10480 8460 10580 8520
rect 10480 8420 10510 8460
rect 10550 8420 10580 8460
rect 10480 8360 10580 8420
rect 10480 8320 10510 8360
rect 10550 8320 10580 8360
rect 10480 8290 10580 8320
rect 7300 6030 7400 6060
rect 7300 5980 7330 6030
rect 7370 5980 7400 6030
rect 7300 5890 7400 5980
rect 7300 5840 7330 5890
rect 7370 5840 7400 5890
rect 7300 5810 7400 5840
rect 9500 6030 9600 6060
rect 9500 5980 9530 6030
rect 9570 5980 9600 6030
rect 9500 5890 9600 5980
rect 9500 5840 9530 5890
rect 9570 5840 9600 5890
rect 9500 5810 9600 5840
rect 7350 5340 7450 5370
rect 7350 5300 7380 5340
rect 7420 5300 7450 5340
rect 7350 5270 7450 5300
rect 8330 5340 8430 5370
rect 8330 5300 8360 5340
rect 8400 5300 8430 5340
rect 8330 5270 8430 5300
rect 9630 5340 9730 5370
rect 9630 5300 9660 5340
rect 9700 5300 9730 5340
rect 9630 5270 9730 5300
rect 10610 5340 10710 5370
rect 10610 5300 10640 5340
rect 10680 5300 10710 5340
rect 10610 5270 10710 5300
rect 810 3810 890 3840
rect 810 3770 830 3810
rect 870 3770 890 3810
rect 810 3730 890 3770
rect 810 3690 830 3730
rect 870 3690 890 3730
rect 810 3650 890 3690
rect 810 3610 830 3650
rect 870 3610 890 3650
rect 810 3580 890 3610
rect 1690 3810 1770 3840
rect 1690 3770 1710 3810
rect 1750 3770 1770 3810
rect 1690 3730 1770 3770
rect 1690 3690 1710 3730
rect 1750 3690 1770 3730
rect 1690 3650 1770 3690
rect 1690 3610 1710 3650
rect 1750 3610 1770 3650
rect 1690 3580 1770 3610
rect -90 3130 -10 3160
rect -90 3090 -70 3130
rect -30 3090 -10 3130
rect -90 3030 -10 3090
rect -90 2990 -70 3030
rect -30 2990 -10 3030
rect -90 2930 -10 2990
rect -90 2890 -70 2930
rect -30 2890 -10 2930
rect -90 2830 -10 2890
rect -90 2790 -70 2830
rect -30 2790 -10 2830
rect -90 2730 -10 2790
rect -90 2690 -70 2730
rect -30 2690 -10 2730
rect -90 2660 -10 2690
rect 2590 3130 2670 3160
rect 2590 3090 2610 3130
rect 2650 3090 2670 3130
rect 2590 3030 2670 3090
rect 2590 2990 2610 3030
rect 2650 2990 2670 3030
rect 2590 2930 2670 2990
rect 2590 2890 2610 2930
rect 2650 2890 2670 2930
rect 2590 2830 2670 2890
rect 2590 2790 2610 2830
rect 2650 2790 2670 2830
rect 2590 2730 2670 2790
rect 2590 2690 2610 2730
rect 2650 2690 2670 2730
rect 2590 2670 2670 2690
rect 3410 2220 3490 2250
rect 3410 2180 3430 2220
rect 3470 2180 3490 2220
rect 3410 2120 3490 2180
rect 3410 2080 3430 2120
rect 3470 2080 3490 2120
rect 3410 2050 3490 2080
rect -714 1519 574 1554
rect -714 1496 -580 1519
rect -714 1462 -681 1496
rect -647 1485 -580 1496
rect -546 1485 -490 1519
rect -456 1485 -400 1519
rect -366 1485 -310 1519
rect -276 1485 -220 1519
rect -186 1485 -130 1519
rect -96 1485 -40 1519
rect -6 1485 50 1519
rect 84 1485 140 1519
rect 174 1485 230 1519
rect 264 1485 320 1519
rect 354 1485 410 1519
rect 444 1496 574 1519
rect 444 1485 506 1496
rect -647 1462 506 1485
rect 540 1462 574 1496
rect -714 1453 574 1462
rect -714 1406 -613 1453
rect -714 1372 -681 1406
rect -647 1372 -613 1406
rect 473 1406 574 1453
rect -714 1316 -613 1372
rect -714 1282 -681 1316
rect -647 1282 -613 1316
rect -714 1226 -613 1282
rect -714 1192 -681 1226
rect -647 1192 -613 1226
rect -714 1136 -613 1192
rect -714 1102 -681 1136
rect -647 1102 -613 1136
rect -714 1046 -613 1102
rect -714 1012 -681 1046
rect -647 1012 -613 1046
rect -714 956 -613 1012
rect -714 922 -681 956
rect -647 922 -613 956
rect -714 866 -613 922
rect -714 832 -681 866
rect -647 832 -613 866
rect -714 776 -613 832
rect -714 742 -681 776
rect -647 742 -613 776
rect -714 686 -613 742
rect -714 652 -681 686
rect -647 652 -613 686
rect -714 596 -613 652
rect -714 562 -681 596
rect -647 562 -613 596
rect -714 506 -613 562
rect -714 472 -681 506
rect -647 472 -613 506
rect -714 416 -613 472
rect 473 1372 506 1406
rect 540 1372 574 1406
rect 473 1316 574 1372
rect 473 1282 506 1316
rect 540 1282 574 1316
rect 473 1226 574 1282
rect 473 1192 506 1226
rect 540 1192 574 1226
rect 473 1136 574 1192
rect 473 1102 506 1136
rect 540 1102 574 1136
rect 473 1046 574 1102
rect 473 1012 506 1046
rect 540 1012 574 1046
rect 473 956 574 1012
rect 473 922 506 956
rect 540 922 574 956
rect 473 866 574 922
rect 473 832 506 866
rect 540 832 574 866
rect 473 776 574 832
rect 473 742 506 776
rect 540 742 574 776
rect 473 686 574 742
rect 473 652 506 686
rect 540 652 574 686
rect 473 596 574 652
rect 473 562 506 596
rect 540 562 574 596
rect 473 506 574 562
rect 473 472 506 506
rect 540 472 574 506
rect -714 382 -681 416
rect -647 382 -613 416
rect -714 367 -613 382
rect 473 416 574 472
rect 473 382 506 416
rect 540 382 574 416
rect 473 367 574 382
rect -714 332 574 367
rect -714 298 -580 332
rect -546 298 -490 332
rect -456 298 -400 332
rect -366 298 -310 332
rect -276 298 -220 332
rect -186 298 -130 332
rect -96 298 -40 332
rect -6 298 50 332
rect 84 298 140 332
rect 174 298 230 332
rect 264 298 320 332
rect 354 298 410 332
rect 444 298 574 332
rect -714 266 574 298
rect 646 1519 1934 1554
rect 646 1496 780 1519
rect 646 1462 679 1496
rect 713 1485 780 1496
rect 814 1485 870 1519
rect 904 1485 960 1519
rect 994 1485 1050 1519
rect 1084 1485 1140 1519
rect 1174 1485 1230 1519
rect 1264 1485 1320 1519
rect 1354 1485 1410 1519
rect 1444 1485 1500 1519
rect 1534 1485 1590 1519
rect 1624 1485 1680 1519
rect 1714 1485 1770 1519
rect 1804 1496 1934 1519
rect 1804 1485 1866 1496
rect 713 1462 1866 1485
rect 1900 1462 1934 1496
rect 646 1453 1934 1462
rect 646 1406 747 1453
rect 646 1372 679 1406
rect 713 1372 747 1406
rect 1833 1406 1934 1453
rect 646 1316 747 1372
rect 646 1282 679 1316
rect 713 1282 747 1316
rect 646 1226 747 1282
rect 646 1192 679 1226
rect 713 1192 747 1226
rect 646 1136 747 1192
rect 646 1102 679 1136
rect 713 1102 747 1136
rect 646 1046 747 1102
rect 646 1012 679 1046
rect 713 1012 747 1046
rect 646 956 747 1012
rect 646 922 679 956
rect 713 922 747 956
rect 646 866 747 922
rect 646 832 679 866
rect 713 832 747 866
rect 646 776 747 832
rect 646 742 679 776
rect 713 742 747 776
rect 646 686 747 742
rect 646 652 679 686
rect 713 652 747 686
rect 646 596 747 652
rect 646 562 679 596
rect 713 562 747 596
rect 646 506 747 562
rect 646 472 679 506
rect 713 472 747 506
rect 646 416 747 472
rect 1833 1372 1866 1406
rect 1900 1372 1934 1406
rect 1833 1316 1934 1372
rect 1833 1282 1866 1316
rect 1900 1282 1934 1316
rect 1833 1226 1934 1282
rect 1833 1192 1866 1226
rect 1900 1192 1934 1226
rect 1833 1136 1934 1192
rect 1833 1102 1866 1136
rect 1900 1102 1934 1136
rect 1833 1046 1934 1102
rect 1833 1012 1866 1046
rect 1900 1012 1934 1046
rect 1833 956 1934 1012
rect 1833 922 1866 956
rect 1900 922 1934 956
rect 1833 866 1934 922
rect 1833 832 1866 866
rect 1900 832 1934 866
rect 1833 776 1934 832
rect 1833 742 1866 776
rect 1900 742 1934 776
rect 1833 686 1934 742
rect 1833 652 1866 686
rect 1900 652 1934 686
rect 1833 596 1934 652
rect 1833 562 1866 596
rect 1900 562 1934 596
rect 1833 506 1934 562
rect 1833 472 1866 506
rect 1900 472 1934 506
rect 646 382 679 416
rect 713 382 747 416
rect 646 367 747 382
rect 1833 416 1934 472
rect 1833 382 1866 416
rect 1900 382 1934 416
rect 1833 367 1934 382
rect 646 332 1934 367
rect 646 298 780 332
rect 814 298 870 332
rect 904 298 960 332
rect 994 298 1050 332
rect 1084 298 1140 332
rect 1174 298 1230 332
rect 1264 298 1320 332
rect 1354 298 1410 332
rect 1444 298 1500 332
rect 1534 298 1590 332
rect 1624 298 1680 332
rect 1714 298 1770 332
rect 1804 298 1934 332
rect 646 266 1934 298
rect 2006 1519 3294 1554
rect 2006 1496 2140 1519
rect 2006 1462 2039 1496
rect 2073 1485 2140 1496
rect 2174 1485 2230 1519
rect 2264 1485 2320 1519
rect 2354 1485 2410 1519
rect 2444 1485 2500 1519
rect 2534 1485 2590 1519
rect 2624 1485 2680 1519
rect 2714 1485 2770 1519
rect 2804 1485 2860 1519
rect 2894 1485 2950 1519
rect 2984 1485 3040 1519
rect 3074 1485 3130 1519
rect 3164 1496 3294 1519
rect 3164 1485 3226 1496
rect 2073 1462 3226 1485
rect 3260 1462 3294 1496
rect 2006 1453 3294 1462
rect 2006 1406 2107 1453
rect 2006 1372 2039 1406
rect 2073 1372 2107 1406
rect 3193 1406 3294 1453
rect 2006 1316 2107 1372
rect 2006 1282 2039 1316
rect 2073 1282 2107 1316
rect 2006 1226 2107 1282
rect 2006 1192 2039 1226
rect 2073 1192 2107 1226
rect 2006 1136 2107 1192
rect 2006 1102 2039 1136
rect 2073 1102 2107 1136
rect 2006 1046 2107 1102
rect 2006 1012 2039 1046
rect 2073 1012 2107 1046
rect 2006 956 2107 1012
rect 2006 922 2039 956
rect 2073 922 2107 956
rect 2006 866 2107 922
rect 2006 832 2039 866
rect 2073 832 2107 866
rect 2006 776 2107 832
rect 2006 742 2039 776
rect 2073 742 2107 776
rect 2006 686 2107 742
rect 2006 652 2039 686
rect 2073 652 2107 686
rect 2006 596 2107 652
rect 2006 562 2039 596
rect 2073 562 2107 596
rect 2006 506 2107 562
rect 2006 472 2039 506
rect 2073 472 2107 506
rect 2006 416 2107 472
rect 3193 1372 3226 1406
rect 3260 1372 3294 1406
rect 3193 1316 3294 1372
rect 3193 1282 3226 1316
rect 3260 1282 3294 1316
rect 3193 1226 3294 1282
rect 3193 1192 3226 1226
rect 3260 1192 3294 1226
rect 3193 1136 3294 1192
rect 3193 1102 3226 1136
rect 3260 1102 3294 1136
rect 3193 1046 3294 1102
rect 3193 1012 3226 1046
rect 3260 1012 3294 1046
rect 3193 956 3294 1012
rect 3193 922 3226 956
rect 3260 922 3294 956
rect 3193 866 3294 922
rect 3193 832 3226 866
rect 3260 832 3294 866
rect 3193 776 3294 832
rect 3193 742 3226 776
rect 3260 742 3294 776
rect 3193 686 3294 742
rect 3193 652 3226 686
rect 3260 652 3294 686
rect 3193 596 3294 652
rect 3193 562 3226 596
rect 3260 562 3294 596
rect 3193 506 3294 562
rect 3193 472 3226 506
rect 3260 472 3294 506
rect 2006 382 2039 416
rect 2073 382 2107 416
rect 2006 367 2107 382
rect 3193 416 3294 472
rect 3193 382 3226 416
rect 3260 382 3294 416
rect 3193 367 3294 382
rect 2006 332 3294 367
rect 2006 298 2140 332
rect 2174 298 2230 332
rect 2264 298 2320 332
rect 2354 298 2410 332
rect 2444 298 2500 332
rect 2534 298 2590 332
rect 2624 298 2680 332
rect 2714 298 2770 332
rect 2804 298 2860 332
rect 2894 298 2950 332
rect 2984 298 3040 332
rect 3074 298 3130 332
rect 3164 298 3294 332
rect 2006 266 3294 298
rect -714 159 574 194
rect -714 136 -580 159
rect -714 102 -681 136
rect -647 125 -580 136
rect -546 125 -490 159
rect -456 125 -400 159
rect -366 125 -310 159
rect -276 125 -220 159
rect -186 125 -130 159
rect -96 125 -40 159
rect -6 125 50 159
rect 84 125 140 159
rect 174 125 230 159
rect 264 125 320 159
rect 354 125 410 159
rect 444 136 574 159
rect 444 125 506 136
rect -647 102 506 125
rect 540 102 574 136
rect -714 93 574 102
rect -714 46 -613 93
rect -714 12 -681 46
rect -647 12 -613 46
rect 473 46 574 93
rect -714 -44 -613 12
rect -714 -78 -681 -44
rect -647 -78 -613 -44
rect -714 -134 -613 -78
rect -714 -168 -681 -134
rect -647 -168 -613 -134
rect -714 -224 -613 -168
rect -714 -258 -681 -224
rect -647 -258 -613 -224
rect -714 -314 -613 -258
rect -714 -348 -681 -314
rect -647 -348 -613 -314
rect -714 -404 -613 -348
rect -714 -438 -681 -404
rect -647 -438 -613 -404
rect -714 -494 -613 -438
rect -714 -528 -681 -494
rect -647 -528 -613 -494
rect -714 -584 -613 -528
rect -714 -618 -681 -584
rect -647 -618 -613 -584
rect -714 -674 -613 -618
rect -714 -708 -681 -674
rect -647 -708 -613 -674
rect -714 -764 -613 -708
rect -714 -798 -681 -764
rect -647 -798 -613 -764
rect -714 -854 -613 -798
rect -714 -888 -681 -854
rect -647 -888 -613 -854
rect -714 -944 -613 -888
rect 473 12 506 46
rect 540 12 574 46
rect 473 -44 574 12
rect 473 -78 506 -44
rect 540 -78 574 -44
rect 473 -134 574 -78
rect 473 -168 506 -134
rect 540 -168 574 -134
rect 473 -224 574 -168
rect 473 -258 506 -224
rect 540 -258 574 -224
rect 473 -314 574 -258
rect 473 -348 506 -314
rect 540 -348 574 -314
rect 473 -404 574 -348
rect 473 -438 506 -404
rect 540 -438 574 -404
rect 473 -494 574 -438
rect 473 -528 506 -494
rect 540 -528 574 -494
rect 473 -584 574 -528
rect 473 -618 506 -584
rect 540 -618 574 -584
rect 473 -674 574 -618
rect 473 -708 506 -674
rect 540 -708 574 -674
rect 473 -764 574 -708
rect 473 -798 506 -764
rect 540 -798 574 -764
rect 473 -854 574 -798
rect 473 -888 506 -854
rect 540 -888 574 -854
rect -714 -978 -681 -944
rect -647 -978 -613 -944
rect -714 -993 -613 -978
rect 473 -944 574 -888
rect 473 -978 506 -944
rect 540 -978 574 -944
rect 473 -993 574 -978
rect -714 -1028 574 -993
rect -714 -1062 -580 -1028
rect -546 -1062 -490 -1028
rect -456 -1062 -400 -1028
rect -366 -1062 -310 -1028
rect -276 -1062 -220 -1028
rect -186 -1062 -130 -1028
rect -96 -1062 -40 -1028
rect -6 -1062 50 -1028
rect 84 -1062 140 -1028
rect 174 -1062 230 -1028
rect 264 -1062 320 -1028
rect 354 -1062 410 -1028
rect 444 -1062 574 -1028
rect -714 -1094 574 -1062
rect 646 159 1934 194
rect 646 136 780 159
rect 646 102 679 136
rect 713 125 780 136
rect 814 125 870 159
rect 904 125 960 159
rect 994 125 1050 159
rect 1084 125 1140 159
rect 1174 125 1230 159
rect 1264 125 1320 159
rect 1354 125 1410 159
rect 1444 125 1500 159
rect 1534 125 1590 159
rect 1624 125 1680 159
rect 1714 125 1770 159
rect 1804 136 1934 159
rect 1804 125 1866 136
rect 713 102 1866 125
rect 1900 102 1934 136
rect 646 93 1934 102
rect 646 46 747 93
rect 646 12 679 46
rect 713 12 747 46
rect 1833 46 1934 93
rect 646 -44 747 12
rect 646 -78 679 -44
rect 713 -78 747 -44
rect 646 -134 747 -78
rect 646 -168 679 -134
rect 713 -168 747 -134
rect 646 -224 747 -168
rect 646 -258 679 -224
rect 713 -258 747 -224
rect 646 -314 747 -258
rect 646 -348 679 -314
rect 713 -348 747 -314
rect 646 -404 747 -348
rect 646 -438 679 -404
rect 713 -438 747 -404
rect 646 -494 747 -438
rect 646 -528 679 -494
rect 713 -528 747 -494
rect 646 -584 747 -528
rect 646 -618 679 -584
rect 713 -618 747 -584
rect 646 -674 747 -618
rect 646 -708 679 -674
rect 713 -708 747 -674
rect 646 -764 747 -708
rect 646 -798 679 -764
rect 713 -798 747 -764
rect 646 -854 747 -798
rect 646 -888 679 -854
rect 713 -888 747 -854
rect 646 -944 747 -888
rect 1833 12 1866 46
rect 1900 12 1934 46
rect 1833 -44 1934 12
rect 1833 -78 1866 -44
rect 1900 -78 1934 -44
rect 1833 -134 1934 -78
rect 1833 -168 1866 -134
rect 1900 -168 1934 -134
rect 1833 -224 1934 -168
rect 1833 -258 1866 -224
rect 1900 -258 1934 -224
rect 1833 -314 1934 -258
rect 1833 -348 1866 -314
rect 1900 -348 1934 -314
rect 1833 -404 1934 -348
rect 1833 -438 1866 -404
rect 1900 -438 1934 -404
rect 1833 -494 1934 -438
rect 1833 -528 1866 -494
rect 1900 -528 1934 -494
rect 1833 -584 1934 -528
rect 1833 -618 1866 -584
rect 1900 -618 1934 -584
rect 1833 -674 1934 -618
rect 1833 -708 1866 -674
rect 1900 -708 1934 -674
rect 1833 -764 1934 -708
rect 1833 -798 1866 -764
rect 1900 -798 1934 -764
rect 1833 -854 1934 -798
rect 1833 -888 1866 -854
rect 1900 -888 1934 -854
rect 646 -978 679 -944
rect 713 -978 747 -944
rect 646 -993 747 -978
rect 1833 -944 1934 -888
rect 1833 -978 1866 -944
rect 1900 -978 1934 -944
rect 1833 -993 1934 -978
rect 646 -1028 1934 -993
rect 646 -1062 780 -1028
rect 814 -1062 870 -1028
rect 904 -1062 960 -1028
rect 994 -1062 1050 -1028
rect 1084 -1062 1140 -1028
rect 1174 -1062 1230 -1028
rect 1264 -1062 1320 -1028
rect 1354 -1062 1410 -1028
rect 1444 -1062 1500 -1028
rect 1534 -1062 1590 -1028
rect 1624 -1062 1680 -1028
rect 1714 -1062 1770 -1028
rect 1804 -1062 1934 -1028
rect 646 -1094 1934 -1062
rect 2006 159 3294 194
rect 2006 136 2140 159
rect 2006 102 2039 136
rect 2073 125 2140 136
rect 2174 125 2230 159
rect 2264 125 2320 159
rect 2354 125 2410 159
rect 2444 125 2500 159
rect 2534 125 2590 159
rect 2624 125 2680 159
rect 2714 125 2770 159
rect 2804 125 2860 159
rect 2894 125 2950 159
rect 2984 125 3040 159
rect 3074 125 3130 159
rect 3164 136 3294 159
rect 3164 125 3226 136
rect 2073 102 3226 125
rect 3260 102 3294 136
rect 2006 93 3294 102
rect 2006 46 2107 93
rect 2006 12 2039 46
rect 2073 12 2107 46
rect 3193 46 3294 93
rect 2006 -44 2107 12
rect 2006 -78 2039 -44
rect 2073 -78 2107 -44
rect 2006 -134 2107 -78
rect 2006 -168 2039 -134
rect 2073 -168 2107 -134
rect 2006 -224 2107 -168
rect 2006 -258 2039 -224
rect 2073 -258 2107 -224
rect 2006 -314 2107 -258
rect 2006 -348 2039 -314
rect 2073 -348 2107 -314
rect 2006 -404 2107 -348
rect 2006 -438 2039 -404
rect 2073 -438 2107 -404
rect 2006 -494 2107 -438
rect 2006 -528 2039 -494
rect 2073 -528 2107 -494
rect 2006 -584 2107 -528
rect 2006 -618 2039 -584
rect 2073 -618 2107 -584
rect 2006 -674 2107 -618
rect 2006 -708 2039 -674
rect 2073 -708 2107 -674
rect 2006 -764 2107 -708
rect 2006 -798 2039 -764
rect 2073 -798 2107 -764
rect 2006 -854 2107 -798
rect 2006 -888 2039 -854
rect 2073 -888 2107 -854
rect 2006 -944 2107 -888
rect 3193 12 3226 46
rect 3260 12 3294 46
rect 3193 -44 3294 12
rect 3193 -78 3226 -44
rect 3260 -78 3294 -44
rect 3193 -134 3294 -78
rect 3193 -168 3226 -134
rect 3260 -168 3294 -134
rect 3193 -224 3294 -168
rect 3193 -258 3226 -224
rect 3260 -258 3294 -224
rect 3193 -314 3294 -258
rect 3193 -348 3226 -314
rect 3260 -348 3294 -314
rect 3193 -404 3294 -348
rect 3193 -438 3226 -404
rect 3260 -438 3294 -404
rect 3193 -494 3294 -438
rect 3193 -528 3226 -494
rect 3260 -528 3294 -494
rect 3193 -584 3294 -528
rect 3193 -618 3226 -584
rect 3260 -618 3294 -584
rect 3193 -674 3294 -618
rect 3193 -708 3226 -674
rect 3260 -708 3294 -674
rect 3193 -764 3294 -708
rect 3193 -798 3226 -764
rect 3260 -798 3294 -764
rect 3193 -854 3294 -798
rect 3193 -888 3226 -854
rect 3260 -888 3294 -854
rect 2006 -978 2039 -944
rect 2073 -978 2107 -944
rect 2006 -993 2107 -978
rect 3193 -944 3294 -888
rect 3193 -978 3226 -944
rect 3260 -978 3294 -944
rect 3193 -993 3294 -978
rect 2006 -1028 3294 -993
rect 2006 -1062 2140 -1028
rect 2174 -1062 2230 -1028
rect 2264 -1062 2320 -1028
rect 2354 -1062 2410 -1028
rect 2444 -1062 2500 -1028
rect 2534 -1062 2590 -1028
rect 2624 -1062 2680 -1028
rect 2714 -1062 2770 -1028
rect 2804 -1062 2860 -1028
rect 2894 -1062 2950 -1028
rect 2984 -1062 3040 -1028
rect 3074 -1062 3130 -1028
rect 3164 -1062 3294 -1028
rect 2006 -1094 3294 -1062
rect -714 -1201 574 -1166
rect -714 -1224 -580 -1201
rect -714 -1258 -681 -1224
rect -647 -1235 -580 -1224
rect -546 -1235 -490 -1201
rect -456 -1235 -400 -1201
rect -366 -1235 -310 -1201
rect -276 -1235 -220 -1201
rect -186 -1235 -130 -1201
rect -96 -1235 -40 -1201
rect -6 -1235 50 -1201
rect 84 -1235 140 -1201
rect 174 -1235 230 -1201
rect 264 -1235 320 -1201
rect 354 -1235 410 -1201
rect 444 -1224 574 -1201
rect 444 -1235 506 -1224
rect -647 -1258 506 -1235
rect 540 -1258 574 -1224
rect -714 -1267 574 -1258
rect -714 -1314 -613 -1267
rect -714 -1348 -681 -1314
rect -647 -1348 -613 -1314
rect 473 -1314 574 -1267
rect -714 -1404 -613 -1348
rect -714 -1438 -681 -1404
rect -647 -1438 -613 -1404
rect -714 -1494 -613 -1438
rect -714 -1528 -681 -1494
rect -647 -1528 -613 -1494
rect -714 -1584 -613 -1528
rect -714 -1618 -681 -1584
rect -647 -1618 -613 -1584
rect -714 -1674 -613 -1618
rect -714 -1708 -681 -1674
rect -647 -1708 -613 -1674
rect -714 -1764 -613 -1708
rect -714 -1798 -681 -1764
rect -647 -1798 -613 -1764
rect -714 -1854 -613 -1798
rect -714 -1888 -681 -1854
rect -647 -1888 -613 -1854
rect -714 -1944 -613 -1888
rect -714 -1978 -681 -1944
rect -647 -1978 -613 -1944
rect -714 -2034 -613 -1978
rect -714 -2068 -681 -2034
rect -647 -2068 -613 -2034
rect -714 -2124 -613 -2068
rect -714 -2158 -681 -2124
rect -647 -2158 -613 -2124
rect -714 -2214 -613 -2158
rect -714 -2248 -681 -2214
rect -647 -2248 -613 -2214
rect -714 -2304 -613 -2248
rect 473 -1348 506 -1314
rect 540 -1348 574 -1314
rect 473 -1404 574 -1348
rect 473 -1438 506 -1404
rect 540 -1438 574 -1404
rect 473 -1494 574 -1438
rect 473 -1528 506 -1494
rect 540 -1528 574 -1494
rect 473 -1584 574 -1528
rect 473 -1618 506 -1584
rect 540 -1618 574 -1584
rect 473 -1674 574 -1618
rect 473 -1708 506 -1674
rect 540 -1708 574 -1674
rect 473 -1764 574 -1708
rect 473 -1798 506 -1764
rect 540 -1798 574 -1764
rect 473 -1854 574 -1798
rect 473 -1888 506 -1854
rect 540 -1888 574 -1854
rect 473 -1944 574 -1888
rect 473 -1978 506 -1944
rect 540 -1978 574 -1944
rect 473 -2034 574 -1978
rect 473 -2068 506 -2034
rect 540 -2068 574 -2034
rect 473 -2124 574 -2068
rect 473 -2158 506 -2124
rect 540 -2158 574 -2124
rect 473 -2214 574 -2158
rect 473 -2248 506 -2214
rect 540 -2248 574 -2214
rect -714 -2338 -681 -2304
rect -647 -2338 -613 -2304
rect -714 -2353 -613 -2338
rect 473 -2304 574 -2248
rect 473 -2338 506 -2304
rect 540 -2338 574 -2304
rect 473 -2353 574 -2338
rect -714 -2388 574 -2353
rect -714 -2422 -580 -2388
rect -546 -2422 -490 -2388
rect -456 -2422 -400 -2388
rect -366 -2422 -310 -2388
rect -276 -2422 -220 -2388
rect -186 -2422 -130 -2388
rect -96 -2422 -40 -2388
rect -6 -2422 50 -2388
rect 84 -2422 140 -2388
rect 174 -2422 230 -2388
rect 264 -2422 320 -2388
rect 354 -2422 410 -2388
rect 444 -2422 574 -2388
rect -714 -2454 574 -2422
rect 646 -1201 1934 -1166
rect 646 -1224 780 -1201
rect 646 -1258 679 -1224
rect 713 -1235 780 -1224
rect 814 -1235 870 -1201
rect 904 -1235 960 -1201
rect 994 -1235 1050 -1201
rect 1084 -1235 1140 -1201
rect 1174 -1235 1230 -1201
rect 1264 -1235 1320 -1201
rect 1354 -1235 1410 -1201
rect 1444 -1235 1500 -1201
rect 1534 -1235 1590 -1201
rect 1624 -1235 1680 -1201
rect 1714 -1235 1770 -1201
rect 1804 -1224 1934 -1201
rect 1804 -1235 1866 -1224
rect 713 -1258 1866 -1235
rect 1900 -1258 1934 -1224
rect 646 -1267 1934 -1258
rect 646 -1314 747 -1267
rect 646 -1348 679 -1314
rect 713 -1348 747 -1314
rect 1833 -1314 1934 -1267
rect 646 -1404 747 -1348
rect 646 -1438 679 -1404
rect 713 -1438 747 -1404
rect 646 -1494 747 -1438
rect 646 -1528 679 -1494
rect 713 -1528 747 -1494
rect 646 -1584 747 -1528
rect 646 -1618 679 -1584
rect 713 -1618 747 -1584
rect 646 -1674 747 -1618
rect 646 -1708 679 -1674
rect 713 -1708 747 -1674
rect 646 -1764 747 -1708
rect 646 -1798 679 -1764
rect 713 -1798 747 -1764
rect 646 -1854 747 -1798
rect 646 -1888 679 -1854
rect 713 -1888 747 -1854
rect 646 -1944 747 -1888
rect 646 -1978 679 -1944
rect 713 -1978 747 -1944
rect 646 -2034 747 -1978
rect 646 -2068 679 -2034
rect 713 -2068 747 -2034
rect 646 -2124 747 -2068
rect 646 -2158 679 -2124
rect 713 -2158 747 -2124
rect 646 -2214 747 -2158
rect 646 -2248 679 -2214
rect 713 -2248 747 -2214
rect 646 -2304 747 -2248
rect 1833 -1348 1866 -1314
rect 1900 -1348 1934 -1314
rect 1833 -1404 1934 -1348
rect 1833 -1438 1866 -1404
rect 1900 -1438 1934 -1404
rect 1833 -1494 1934 -1438
rect 1833 -1528 1866 -1494
rect 1900 -1528 1934 -1494
rect 1833 -1584 1934 -1528
rect 1833 -1618 1866 -1584
rect 1900 -1618 1934 -1584
rect 1833 -1674 1934 -1618
rect 1833 -1708 1866 -1674
rect 1900 -1708 1934 -1674
rect 1833 -1764 1934 -1708
rect 1833 -1798 1866 -1764
rect 1900 -1798 1934 -1764
rect 1833 -1854 1934 -1798
rect 1833 -1888 1866 -1854
rect 1900 -1888 1934 -1854
rect 1833 -1944 1934 -1888
rect 1833 -1978 1866 -1944
rect 1900 -1978 1934 -1944
rect 1833 -2034 1934 -1978
rect 1833 -2068 1866 -2034
rect 1900 -2068 1934 -2034
rect 1833 -2124 1934 -2068
rect 1833 -2158 1866 -2124
rect 1900 -2158 1934 -2124
rect 1833 -2214 1934 -2158
rect 1833 -2248 1866 -2214
rect 1900 -2248 1934 -2214
rect 646 -2338 679 -2304
rect 713 -2338 747 -2304
rect 646 -2353 747 -2338
rect 1833 -2304 1934 -2248
rect 1833 -2338 1866 -2304
rect 1900 -2338 1934 -2304
rect 1833 -2353 1934 -2338
rect 646 -2388 1934 -2353
rect 646 -2422 780 -2388
rect 814 -2422 870 -2388
rect 904 -2422 960 -2388
rect 994 -2422 1050 -2388
rect 1084 -2422 1140 -2388
rect 1174 -2422 1230 -2388
rect 1264 -2422 1320 -2388
rect 1354 -2422 1410 -2388
rect 1444 -2422 1500 -2388
rect 1534 -2422 1590 -2388
rect 1624 -2422 1680 -2388
rect 1714 -2422 1770 -2388
rect 1804 -2422 1934 -2388
rect 646 -2454 1934 -2422
rect 2006 -1201 3294 -1166
rect 2006 -1224 2140 -1201
rect 2006 -1258 2039 -1224
rect 2073 -1235 2140 -1224
rect 2174 -1235 2230 -1201
rect 2264 -1235 2320 -1201
rect 2354 -1235 2410 -1201
rect 2444 -1235 2500 -1201
rect 2534 -1235 2590 -1201
rect 2624 -1235 2680 -1201
rect 2714 -1235 2770 -1201
rect 2804 -1235 2860 -1201
rect 2894 -1235 2950 -1201
rect 2984 -1235 3040 -1201
rect 3074 -1235 3130 -1201
rect 3164 -1224 3294 -1201
rect 3164 -1235 3226 -1224
rect 2073 -1258 3226 -1235
rect 3260 -1258 3294 -1224
rect 2006 -1267 3294 -1258
rect 2006 -1314 2107 -1267
rect 2006 -1348 2039 -1314
rect 2073 -1348 2107 -1314
rect 3193 -1314 3294 -1267
rect 2006 -1404 2107 -1348
rect 2006 -1438 2039 -1404
rect 2073 -1438 2107 -1404
rect 2006 -1494 2107 -1438
rect 2006 -1528 2039 -1494
rect 2073 -1528 2107 -1494
rect 2006 -1584 2107 -1528
rect 2006 -1618 2039 -1584
rect 2073 -1618 2107 -1584
rect 2006 -1674 2107 -1618
rect 2006 -1708 2039 -1674
rect 2073 -1708 2107 -1674
rect 2006 -1764 2107 -1708
rect 2006 -1798 2039 -1764
rect 2073 -1798 2107 -1764
rect 2006 -1854 2107 -1798
rect 2006 -1888 2039 -1854
rect 2073 -1888 2107 -1854
rect 2006 -1944 2107 -1888
rect 2006 -1978 2039 -1944
rect 2073 -1978 2107 -1944
rect 2006 -2034 2107 -1978
rect 2006 -2068 2039 -2034
rect 2073 -2068 2107 -2034
rect 2006 -2124 2107 -2068
rect 2006 -2158 2039 -2124
rect 2073 -2158 2107 -2124
rect 2006 -2214 2107 -2158
rect 2006 -2248 2039 -2214
rect 2073 -2248 2107 -2214
rect 2006 -2304 2107 -2248
rect 3193 -1348 3226 -1314
rect 3260 -1348 3294 -1314
rect 3193 -1404 3294 -1348
rect 3193 -1438 3226 -1404
rect 3260 -1438 3294 -1404
rect 3193 -1494 3294 -1438
rect 3193 -1528 3226 -1494
rect 3260 -1528 3294 -1494
rect 3193 -1584 3294 -1528
rect 3193 -1618 3226 -1584
rect 3260 -1618 3294 -1584
rect 3193 -1674 3294 -1618
rect 3193 -1708 3226 -1674
rect 3260 -1708 3294 -1674
rect 3193 -1764 3294 -1708
rect 3193 -1798 3226 -1764
rect 3260 -1798 3294 -1764
rect 3193 -1854 3294 -1798
rect 3193 -1888 3226 -1854
rect 3260 -1888 3294 -1854
rect 3193 -1944 3294 -1888
rect 3193 -1978 3226 -1944
rect 3260 -1978 3294 -1944
rect 3193 -2034 3294 -1978
rect 3193 -2068 3226 -2034
rect 3260 -2068 3294 -2034
rect 3193 -2124 3294 -2068
rect 3193 -2158 3226 -2124
rect 3260 -2158 3294 -2124
rect 3193 -2214 3294 -2158
rect 3193 -2248 3226 -2214
rect 3260 -2248 3294 -2214
rect 2006 -2338 2039 -2304
rect 2073 -2338 2107 -2304
rect 2006 -2353 2107 -2338
rect 3193 -2304 3294 -2248
rect 3193 -2338 3226 -2304
rect 3260 -2338 3294 -2304
rect 3193 -2353 3294 -2338
rect 2006 -2388 3294 -2353
rect 2006 -2422 2140 -2388
rect 2174 -2422 2230 -2388
rect 2264 -2422 2320 -2388
rect 2354 -2422 2410 -2388
rect 2444 -2422 2500 -2388
rect 2534 -2422 2590 -2388
rect 2624 -2422 2680 -2388
rect 2714 -2422 2770 -2388
rect 2804 -2422 2860 -2388
rect 2894 -2422 2950 -2388
rect 2984 -2422 3040 -2388
rect 3074 -2422 3130 -2388
rect 3164 -2422 3294 -2388
rect 2006 -2454 3294 -2422
rect 1240 -2540 1340 -2510
rect 1240 -2580 1270 -2540
rect 1310 -2580 1340 -2540
rect 1240 -2620 1340 -2580
rect 1240 -2660 1270 -2620
rect 1310 -2660 1340 -2620
rect 1240 -2700 1340 -2660
rect 1240 -2740 1270 -2700
rect 1310 -2740 1340 -2700
rect 1240 -2770 1340 -2740
<< nsubdiff >>
rect 790 12870 870 12900
rect 790 12830 810 12870
rect 850 12830 870 12870
rect 790 12800 870 12830
rect 3160 12870 3240 12900
rect 3160 12830 3180 12870
rect 3220 12830 3240 12870
rect 3160 12800 3240 12830
rect 11100 12910 12120 12950
rect 12280 12910 13330 12950
rect 6030 12870 6110 12900
rect 6030 12830 6050 12870
rect 6090 12830 6110 12870
rect 6030 12800 6110 12830
rect 7330 12870 7410 12900
rect 7330 12830 7350 12870
rect 7390 12830 7410 12870
rect 7330 12800 7410 12830
rect 8630 12870 8710 12900
rect 8630 12830 8650 12870
rect 8690 12830 8710 12870
rect 8630 12800 8710 12830
rect 9930 12870 10010 12900
rect 9930 12830 9950 12870
rect 9990 12830 10010 12870
rect 9930 12800 10010 12830
rect 11100 11600 11140 12910
rect 13290 11600 13330 12910
rect 11100 10840 11140 11270
rect 13290 10840 13330 11270
rect 11100 10800 12120 10840
rect 12280 10800 13160 10840
rect 13230 10800 13330 10840
rect 1180 9790 1260 9820
rect 1180 9750 1200 9790
rect 1240 9750 1260 9790
rect 1180 9690 1260 9750
rect 1180 9650 1200 9690
rect 1240 9650 1260 9690
rect 1180 9590 1260 9650
rect 1180 9550 1200 9590
rect 1240 9550 1260 9590
rect 1180 9490 1260 9550
rect 1180 9450 1200 9490
rect 1240 9450 1260 9490
rect 1180 9420 1260 9450
rect 2080 9790 2160 9820
rect 2080 9750 2100 9790
rect 2140 9750 2160 9790
rect 2080 9690 2160 9750
rect 2080 9650 2100 9690
rect 2140 9650 2160 9690
rect 2080 9590 2160 9650
rect 2080 9550 2100 9590
rect 2140 9550 2160 9590
rect 2080 9490 2160 9550
rect 2080 9450 2100 9490
rect 2140 9450 2160 9490
rect 2080 9420 2160 9450
rect 2980 9790 3060 9820
rect 2980 9750 3000 9790
rect 3040 9750 3060 9790
rect 2980 9690 3060 9750
rect 2980 9650 3000 9690
rect 3040 9650 3060 9690
rect 2980 9590 3060 9650
rect 2980 9550 3000 9590
rect 3040 9550 3060 9590
rect 2980 9490 3060 9550
rect 2980 9450 3000 9490
rect 3040 9450 3060 9490
rect 2980 9420 3060 9450
rect 3120 9790 3200 9820
rect 3120 9750 3140 9790
rect 3180 9750 3200 9790
rect 3120 9690 3200 9750
rect 3120 9650 3140 9690
rect 3180 9650 3200 9690
rect 3120 9590 3200 9650
rect 3120 9550 3140 9590
rect 3180 9550 3200 9590
rect 3120 9490 3200 9550
rect 3120 9450 3140 9490
rect 3180 9450 3200 9490
rect 3120 9430 3200 9450
rect 3120 9420 3180 9430
rect 3560 9790 3640 9820
rect 3560 9750 3580 9790
rect 3620 9750 3640 9790
rect 3560 9690 3640 9750
rect 3560 9650 3580 9690
rect 3620 9650 3640 9690
rect 3560 9590 3640 9650
rect 3560 9550 3580 9590
rect 3620 9550 3640 9590
rect 3560 9490 3640 9550
rect 3560 9450 3580 9490
rect 3620 9450 3640 9490
rect 3560 9420 3640 9450
rect 3890 9790 3970 9820
rect 3890 9750 3910 9790
rect 3950 9750 3970 9790
rect 3890 9690 3970 9750
rect 3890 9650 3910 9690
rect 3950 9650 3970 9690
rect 3890 9590 3970 9650
rect 3890 9550 3910 9590
rect 3950 9550 3970 9590
rect 3890 9490 3970 9550
rect 3890 9450 3910 9490
rect 3950 9450 3970 9490
rect 3890 9420 3970 9450
rect 4290 9790 4390 9820
rect 4290 9750 4320 9790
rect 4360 9750 4390 9790
rect 4290 9690 4390 9750
rect 4290 9650 4320 9690
rect 4360 9650 4390 9690
rect 4290 9590 4390 9650
rect 4290 9550 4320 9590
rect 4360 9550 4390 9590
rect 4290 9490 4390 9550
rect 4290 9450 4320 9490
rect 4360 9450 4390 9490
rect 4290 9420 4390 9450
rect 4680 9790 4780 9820
rect 4680 9750 4710 9790
rect 4750 9750 4780 9790
rect 4680 9690 4780 9750
rect 4680 9650 4710 9690
rect 4750 9650 4780 9690
rect 4680 9590 4780 9650
rect 4680 9550 4710 9590
rect 4750 9550 4780 9590
rect 4680 9490 4780 9550
rect 4680 9450 4710 9490
rect 4750 9450 4780 9490
rect 4680 9420 4780 9450
rect 5070 9790 5170 9820
rect 5070 9750 5100 9790
rect 5140 9750 5170 9790
rect 5070 9690 5170 9750
rect 5070 9650 5100 9690
rect 5140 9650 5170 9690
rect 5070 9590 5170 9650
rect 5070 9550 5100 9590
rect 5140 9550 5170 9590
rect 5070 9490 5170 9550
rect 5070 9450 5100 9490
rect 5140 9450 5170 9490
rect 5070 9420 5170 9450
rect 5750 9790 5850 9820
rect 5750 9750 5780 9790
rect 5820 9750 5850 9790
rect 5750 9690 5850 9750
rect 5750 9650 5780 9690
rect 5820 9650 5850 9690
rect 5750 9590 5850 9650
rect 5750 9550 5780 9590
rect 5820 9550 5850 9590
rect 5750 9490 5850 9550
rect 5750 9450 5780 9490
rect 5820 9450 5850 9490
rect 5750 9420 5850 9450
rect 7440 9760 7540 9790
rect 7440 9720 7470 9760
rect 7510 9720 7540 9760
rect 7440 9660 7540 9720
rect 7440 9620 7470 9660
rect 7510 9620 7540 9660
rect 7440 9560 7540 9620
rect 7440 9520 7470 9560
rect 7510 9520 7540 9560
rect 7440 9460 7540 9520
rect 7440 9420 7470 9460
rect 7510 9420 7540 9460
rect 7440 9390 7540 9420
rect 8960 9760 9060 9790
rect 8960 9720 8990 9760
rect 9030 9720 9060 9760
rect 8960 9660 9060 9720
rect 8960 9620 8990 9660
rect 9030 9620 9060 9660
rect 8960 9560 9060 9620
rect 8960 9520 8990 9560
rect 9030 9520 9060 9560
rect 8960 9460 9060 9520
rect 8960 9420 8990 9460
rect 9030 9420 9060 9460
rect 8960 9390 9060 9420
rect 10480 9760 10580 9790
rect 10480 9720 10510 9760
rect 10550 9720 10580 9760
rect 10480 9660 10580 9720
rect 10480 9620 10510 9660
rect 10550 9620 10580 9660
rect 10480 9560 10580 9620
rect 10480 9520 10510 9560
rect 10550 9520 10580 9560
rect 10480 9460 10580 9520
rect 10480 9420 10510 9460
rect 10550 9420 10580 9460
rect 10480 9390 10580 9420
rect 1180 9030 1260 9060
rect 1180 8990 1200 9030
rect 1240 8990 1260 9030
rect 1180 8930 1260 8990
rect 1180 8890 1200 8930
rect 1240 8890 1260 8930
rect 1180 8830 1260 8890
rect 1180 8790 1200 8830
rect 1240 8790 1260 8830
rect 1180 8730 1260 8790
rect 1180 8690 1200 8730
rect 1240 8690 1260 8730
rect 1180 8660 1260 8690
rect 2080 9030 2160 9060
rect 2080 8990 2100 9030
rect 2140 8990 2160 9030
rect 2080 8930 2160 8990
rect 2080 8890 2100 8930
rect 2140 8890 2160 8930
rect 2080 8830 2160 8890
rect 2080 8790 2100 8830
rect 2140 8790 2160 8830
rect 2080 8730 2160 8790
rect 2080 8690 2100 8730
rect 2140 8690 2160 8730
rect 2080 8660 2160 8690
rect 2980 9030 3060 9060
rect 2980 8990 3000 9030
rect 3040 8990 3060 9030
rect 2980 8930 3060 8990
rect 2980 8890 3000 8930
rect 3040 8890 3060 8930
rect 2980 8830 3060 8890
rect 2980 8790 3000 8830
rect 3040 8790 3060 8830
rect 2980 8730 3060 8790
rect 2980 8690 3000 8730
rect 3040 8690 3060 8730
rect 2980 8660 3060 8690
rect 3380 9030 3460 9060
rect 3380 8990 3400 9030
rect 3440 8990 3460 9030
rect 3380 8930 3460 8990
rect 3380 8890 3400 8930
rect 3440 8890 3460 8930
rect 3380 8830 3460 8890
rect 3380 8790 3400 8830
rect 3440 8790 3460 8830
rect 3380 8730 3460 8790
rect 3380 8690 3400 8730
rect 3440 8690 3460 8730
rect 3380 8660 3460 8690
rect 3710 9030 3790 9060
rect 3710 8990 3730 9030
rect 3770 8990 3790 9030
rect 3710 8930 3790 8990
rect 3710 8890 3730 8930
rect 3770 8890 3790 8930
rect 3710 8830 3790 8890
rect 3710 8790 3730 8830
rect 3770 8790 3790 8830
rect 3710 8730 3790 8790
rect 3710 8690 3730 8730
rect 3770 8690 3790 8730
rect 3710 8660 3790 8690
rect 4040 9030 4120 9060
rect 4040 8990 4060 9030
rect 4100 8990 4120 9030
rect 4040 8930 4120 8990
rect 4040 8890 4060 8930
rect 4100 8890 4120 8930
rect 4040 8830 4120 8890
rect 4040 8790 4060 8830
rect 4100 8790 4120 8830
rect 4040 8730 4120 8790
rect 4040 8690 4060 8730
rect 4100 8690 4120 8730
rect 4040 8660 4120 8690
rect 4290 9030 4390 9060
rect 4290 8990 4320 9030
rect 4360 8990 4390 9030
rect 4290 8930 4390 8990
rect 4290 8890 4320 8930
rect 4360 8890 4390 8930
rect 4290 8830 4390 8890
rect 4290 8790 4320 8830
rect 4360 8790 4390 8830
rect 4290 8730 4390 8790
rect 4290 8690 4320 8730
rect 4360 8690 4390 8730
rect 4290 8660 4390 8690
rect 5070 9030 5170 9060
rect 5070 8990 5100 9030
rect 5140 8990 5170 9030
rect 5070 8930 5170 8990
rect 5070 8890 5100 8930
rect 5140 8890 5170 8930
rect 5070 8830 5170 8890
rect 5070 8790 5100 8830
rect 5140 8790 5170 8830
rect 5070 8730 5170 8790
rect 5070 8690 5100 8730
rect 5140 8690 5170 8730
rect 5070 8660 5170 8690
rect -440 6840 -360 6870
rect -440 6800 -420 6840
rect -380 6800 -360 6840
rect -440 6740 -360 6800
rect -440 6700 -420 6740
rect -380 6700 -360 6740
rect -440 6670 -360 6700
rect 1040 6840 1120 6870
rect 1040 6800 1060 6840
rect 1100 6800 1120 6840
rect 1040 6740 1120 6800
rect 1040 6700 1060 6740
rect 1100 6700 1120 6740
rect 1040 6670 1120 6700
rect 1460 6840 1540 6870
rect 1460 6800 1480 6840
rect 1520 6800 1540 6840
rect 1460 6740 1540 6800
rect 1460 6700 1480 6740
rect 1520 6700 1540 6740
rect 1460 6670 1540 6700
rect 2940 6840 3020 6870
rect 2940 6800 2960 6840
rect 3000 6800 3020 6840
rect 2940 6740 3020 6800
rect 2940 6700 2960 6740
rect 3000 6700 3020 6740
rect 2940 6670 3020 6700
rect 11043 6811 11139 6845
rect 11399 6811 11495 6845
rect 11043 6749 11077 6811
rect -450 6240 -370 6270
rect -450 6200 -430 6240
rect -390 6200 -370 6240
rect -450 6140 -370 6200
rect -450 6100 -430 6140
rect -390 6100 -370 6140
rect -450 6040 -370 6100
rect -450 6000 -430 6040
rect -390 6000 -370 6040
rect -450 5940 -370 6000
rect -450 5900 -430 5940
rect -390 5900 -370 5940
rect -450 5840 -370 5900
rect -450 5800 -430 5840
rect -390 5800 -370 5840
rect -450 5740 -370 5800
rect -450 5700 -430 5740
rect -390 5700 -370 5740
rect -450 5670 -370 5700
rect 2950 6240 3030 6270
rect 2950 6200 2970 6240
rect 3010 6200 3030 6240
rect 2950 6140 3030 6200
rect 2950 6100 2970 6140
rect 3010 6100 3030 6140
rect 2950 6040 3030 6100
rect 2950 6000 2970 6040
rect 3010 6000 3030 6040
rect 2950 5940 3030 6000
rect 2950 5900 2970 5940
rect 3010 5900 3030 5940
rect 2950 5840 3030 5900
rect 3410 6040 3490 6070
rect 3410 6000 3430 6040
rect 3470 6000 3490 6040
rect 3410 5940 3490 6000
rect 3410 5900 3430 5940
rect 3470 5900 3490 5940
rect 3410 5870 3490 5900
rect 4020 6040 4100 6070
rect 4020 6000 4040 6040
rect 4080 6000 4100 6040
rect 4020 5940 4100 6000
rect 4020 5900 4040 5940
rect 4080 5900 4100 5940
rect 4020 5870 4100 5900
rect 2950 5800 2970 5840
rect 3010 5800 3030 5840
rect 2950 5740 3030 5800
rect 2950 5700 2970 5740
rect 3010 5700 3030 5740
rect 2950 5670 3030 5700
rect 11461 6749 11495 6811
rect 11043 5597 11077 5659
rect 11461 5597 11495 5659
rect 11043 5563 11139 5597
rect 11399 5563 11495 5597
rect -1550 4680 -1470 4710
rect -1550 4640 -1530 4680
rect -1490 4640 -1470 4680
rect -1550 4580 -1470 4640
rect -1550 4540 -1530 4580
rect -1490 4540 -1470 4580
rect -1550 4510 -1470 4540
rect 1010 4680 1090 4710
rect 1010 4640 1030 4680
rect 1070 4640 1090 4680
rect 1010 4580 1090 4640
rect 1010 4540 1030 4580
rect 1070 4540 1090 4580
rect 1010 4510 1090 4540
rect 1490 4680 1570 4710
rect 1490 4640 1510 4680
rect 1550 4640 1570 4680
rect 1490 4580 1570 4640
rect 1490 4540 1510 4580
rect 1550 4540 1570 4580
rect 1490 4510 1570 4540
rect 4050 4680 4130 4710
rect 4050 4640 4070 4680
rect 4110 4640 4130 4680
rect 4050 4580 4130 4640
rect 8490 4760 8590 4790
rect 8490 4720 8520 4760
rect 8560 4720 8590 4760
rect 8490 4660 8590 4720
rect 8490 4620 8520 4660
rect 8560 4620 8590 4660
rect 8490 4590 8590 4620
rect 9470 4760 9570 4790
rect 9470 4720 9500 4760
rect 9540 4720 9570 4760
rect 9470 4660 9570 4720
rect 9470 4620 9500 4660
rect 9540 4620 9570 4660
rect 9470 4590 9570 4620
rect 9630 4760 9730 4790
rect 9630 4720 9660 4760
rect 9700 4720 9730 4760
rect 9630 4660 9730 4720
rect 9630 4620 9660 4660
rect 9700 4620 9730 4660
rect 9630 4590 9730 4620
rect 10610 4760 10710 4790
rect 10610 4720 10640 4760
rect 10680 4720 10710 4760
rect 10610 4660 10710 4720
rect 10610 4620 10640 4660
rect 10680 4620 10710 4660
rect 10610 4590 10710 4620
rect 4050 4540 4070 4580
rect 4110 4540 4130 4580
rect 4050 4510 4130 4540
rect 11043 4347 11139 4381
rect 11399 4347 11495 4381
rect 11043 4285 11077 4347
rect 7420 4110 7520 4140
rect 7420 4070 7450 4110
rect 7490 4070 7520 4110
rect 7420 4010 7520 4070
rect 7420 3970 7450 4010
rect 7490 3970 7520 4010
rect 7420 3910 7520 3970
rect 7420 3870 7450 3910
rect 7490 3870 7520 3910
rect 7420 3810 7520 3870
rect 7420 3770 7450 3810
rect 7490 3770 7520 3810
rect 7420 3710 7520 3770
rect 7420 3670 7450 3710
rect 7490 3670 7520 3710
rect 7420 3640 7520 3670
rect 9620 4110 9720 4140
rect 9620 4070 9650 4110
rect 9690 4070 9720 4110
rect 9620 4010 9720 4070
rect 9620 3970 9650 4010
rect 9690 3970 9720 4010
rect 9620 3910 9720 3970
rect 9620 3870 9650 3910
rect 9690 3870 9720 3910
rect 9620 3810 9720 3870
rect 9620 3770 9650 3810
rect 9690 3770 9720 3810
rect 9620 3710 9720 3770
rect 9620 3670 9650 3710
rect 9690 3670 9720 3710
rect 9620 3640 9720 3670
rect 11461 4285 11495 4347
rect 11043 3077 11077 3139
rect 11461 3077 11495 3139
rect 11043 3043 11139 3077
rect 11399 3043 11495 3077
rect -551 1372 411 1391
rect -551 1338 -474 1372
rect -440 1338 -384 1372
rect -350 1338 -294 1372
rect -260 1338 -204 1372
rect -170 1338 -114 1372
rect -80 1338 -24 1372
rect 10 1338 66 1372
rect 100 1338 156 1372
rect 190 1338 246 1372
rect 280 1338 411 1372
rect -551 1319 411 1338
rect -551 1296 -479 1319
rect -551 1262 -532 1296
rect -498 1262 -479 1296
rect -551 1206 -479 1262
rect 339 1315 411 1319
rect 339 1281 358 1315
rect 392 1281 411 1315
rect -551 1172 -532 1206
rect -498 1172 -479 1206
rect -551 1116 -479 1172
rect -551 1082 -532 1116
rect -498 1082 -479 1116
rect -551 1026 -479 1082
rect -551 992 -532 1026
rect -498 992 -479 1026
rect -551 936 -479 992
rect -551 902 -532 936
rect -498 902 -479 936
rect -551 846 -479 902
rect -551 812 -532 846
rect -498 812 -479 846
rect -551 756 -479 812
rect -551 722 -532 756
rect -498 722 -479 756
rect -551 666 -479 722
rect -551 632 -532 666
rect -498 632 -479 666
rect -551 576 -479 632
rect -551 542 -532 576
rect -498 542 -479 576
rect 339 1225 411 1281
rect 339 1191 358 1225
rect 392 1191 411 1225
rect 339 1135 411 1191
rect 339 1101 358 1135
rect 392 1101 411 1135
rect 339 1045 411 1101
rect 339 1011 358 1045
rect 392 1011 411 1045
rect 339 955 411 1011
rect 339 921 358 955
rect 392 921 411 955
rect 339 865 411 921
rect 339 831 358 865
rect 392 831 411 865
rect 339 775 411 831
rect 339 741 358 775
rect 392 741 411 775
rect 339 685 411 741
rect 339 651 358 685
rect 392 651 411 685
rect 339 595 411 651
rect -551 501 -479 542
rect 339 561 358 595
rect 392 561 411 595
rect 339 501 411 561
rect -551 482 411 501
rect -551 448 -440 482
rect -406 448 -350 482
rect -316 448 -260 482
rect -226 448 -170 482
rect -136 448 -80 482
rect -46 448 10 482
rect 44 448 100 482
rect 134 448 190 482
rect 224 448 280 482
rect 314 448 411 482
rect -551 429 411 448
rect 809 1372 1771 1391
rect 809 1338 886 1372
rect 920 1338 976 1372
rect 1010 1338 1066 1372
rect 1100 1338 1156 1372
rect 1190 1338 1246 1372
rect 1280 1338 1336 1372
rect 1370 1338 1426 1372
rect 1460 1338 1516 1372
rect 1550 1338 1606 1372
rect 1640 1338 1771 1372
rect 809 1319 1771 1338
rect 809 1296 881 1319
rect 809 1262 828 1296
rect 862 1262 881 1296
rect 809 1206 881 1262
rect 1699 1315 1771 1319
rect 1699 1281 1718 1315
rect 1752 1281 1771 1315
rect 809 1172 828 1206
rect 862 1172 881 1206
rect 809 1116 881 1172
rect 809 1082 828 1116
rect 862 1082 881 1116
rect 809 1026 881 1082
rect 809 992 828 1026
rect 862 992 881 1026
rect 809 936 881 992
rect 809 902 828 936
rect 862 902 881 936
rect 809 846 881 902
rect 809 812 828 846
rect 862 812 881 846
rect 809 756 881 812
rect 809 722 828 756
rect 862 722 881 756
rect 809 666 881 722
rect 809 632 828 666
rect 862 632 881 666
rect 809 576 881 632
rect 809 542 828 576
rect 862 542 881 576
rect 1699 1225 1771 1281
rect 1699 1191 1718 1225
rect 1752 1191 1771 1225
rect 1699 1135 1771 1191
rect 1699 1101 1718 1135
rect 1752 1101 1771 1135
rect 1699 1045 1771 1101
rect 1699 1011 1718 1045
rect 1752 1011 1771 1045
rect 1699 955 1771 1011
rect 1699 921 1718 955
rect 1752 921 1771 955
rect 1699 865 1771 921
rect 1699 831 1718 865
rect 1752 831 1771 865
rect 1699 775 1771 831
rect 1699 741 1718 775
rect 1752 741 1771 775
rect 1699 685 1771 741
rect 1699 651 1718 685
rect 1752 651 1771 685
rect 1699 595 1771 651
rect 809 501 881 542
rect 1699 561 1718 595
rect 1752 561 1771 595
rect 1699 501 1771 561
rect 809 482 1771 501
rect 809 448 920 482
rect 954 448 1010 482
rect 1044 448 1100 482
rect 1134 448 1190 482
rect 1224 448 1280 482
rect 1314 448 1370 482
rect 1404 448 1460 482
rect 1494 448 1550 482
rect 1584 448 1640 482
rect 1674 448 1771 482
rect 809 429 1771 448
rect 2169 1372 3131 1391
rect 2169 1338 2246 1372
rect 2280 1338 2336 1372
rect 2370 1338 2426 1372
rect 2460 1338 2516 1372
rect 2550 1338 2606 1372
rect 2640 1338 2696 1372
rect 2730 1338 2786 1372
rect 2820 1338 2876 1372
rect 2910 1338 2966 1372
rect 3000 1338 3131 1372
rect 2169 1319 3131 1338
rect 2169 1296 2241 1319
rect 2169 1262 2188 1296
rect 2222 1262 2241 1296
rect 2169 1206 2241 1262
rect 3059 1315 3131 1319
rect 3059 1281 3078 1315
rect 3112 1281 3131 1315
rect 2169 1172 2188 1206
rect 2222 1172 2241 1206
rect 2169 1116 2241 1172
rect 2169 1082 2188 1116
rect 2222 1082 2241 1116
rect 2169 1026 2241 1082
rect 2169 992 2188 1026
rect 2222 992 2241 1026
rect 2169 936 2241 992
rect 2169 902 2188 936
rect 2222 902 2241 936
rect 2169 846 2241 902
rect 2169 812 2188 846
rect 2222 812 2241 846
rect 2169 756 2241 812
rect 2169 722 2188 756
rect 2222 722 2241 756
rect 2169 666 2241 722
rect 2169 632 2188 666
rect 2222 632 2241 666
rect 2169 576 2241 632
rect 2169 542 2188 576
rect 2222 542 2241 576
rect 3059 1225 3131 1281
rect 3059 1191 3078 1225
rect 3112 1191 3131 1225
rect 3059 1135 3131 1191
rect 3059 1101 3078 1135
rect 3112 1101 3131 1135
rect 3059 1045 3131 1101
rect 3059 1011 3078 1045
rect 3112 1011 3131 1045
rect 3059 955 3131 1011
rect 3059 921 3078 955
rect 3112 921 3131 955
rect 3059 865 3131 921
rect 3059 831 3078 865
rect 3112 831 3131 865
rect 3059 775 3131 831
rect 3059 741 3078 775
rect 3112 741 3131 775
rect 3059 685 3131 741
rect 3059 651 3078 685
rect 3112 651 3131 685
rect 3059 595 3131 651
rect 2169 501 2241 542
rect 3059 561 3078 595
rect 3112 561 3131 595
rect 3059 501 3131 561
rect 2169 482 3131 501
rect 2169 448 2280 482
rect 2314 448 2370 482
rect 2404 448 2460 482
rect 2494 448 2550 482
rect 2584 448 2640 482
rect 2674 448 2730 482
rect 2764 448 2820 482
rect 2854 448 2910 482
rect 2944 448 3000 482
rect 3034 448 3131 482
rect 2169 429 3131 448
rect -1827 149 -1731 183
rect -1139 149 -1043 183
rect -1827 87 -1793 149
rect -2940 -382 -2844 -348
rect -2252 -382 -2156 -348
rect -2940 -444 -2906 -382
rect -3727 -781 -3631 -747
rect -3371 -781 -3275 -747
rect -3727 -843 -3693 -781
rect -3309 -843 -3275 -781
rect -3727 -2233 -3693 -2171
rect -3309 -2233 -3275 -2171
rect -3727 -2267 -3631 -2233
rect -3371 -2267 -3275 -2233
rect -2190 -444 -2156 -382
rect -2940 -2236 -2906 -2174
rect -2190 -2236 -2156 -2174
rect -2940 -2270 -2844 -2236
rect -2252 -2270 -2156 -2236
rect -1077 87 -1043 149
rect -1827 -2233 -1793 -2171
rect -551 12 411 31
rect -551 -22 -474 12
rect -440 -22 -384 12
rect -350 -22 -294 12
rect -260 -22 -204 12
rect -170 -22 -114 12
rect -80 -22 -24 12
rect 10 -22 66 12
rect 100 -22 156 12
rect 190 -22 246 12
rect 280 -22 411 12
rect -551 -41 411 -22
rect -551 -64 -479 -41
rect -551 -98 -532 -64
rect -498 -98 -479 -64
rect -551 -154 -479 -98
rect 339 -45 411 -41
rect 339 -79 358 -45
rect 392 -79 411 -45
rect -551 -188 -532 -154
rect -498 -188 -479 -154
rect -551 -244 -479 -188
rect -551 -278 -532 -244
rect -498 -278 -479 -244
rect -551 -334 -479 -278
rect -551 -368 -532 -334
rect -498 -368 -479 -334
rect -551 -424 -479 -368
rect -551 -458 -532 -424
rect -498 -458 -479 -424
rect -551 -514 -479 -458
rect -551 -548 -532 -514
rect -498 -548 -479 -514
rect -551 -604 -479 -548
rect -551 -638 -532 -604
rect -498 -638 -479 -604
rect -551 -694 -479 -638
rect -551 -728 -532 -694
rect -498 -728 -479 -694
rect -551 -784 -479 -728
rect -551 -818 -532 -784
rect -498 -818 -479 -784
rect 339 -135 411 -79
rect 339 -169 358 -135
rect 392 -169 411 -135
rect 339 -225 411 -169
rect 339 -259 358 -225
rect 392 -259 411 -225
rect 339 -315 411 -259
rect 339 -349 358 -315
rect 392 -349 411 -315
rect 339 -405 411 -349
rect 339 -439 358 -405
rect 392 -439 411 -405
rect 339 -495 411 -439
rect 339 -529 358 -495
rect 392 -529 411 -495
rect 339 -585 411 -529
rect 339 -619 358 -585
rect 392 -619 411 -585
rect 339 -675 411 -619
rect 339 -709 358 -675
rect 392 -709 411 -675
rect 339 -765 411 -709
rect -551 -859 -479 -818
rect 339 -799 358 -765
rect 392 -799 411 -765
rect 339 -859 411 -799
rect -551 -878 411 -859
rect -551 -912 -440 -878
rect -406 -912 -350 -878
rect -316 -912 -260 -878
rect -226 -912 -170 -878
rect -136 -912 -80 -878
rect -46 -912 10 -878
rect 44 -912 100 -878
rect 134 -912 190 -878
rect 224 -912 280 -878
rect 314 -912 411 -878
rect -551 -931 411 -912
rect 809 12 1771 31
rect 809 -22 886 12
rect 920 -22 976 12
rect 1010 -22 1066 12
rect 1100 -22 1156 12
rect 1190 -22 1246 12
rect 1280 -22 1336 12
rect 1370 -22 1426 12
rect 1460 -22 1516 12
rect 1550 -22 1606 12
rect 1640 -22 1771 12
rect 809 -41 1771 -22
rect 809 -64 881 -41
rect 809 -98 828 -64
rect 862 -98 881 -64
rect 809 -154 881 -98
rect 1699 -45 1771 -41
rect 1699 -79 1718 -45
rect 1752 -79 1771 -45
rect 809 -188 828 -154
rect 862 -188 881 -154
rect 809 -244 881 -188
rect 809 -278 828 -244
rect 862 -278 881 -244
rect 809 -334 881 -278
rect 809 -368 828 -334
rect 862 -368 881 -334
rect 809 -424 881 -368
rect 809 -458 828 -424
rect 862 -458 881 -424
rect 809 -514 881 -458
rect 809 -548 828 -514
rect 862 -548 881 -514
rect 809 -604 881 -548
rect 809 -638 828 -604
rect 862 -638 881 -604
rect 809 -694 881 -638
rect 809 -728 828 -694
rect 862 -728 881 -694
rect 809 -784 881 -728
rect 809 -818 828 -784
rect 862 -818 881 -784
rect 1699 -135 1771 -79
rect 1699 -169 1718 -135
rect 1752 -169 1771 -135
rect 1699 -225 1771 -169
rect 1699 -259 1718 -225
rect 1752 -259 1771 -225
rect 1699 -315 1771 -259
rect 1699 -349 1718 -315
rect 1752 -349 1771 -315
rect 1699 -405 1771 -349
rect 1699 -439 1718 -405
rect 1752 -439 1771 -405
rect 1699 -495 1771 -439
rect 1699 -529 1718 -495
rect 1752 -529 1771 -495
rect 1699 -585 1771 -529
rect 1699 -619 1718 -585
rect 1752 -619 1771 -585
rect 1699 -675 1771 -619
rect 1699 -709 1718 -675
rect 1752 -709 1771 -675
rect 1699 -765 1771 -709
rect 809 -859 881 -818
rect 1699 -799 1718 -765
rect 1752 -799 1771 -765
rect 1699 -859 1771 -799
rect 809 -878 1771 -859
rect 809 -912 920 -878
rect 954 -912 1010 -878
rect 1044 -912 1100 -878
rect 1134 -912 1190 -878
rect 1224 -912 1280 -878
rect 1314 -912 1370 -878
rect 1404 -912 1460 -878
rect 1494 -912 1550 -878
rect 1584 -912 1640 -878
rect 1674 -912 1771 -878
rect 809 -931 1771 -912
rect 2169 12 3131 31
rect 2169 -22 2246 12
rect 2280 -22 2336 12
rect 2370 -22 2426 12
rect 2460 -22 2516 12
rect 2550 -22 2606 12
rect 2640 -22 2696 12
rect 2730 -22 2786 12
rect 2820 -22 2876 12
rect 2910 -22 2966 12
rect 3000 -22 3131 12
rect 2169 -41 3131 -22
rect 2169 -64 2241 -41
rect 2169 -98 2188 -64
rect 2222 -98 2241 -64
rect 2169 -154 2241 -98
rect 3059 -45 3131 -41
rect 3059 -79 3078 -45
rect 3112 -79 3131 -45
rect 2169 -188 2188 -154
rect 2222 -188 2241 -154
rect 2169 -244 2241 -188
rect 2169 -278 2188 -244
rect 2222 -278 2241 -244
rect 2169 -334 2241 -278
rect 2169 -368 2188 -334
rect 2222 -368 2241 -334
rect 2169 -424 2241 -368
rect 2169 -458 2188 -424
rect 2222 -458 2241 -424
rect 2169 -514 2241 -458
rect 2169 -548 2188 -514
rect 2222 -548 2241 -514
rect 2169 -604 2241 -548
rect 2169 -638 2188 -604
rect 2222 -638 2241 -604
rect 2169 -694 2241 -638
rect 2169 -728 2188 -694
rect 2222 -728 2241 -694
rect 2169 -784 2241 -728
rect 2169 -818 2188 -784
rect 2222 -818 2241 -784
rect 3059 -135 3131 -79
rect 3059 -169 3078 -135
rect 3112 -169 3131 -135
rect 3059 -225 3131 -169
rect 3059 -259 3078 -225
rect 3112 -259 3131 -225
rect 3059 -315 3131 -259
rect 3059 -349 3078 -315
rect 3112 -349 3131 -315
rect 3059 -405 3131 -349
rect 3059 -439 3078 -405
rect 3112 -439 3131 -405
rect 3059 -495 3131 -439
rect 3059 -529 3078 -495
rect 3112 -529 3131 -495
rect 3059 -585 3131 -529
rect 3059 -619 3078 -585
rect 3112 -619 3131 -585
rect 3059 -675 3131 -619
rect 3059 -709 3078 -675
rect 3112 -709 3131 -675
rect 3059 -765 3131 -709
rect 2169 -859 2241 -818
rect 3059 -799 3078 -765
rect 3112 -799 3131 -765
rect 3059 -859 3131 -799
rect 2169 -878 3131 -859
rect 2169 -912 2280 -878
rect 2314 -912 2370 -878
rect 2404 -912 2460 -878
rect 2494 -912 2550 -878
rect 2584 -912 2640 -878
rect 2674 -912 2730 -878
rect 2764 -912 2820 -878
rect 2854 -912 2910 -878
rect 2944 -912 3000 -878
rect 3034 -912 3131 -878
rect 2169 -931 3131 -912
rect 3493 149 3589 183
rect 4181 149 4277 183
rect 3493 87 3527 149
rect -1077 -2233 -1043 -2171
rect -1827 -2267 -1731 -2233
rect -1139 -2267 -1043 -2233
rect -551 -1348 411 -1329
rect -551 -1382 -474 -1348
rect -440 -1382 -384 -1348
rect -350 -1382 -294 -1348
rect -260 -1382 -204 -1348
rect -170 -1382 -114 -1348
rect -80 -1382 -24 -1348
rect 10 -1382 66 -1348
rect 100 -1382 156 -1348
rect 190 -1382 246 -1348
rect 280 -1382 411 -1348
rect -551 -1401 411 -1382
rect -551 -1424 -479 -1401
rect -551 -1458 -532 -1424
rect -498 -1458 -479 -1424
rect -551 -1514 -479 -1458
rect 339 -1405 411 -1401
rect 339 -1439 358 -1405
rect 392 -1439 411 -1405
rect -551 -1548 -532 -1514
rect -498 -1548 -479 -1514
rect -551 -1604 -479 -1548
rect -551 -1638 -532 -1604
rect -498 -1638 -479 -1604
rect -551 -1694 -479 -1638
rect -551 -1728 -532 -1694
rect -498 -1728 -479 -1694
rect -551 -1784 -479 -1728
rect -551 -1818 -532 -1784
rect -498 -1818 -479 -1784
rect -551 -1874 -479 -1818
rect -551 -1908 -532 -1874
rect -498 -1908 -479 -1874
rect -551 -1964 -479 -1908
rect -551 -1998 -532 -1964
rect -498 -1998 -479 -1964
rect -551 -2054 -479 -1998
rect -551 -2088 -532 -2054
rect -498 -2088 -479 -2054
rect -551 -2144 -479 -2088
rect -551 -2178 -532 -2144
rect -498 -2178 -479 -2144
rect 339 -1495 411 -1439
rect 339 -1529 358 -1495
rect 392 -1529 411 -1495
rect 339 -1585 411 -1529
rect 339 -1619 358 -1585
rect 392 -1619 411 -1585
rect 339 -1675 411 -1619
rect 339 -1709 358 -1675
rect 392 -1709 411 -1675
rect 339 -1765 411 -1709
rect 339 -1799 358 -1765
rect 392 -1799 411 -1765
rect 339 -1855 411 -1799
rect 339 -1889 358 -1855
rect 392 -1889 411 -1855
rect 339 -1945 411 -1889
rect 339 -1979 358 -1945
rect 392 -1979 411 -1945
rect 339 -2035 411 -1979
rect 339 -2069 358 -2035
rect 392 -2069 411 -2035
rect 339 -2125 411 -2069
rect -551 -2219 -479 -2178
rect 339 -2159 358 -2125
rect 392 -2159 411 -2125
rect 339 -2219 411 -2159
rect -551 -2238 411 -2219
rect -551 -2272 -440 -2238
rect -406 -2272 -350 -2238
rect -316 -2272 -260 -2238
rect -226 -2272 -170 -2238
rect -136 -2272 -80 -2238
rect -46 -2272 10 -2238
rect 44 -2272 100 -2238
rect 134 -2272 190 -2238
rect 224 -2272 280 -2238
rect 314 -2272 411 -2238
rect -551 -2291 411 -2272
rect 809 -1348 1771 -1329
rect 809 -1382 886 -1348
rect 920 -1382 976 -1348
rect 1010 -1382 1066 -1348
rect 1100 -1382 1156 -1348
rect 1190 -1382 1246 -1348
rect 1280 -1382 1336 -1348
rect 1370 -1382 1426 -1348
rect 1460 -1382 1516 -1348
rect 1550 -1382 1606 -1348
rect 1640 -1382 1771 -1348
rect 809 -1401 1771 -1382
rect 809 -1424 881 -1401
rect 809 -1458 828 -1424
rect 862 -1458 881 -1424
rect 809 -1514 881 -1458
rect 1699 -1405 1771 -1401
rect 1699 -1439 1718 -1405
rect 1752 -1439 1771 -1405
rect 809 -1548 828 -1514
rect 862 -1548 881 -1514
rect 809 -1604 881 -1548
rect 809 -1638 828 -1604
rect 862 -1638 881 -1604
rect 809 -1694 881 -1638
rect 809 -1728 828 -1694
rect 862 -1728 881 -1694
rect 809 -1784 881 -1728
rect 809 -1818 828 -1784
rect 862 -1818 881 -1784
rect 809 -1874 881 -1818
rect 809 -1908 828 -1874
rect 862 -1908 881 -1874
rect 809 -1964 881 -1908
rect 809 -1998 828 -1964
rect 862 -1998 881 -1964
rect 809 -2054 881 -1998
rect 809 -2088 828 -2054
rect 862 -2088 881 -2054
rect 809 -2144 881 -2088
rect 809 -2178 828 -2144
rect 862 -2178 881 -2144
rect 1699 -1495 1771 -1439
rect 1699 -1529 1718 -1495
rect 1752 -1529 1771 -1495
rect 1699 -1585 1771 -1529
rect 1699 -1619 1718 -1585
rect 1752 -1619 1771 -1585
rect 1699 -1675 1771 -1619
rect 1699 -1709 1718 -1675
rect 1752 -1709 1771 -1675
rect 1699 -1765 1771 -1709
rect 1699 -1799 1718 -1765
rect 1752 -1799 1771 -1765
rect 1699 -1855 1771 -1799
rect 1699 -1889 1718 -1855
rect 1752 -1889 1771 -1855
rect 1699 -1945 1771 -1889
rect 1699 -1979 1718 -1945
rect 1752 -1979 1771 -1945
rect 1699 -2035 1771 -1979
rect 1699 -2069 1718 -2035
rect 1752 -2069 1771 -2035
rect 1699 -2125 1771 -2069
rect 809 -2219 881 -2178
rect 1699 -2159 1718 -2125
rect 1752 -2159 1771 -2125
rect 1699 -2219 1771 -2159
rect 809 -2238 1771 -2219
rect 809 -2272 920 -2238
rect 954 -2272 1010 -2238
rect 1044 -2272 1100 -2238
rect 1134 -2272 1190 -2238
rect 1224 -2272 1280 -2238
rect 1314 -2272 1370 -2238
rect 1404 -2272 1460 -2238
rect 1494 -2272 1550 -2238
rect 1584 -2272 1640 -2238
rect 1674 -2272 1771 -2238
rect 809 -2291 1771 -2272
rect 2169 -1348 3131 -1329
rect 2169 -1382 2246 -1348
rect 2280 -1382 2336 -1348
rect 2370 -1382 2426 -1348
rect 2460 -1382 2516 -1348
rect 2550 -1382 2606 -1348
rect 2640 -1382 2696 -1348
rect 2730 -1382 2786 -1348
rect 2820 -1382 2876 -1348
rect 2910 -1382 2966 -1348
rect 3000 -1382 3131 -1348
rect 2169 -1401 3131 -1382
rect 2169 -1424 2241 -1401
rect 2169 -1458 2188 -1424
rect 2222 -1458 2241 -1424
rect 2169 -1514 2241 -1458
rect 3059 -1405 3131 -1401
rect 3059 -1439 3078 -1405
rect 3112 -1439 3131 -1405
rect 2169 -1548 2188 -1514
rect 2222 -1548 2241 -1514
rect 2169 -1604 2241 -1548
rect 2169 -1638 2188 -1604
rect 2222 -1638 2241 -1604
rect 2169 -1694 2241 -1638
rect 2169 -1728 2188 -1694
rect 2222 -1728 2241 -1694
rect 2169 -1784 2241 -1728
rect 2169 -1818 2188 -1784
rect 2222 -1818 2241 -1784
rect 2169 -1874 2241 -1818
rect 2169 -1908 2188 -1874
rect 2222 -1908 2241 -1874
rect 2169 -1964 2241 -1908
rect 2169 -1998 2188 -1964
rect 2222 -1998 2241 -1964
rect 2169 -2054 2241 -1998
rect 2169 -2088 2188 -2054
rect 2222 -2088 2241 -2054
rect 2169 -2144 2241 -2088
rect 2169 -2178 2188 -2144
rect 2222 -2178 2241 -2144
rect 3059 -1495 3131 -1439
rect 3059 -1529 3078 -1495
rect 3112 -1529 3131 -1495
rect 3059 -1585 3131 -1529
rect 3059 -1619 3078 -1585
rect 3112 -1619 3131 -1585
rect 3059 -1675 3131 -1619
rect 3059 -1709 3078 -1675
rect 3112 -1709 3131 -1675
rect 3059 -1765 3131 -1709
rect 3059 -1799 3078 -1765
rect 3112 -1799 3131 -1765
rect 3059 -1855 3131 -1799
rect 3059 -1889 3078 -1855
rect 3112 -1889 3131 -1855
rect 3059 -1945 3131 -1889
rect 3059 -1979 3078 -1945
rect 3112 -1979 3131 -1945
rect 3059 -2035 3131 -1979
rect 3059 -2069 3078 -2035
rect 3112 -2069 3131 -2035
rect 3059 -2125 3131 -2069
rect 2169 -2219 2241 -2178
rect 3059 -2159 3078 -2125
rect 3112 -2159 3131 -2125
rect 3059 -2219 3131 -2159
rect 2169 -2238 3131 -2219
rect 2169 -2272 2280 -2238
rect 2314 -2272 2370 -2238
rect 2404 -2272 2460 -2238
rect 2494 -2272 2550 -2238
rect 2584 -2272 2640 -2238
rect 2674 -2272 2730 -2238
rect 2764 -2272 2820 -2238
rect 2854 -2272 2910 -2238
rect 2944 -2272 3000 -2238
rect 3034 -2272 3131 -2238
rect 2169 -2291 3131 -2272
rect 4243 87 4277 149
rect 3493 -2233 3527 -2171
rect 5393 -781 5489 -747
rect 5749 -781 5845 -747
rect 5393 -843 5427 -781
rect 4243 -2233 4277 -2171
rect 3493 -2267 3589 -2233
rect 4181 -2267 4277 -2233
rect 4606 -988 4702 -954
rect 4962 -988 5058 -954
rect 4606 -1050 4640 -988
rect 5024 -1050 5058 -988
rect 4606 -2230 4640 -2168
rect 5024 -2230 5058 -2168
rect 4606 -2264 4702 -2230
rect 4962 -2264 5058 -2230
rect 5811 -843 5845 -781
rect 5393 -2233 5427 -2171
rect 5811 -2233 5845 -2171
rect 5393 -2267 5489 -2233
rect 5749 -2267 5845 -2233
rect 2863 -2949 2959 -2915
rect 5381 -2949 5477 -2915
rect 2863 -3011 2897 -2949
rect 5443 -3011 5477 -2949
rect 2863 -3333 2897 -3271
rect 5443 -3333 5477 -3271
rect 2863 -3367 2959 -3333
rect 5381 -3367 5477 -3333
<< psubdiffcont >>
rect 12240 14410 12380 14450
rect 11100 13670 11140 13880
rect 13100 13670 13140 13880
rect 6950 13240 6990 13280
rect 3710 13150 3750 13190
rect 5160 13150 5200 13190
rect 8250 13240 8290 13280
rect 9550 13240 9590 13280
rect 12240 13110 12380 13150
rect 1200 10170 1240 10210
rect 1200 10070 1240 10110
rect 2100 10170 2140 10210
rect 2100 10070 2140 10110
rect 3000 10170 3040 10210
rect 3000 10070 3040 10110
rect 3140 10170 3180 10210
rect 3140 10070 3180 10110
rect 3580 10170 3620 10210
rect 3580 10070 3620 10110
rect 3910 10170 3950 10210
rect 3910 10070 3950 10110
rect 4330 10170 4370 10210
rect 4330 10070 4370 10110
rect 4720 10170 4760 10210
rect 4720 10070 4760 10110
rect 5110 10170 5150 10210
rect 5110 10070 5150 10110
rect 7270 8620 7310 8660
rect 7270 8520 7310 8560
rect 1200 8370 1240 8410
rect 1200 8270 1240 8310
rect 2100 8370 2140 8410
rect 2100 8270 2140 8310
rect 3000 8370 3040 8410
rect 3000 8270 3040 8310
rect 3400 8370 3440 8410
rect 3400 8270 3440 8310
rect 3730 8370 3770 8410
rect 3730 8270 3770 8310
rect 4060 8370 4100 8410
rect 4060 8270 4100 8310
rect 4320 8370 4360 8410
rect 4320 8270 4360 8310
rect 5100 8370 5140 8410
rect 5100 8270 5140 8310
rect 5780 8370 5820 8410
rect 5780 8270 5820 8310
rect 7270 8420 7310 8460
rect 7270 8320 7310 8360
rect 8350 8620 8390 8660
rect 8350 8520 8390 8560
rect 8350 8420 8390 8460
rect 8350 8320 8390 8360
rect 9430 8620 9470 8660
rect 9430 8520 9470 8560
rect 9430 8420 9470 8460
rect 9430 8320 9470 8360
rect 10510 8620 10550 8660
rect 10510 8520 10550 8560
rect 10510 8420 10550 8460
rect 10510 8320 10550 8360
rect 7330 5980 7370 6030
rect 7330 5840 7370 5890
rect 9530 5980 9570 6030
rect 9530 5840 9570 5890
rect 7380 5300 7420 5340
rect 8360 5300 8400 5340
rect 9660 5300 9700 5340
rect 10640 5300 10680 5340
rect 830 3770 870 3810
rect 830 3690 870 3730
rect 830 3610 870 3650
rect 1710 3770 1750 3810
rect 1710 3690 1750 3730
rect 1710 3610 1750 3650
rect -70 3090 -30 3130
rect -70 2990 -30 3030
rect -70 2890 -30 2930
rect -70 2790 -30 2830
rect -70 2690 -30 2730
rect 2610 3090 2650 3130
rect 2610 2990 2650 3030
rect 2610 2890 2650 2930
rect 2610 2790 2650 2830
rect 2610 2690 2650 2730
rect 3430 2180 3470 2220
rect 3430 2080 3470 2120
rect -681 1462 -647 1496
rect -580 1485 -546 1519
rect -490 1485 -456 1519
rect -400 1485 -366 1519
rect -310 1485 -276 1519
rect -220 1485 -186 1519
rect -130 1485 -96 1519
rect -40 1485 -6 1519
rect 50 1485 84 1519
rect 140 1485 174 1519
rect 230 1485 264 1519
rect 320 1485 354 1519
rect 410 1485 444 1519
rect 506 1462 540 1496
rect -681 1372 -647 1406
rect -681 1282 -647 1316
rect -681 1192 -647 1226
rect -681 1102 -647 1136
rect -681 1012 -647 1046
rect -681 922 -647 956
rect -681 832 -647 866
rect -681 742 -647 776
rect -681 652 -647 686
rect -681 562 -647 596
rect -681 472 -647 506
rect 506 1372 540 1406
rect 506 1282 540 1316
rect 506 1192 540 1226
rect 506 1102 540 1136
rect 506 1012 540 1046
rect 506 922 540 956
rect 506 832 540 866
rect 506 742 540 776
rect 506 652 540 686
rect 506 562 540 596
rect 506 472 540 506
rect -681 382 -647 416
rect 506 382 540 416
rect -580 298 -546 332
rect -490 298 -456 332
rect -400 298 -366 332
rect -310 298 -276 332
rect -220 298 -186 332
rect -130 298 -96 332
rect -40 298 -6 332
rect 50 298 84 332
rect 140 298 174 332
rect 230 298 264 332
rect 320 298 354 332
rect 410 298 444 332
rect 679 1462 713 1496
rect 780 1485 814 1519
rect 870 1485 904 1519
rect 960 1485 994 1519
rect 1050 1485 1084 1519
rect 1140 1485 1174 1519
rect 1230 1485 1264 1519
rect 1320 1485 1354 1519
rect 1410 1485 1444 1519
rect 1500 1485 1534 1519
rect 1590 1485 1624 1519
rect 1680 1485 1714 1519
rect 1770 1485 1804 1519
rect 1866 1462 1900 1496
rect 679 1372 713 1406
rect 679 1282 713 1316
rect 679 1192 713 1226
rect 679 1102 713 1136
rect 679 1012 713 1046
rect 679 922 713 956
rect 679 832 713 866
rect 679 742 713 776
rect 679 652 713 686
rect 679 562 713 596
rect 679 472 713 506
rect 1866 1372 1900 1406
rect 1866 1282 1900 1316
rect 1866 1192 1900 1226
rect 1866 1102 1900 1136
rect 1866 1012 1900 1046
rect 1866 922 1900 956
rect 1866 832 1900 866
rect 1866 742 1900 776
rect 1866 652 1900 686
rect 1866 562 1900 596
rect 1866 472 1900 506
rect 679 382 713 416
rect 1866 382 1900 416
rect 780 298 814 332
rect 870 298 904 332
rect 960 298 994 332
rect 1050 298 1084 332
rect 1140 298 1174 332
rect 1230 298 1264 332
rect 1320 298 1354 332
rect 1410 298 1444 332
rect 1500 298 1534 332
rect 1590 298 1624 332
rect 1680 298 1714 332
rect 1770 298 1804 332
rect 2039 1462 2073 1496
rect 2140 1485 2174 1519
rect 2230 1485 2264 1519
rect 2320 1485 2354 1519
rect 2410 1485 2444 1519
rect 2500 1485 2534 1519
rect 2590 1485 2624 1519
rect 2680 1485 2714 1519
rect 2770 1485 2804 1519
rect 2860 1485 2894 1519
rect 2950 1485 2984 1519
rect 3040 1485 3074 1519
rect 3130 1485 3164 1519
rect 3226 1462 3260 1496
rect 2039 1372 2073 1406
rect 2039 1282 2073 1316
rect 2039 1192 2073 1226
rect 2039 1102 2073 1136
rect 2039 1012 2073 1046
rect 2039 922 2073 956
rect 2039 832 2073 866
rect 2039 742 2073 776
rect 2039 652 2073 686
rect 2039 562 2073 596
rect 2039 472 2073 506
rect 3226 1372 3260 1406
rect 3226 1282 3260 1316
rect 3226 1192 3260 1226
rect 3226 1102 3260 1136
rect 3226 1012 3260 1046
rect 3226 922 3260 956
rect 3226 832 3260 866
rect 3226 742 3260 776
rect 3226 652 3260 686
rect 3226 562 3260 596
rect 3226 472 3260 506
rect 2039 382 2073 416
rect 3226 382 3260 416
rect 2140 298 2174 332
rect 2230 298 2264 332
rect 2320 298 2354 332
rect 2410 298 2444 332
rect 2500 298 2534 332
rect 2590 298 2624 332
rect 2680 298 2714 332
rect 2770 298 2804 332
rect 2860 298 2894 332
rect 2950 298 2984 332
rect 3040 298 3074 332
rect 3130 298 3164 332
rect -681 102 -647 136
rect -580 125 -546 159
rect -490 125 -456 159
rect -400 125 -366 159
rect -310 125 -276 159
rect -220 125 -186 159
rect -130 125 -96 159
rect -40 125 -6 159
rect 50 125 84 159
rect 140 125 174 159
rect 230 125 264 159
rect 320 125 354 159
rect 410 125 444 159
rect 506 102 540 136
rect -681 12 -647 46
rect -681 -78 -647 -44
rect -681 -168 -647 -134
rect -681 -258 -647 -224
rect -681 -348 -647 -314
rect -681 -438 -647 -404
rect -681 -528 -647 -494
rect -681 -618 -647 -584
rect -681 -708 -647 -674
rect -681 -798 -647 -764
rect -681 -888 -647 -854
rect 506 12 540 46
rect 506 -78 540 -44
rect 506 -168 540 -134
rect 506 -258 540 -224
rect 506 -348 540 -314
rect 506 -438 540 -404
rect 506 -528 540 -494
rect 506 -618 540 -584
rect 506 -708 540 -674
rect 506 -798 540 -764
rect 506 -888 540 -854
rect -681 -978 -647 -944
rect 506 -978 540 -944
rect -580 -1062 -546 -1028
rect -490 -1062 -456 -1028
rect -400 -1062 -366 -1028
rect -310 -1062 -276 -1028
rect -220 -1062 -186 -1028
rect -130 -1062 -96 -1028
rect -40 -1062 -6 -1028
rect 50 -1062 84 -1028
rect 140 -1062 174 -1028
rect 230 -1062 264 -1028
rect 320 -1062 354 -1028
rect 410 -1062 444 -1028
rect 679 102 713 136
rect 780 125 814 159
rect 870 125 904 159
rect 960 125 994 159
rect 1050 125 1084 159
rect 1140 125 1174 159
rect 1230 125 1264 159
rect 1320 125 1354 159
rect 1410 125 1444 159
rect 1500 125 1534 159
rect 1590 125 1624 159
rect 1680 125 1714 159
rect 1770 125 1804 159
rect 1866 102 1900 136
rect 679 12 713 46
rect 679 -78 713 -44
rect 679 -168 713 -134
rect 679 -258 713 -224
rect 679 -348 713 -314
rect 679 -438 713 -404
rect 679 -528 713 -494
rect 679 -618 713 -584
rect 679 -708 713 -674
rect 679 -798 713 -764
rect 679 -888 713 -854
rect 1866 12 1900 46
rect 1866 -78 1900 -44
rect 1866 -168 1900 -134
rect 1866 -258 1900 -224
rect 1866 -348 1900 -314
rect 1866 -438 1900 -404
rect 1866 -528 1900 -494
rect 1866 -618 1900 -584
rect 1866 -708 1900 -674
rect 1866 -798 1900 -764
rect 1866 -888 1900 -854
rect 679 -978 713 -944
rect 1866 -978 1900 -944
rect 780 -1062 814 -1028
rect 870 -1062 904 -1028
rect 960 -1062 994 -1028
rect 1050 -1062 1084 -1028
rect 1140 -1062 1174 -1028
rect 1230 -1062 1264 -1028
rect 1320 -1062 1354 -1028
rect 1410 -1062 1444 -1028
rect 1500 -1062 1534 -1028
rect 1590 -1062 1624 -1028
rect 1680 -1062 1714 -1028
rect 1770 -1062 1804 -1028
rect 2039 102 2073 136
rect 2140 125 2174 159
rect 2230 125 2264 159
rect 2320 125 2354 159
rect 2410 125 2444 159
rect 2500 125 2534 159
rect 2590 125 2624 159
rect 2680 125 2714 159
rect 2770 125 2804 159
rect 2860 125 2894 159
rect 2950 125 2984 159
rect 3040 125 3074 159
rect 3130 125 3164 159
rect 3226 102 3260 136
rect 2039 12 2073 46
rect 2039 -78 2073 -44
rect 2039 -168 2073 -134
rect 2039 -258 2073 -224
rect 2039 -348 2073 -314
rect 2039 -438 2073 -404
rect 2039 -528 2073 -494
rect 2039 -618 2073 -584
rect 2039 -708 2073 -674
rect 2039 -798 2073 -764
rect 2039 -888 2073 -854
rect 3226 12 3260 46
rect 3226 -78 3260 -44
rect 3226 -168 3260 -134
rect 3226 -258 3260 -224
rect 3226 -348 3260 -314
rect 3226 -438 3260 -404
rect 3226 -528 3260 -494
rect 3226 -618 3260 -584
rect 3226 -708 3260 -674
rect 3226 -798 3260 -764
rect 3226 -888 3260 -854
rect 2039 -978 2073 -944
rect 3226 -978 3260 -944
rect 2140 -1062 2174 -1028
rect 2230 -1062 2264 -1028
rect 2320 -1062 2354 -1028
rect 2410 -1062 2444 -1028
rect 2500 -1062 2534 -1028
rect 2590 -1062 2624 -1028
rect 2680 -1062 2714 -1028
rect 2770 -1062 2804 -1028
rect 2860 -1062 2894 -1028
rect 2950 -1062 2984 -1028
rect 3040 -1062 3074 -1028
rect 3130 -1062 3164 -1028
rect -681 -1258 -647 -1224
rect -580 -1235 -546 -1201
rect -490 -1235 -456 -1201
rect -400 -1235 -366 -1201
rect -310 -1235 -276 -1201
rect -220 -1235 -186 -1201
rect -130 -1235 -96 -1201
rect -40 -1235 -6 -1201
rect 50 -1235 84 -1201
rect 140 -1235 174 -1201
rect 230 -1235 264 -1201
rect 320 -1235 354 -1201
rect 410 -1235 444 -1201
rect 506 -1258 540 -1224
rect -681 -1348 -647 -1314
rect -681 -1438 -647 -1404
rect -681 -1528 -647 -1494
rect -681 -1618 -647 -1584
rect -681 -1708 -647 -1674
rect -681 -1798 -647 -1764
rect -681 -1888 -647 -1854
rect -681 -1978 -647 -1944
rect -681 -2068 -647 -2034
rect -681 -2158 -647 -2124
rect -681 -2248 -647 -2214
rect 506 -1348 540 -1314
rect 506 -1438 540 -1404
rect 506 -1528 540 -1494
rect 506 -1618 540 -1584
rect 506 -1708 540 -1674
rect 506 -1798 540 -1764
rect 506 -1888 540 -1854
rect 506 -1978 540 -1944
rect 506 -2068 540 -2034
rect 506 -2158 540 -2124
rect 506 -2248 540 -2214
rect -681 -2338 -647 -2304
rect 506 -2338 540 -2304
rect -580 -2422 -546 -2388
rect -490 -2422 -456 -2388
rect -400 -2422 -366 -2388
rect -310 -2422 -276 -2388
rect -220 -2422 -186 -2388
rect -130 -2422 -96 -2388
rect -40 -2422 -6 -2388
rect 50 -2422 84 -2388
rect 140 -2422 174 -2388
rect 230 -2422 264 -2388
rect 320 -2422 354 -2388
rect 410 -2422 444 -2388
rect 679 -1258 713 -1224
rect 780 -1235 814 -1201
rect 870 -1235 904 -1201
rect 960 -1235 994 -1201
rect 1050 -1235 1084 -1201
rect 1140 -1235 1174 -1201
rect 1230 -1235 1264 -1201
rect 1320 -1235 1354 -1201
rect 1410 -1235 1444 -1201
rect 1500 -1235 1534 -1201
rect 1590 -1235 1624 -1201
rect 1680 -1235 1714 -1201
rect 1770 -1235 1804 -1201
rect 1866 -1258 1900 -1224
rect 679 -1348 713 -1314
rect 679 -1438 713 -1404
rect 679 -1528 713 -1494
rect 679 -1618 713 -1584
rect 679 -1708 713 -1674
rect 679 -1798 713 -1764
rect 679 -1888 713 -1854
rect 679 -1978 713 -1944
rect 679 -2068 713 -2034
rect 679 -2158 713 -2124
rect 679 -2248 713 -2214
rect 1866 -1348 1900 -1314
rect 1866 -1438 1900 -1404
rect 1866 -1528 1900 -1494
rect 1866 -1618 1900 -1584
rect 1866 -1708 1900 -1674
rect 1866 -1798 1900 -1764
rect 1866 -1888 1900 -1854
rect 1866 -1978 1900 -1944
rect 1866 -2068 1900 -2034
rect 1866 -2158 1900 -2124
rect 1866 -2248 1900 -2214
rect 679 -2338 713 -2304
rect 1866 -2338 1900 -2304
rect 780 -2422 814 -2388
rect 870 -2422 904 -2388
rect 960 -2422 994 -2388
rect 1050 -2422 1084 -2388
rect 1140 -2422 1174 -2388
rect 1230 -2422 1264 -2388
rect 1320 -2422 1354 -2388
rect 1410 -2422 1444 -2388
rect 1500 -2422 1534 -2388
rect 1590 -2422 1624 -2388
rect 1680 -2422 1714 -2388
rect 1770 -2422 1804 -2388
rect 2039 -1258 2073 -1224
rect 2140 -1235 2174 -1201
rect 2230 -1235 2264 -1201
rect 2320 -1235 2354 -1201
rect 2410 -1235 2444 -1201
rect 2500 -1235 2534 -1201
rect 2590 -1235 2624 -1201
rect 2680 -1235 2714 -1201
rect 2770 -1235 2804 -1201
rect 2860 -1235 2894 -1201
rect 2950 -1235 2984 -1201
rect 3040 -1235 3074 -1201
rect 3130 -1235 3164 -1201
rect 3226 -1258 3260 -1224
rect 2039 -1348 2073 -1314
rect 2039 -1438 2073 -1404
rect 2039 -1528 2073 -1494
rect 2039 -1618 2073 -1584
rect 2039 -1708 2073 -1674
rect 2039 -1798 2073 -1764
rect 2039 -1888 2073 -1854
rect 2039 -1978 2073 -1944
rect 2039 -2068 2073 -2034
rect 2039 -2158 2073 -2124
rect 2039 -2248 2073 -2214
rect 3226 -1348 3260 -1314
rect 3226 -1438 3260 -1404
rect 3226 -1528 3260 -1494
rect 3226 -1618 3260 -1584
rect 3226 -1708 3260 -1674
rect 3226 -1798 3260 -1764
rect 3226 -1888 3260 -1854
rect 3226 -1978 3260 -1944
rect 3226 -2068 3260 -2034
rect 3226 -2158 3260 -2124
rect 3226 -2248 3260 -2214
rect 2039 -2338 2073 -2304
rect 3226 -2338 3260 -2304
rect 2140 -2422 2174 -2388
rect 2230 -2422 2264 -2388
rect 2320 -2422 2354 -2388
rect 2410 -2422 2444 -2388
rect 2500 -2422 2534 -2388
rect 2590 -2422 2624 -2388
rect 2680 -2422 2714 -2388
rect 2770 -2422 2804 -2388
rect 2860 -2422 2894 -2388
rect 2950 -2422 2984 -2388
rect 3040 -2422 3074 -2388
rect 3130 -2422 3164 -2388
rect 1270 -2580 1310 -2540
rect 1270 -2660 1310 -2620
rect 1270 -2740 1310 -2700
<< nsubdiffcont >>
rect 810 12830 850 12870
rect 3180 12830 3220 12870
rect 12120 12910 12280 12950
rect 6050 12830 6090 12870
rect 7350 12830 7390 12870
rect 8650 12830 8690 12870
rect 9950 12830 9990 12870
rect 11100 11270 11140 11600
rect 13290 11270 13330 11600
rect 12120 10800 12280 10840
rect 13160 10800 13230 10840
rect 1200 9750 1240 9790
rect 1200 9650 1240 9690
rect 1200 9550 1240 9590
rect 1200 9450 1240 9490
rect 2100 9750 2140 9790
rect 2100 9650 2140 9690
rect 2100 9550 2140 9590
rect 2100 9450 2140 9490
rect 3000 9750 3040 9790
rect 3000 9650 3040 9690
rect 3000 9550 3040 9590
rect 3000 9450 3040 9490
rect 3140 9750 3180 9790
rect 3140 9650 3180 9690
rect 3140 9550 3180 9590
rect 3140 9450 3180 9490
rect 3580 9750 3620 9790
rect 3580 9650 3620 9690
rect 3580 9550 3620 9590
rect 3580 9450 3620 9490
rect 3910 9750 3950 9790
rect 3910 9650 3950 9690
rect 3910 9550 3950 9590
rect 3910 9450 3950 9490
rect 4320 9750 4360 9790
rect 4320 9650 4360 9690
rect 4320 9550 4360 9590
rect 4320 9450 4360 9490
rect 4710 9750 4750 9790
rect 4710 9650 4750 9690
rect 4710 9550 4750 9590
rect 4710 9450 4750 9490
rect 5100 9750 5140 9790
rect 5100 9650 5140 9690
rect 5100 9550 5140 9590
rect 5100 9450 5140 9490
rect 5780 9750 5820 9790
rect 5780 9650 5820 9690
rect 5780 9550 5820 9590
rect 5780 9450 5820 9490
rect 7470 9720 7510 9760
rect 7470 9620 7510 9660
rect 7470 9520 7510 9560
rect 7470 9420 7510 9460
rect 8990 9720 9030 9760
rect 8990 9620 9030 9660
rect 8990 9520 9030 9560
rect 8990 9420 9030 9460
rect 10510 9720 10550 9760
rect 10510 9620 10550 9660
rect 10510 9520 10550 9560
rect 10510 9420 10550 9460
rect 1200 8990 1240 9030
rect 1200 8890 1240 8930
rect 1200 8790 1240 8830
rect 1200 8690 1240 8730
rect 2100 8990 2140 9030
rect 2100 8890 2140 8930
rect 2100 8790 2140 8830
rect 2100 8690 2140 8730
rect 3000 8990 3040 9030
rect 3000 8890 3040 8930
rect 3000 8790 3040 8830
rect 3000 8690 3040 8730
rect 3400 8990 3440 9030
rect 3400 8890 3440 8930
rect 3400 8790 3440 8830
rect 3400 8690 3440 8730
rect 3730 8990 3770 9030
rect 3730 8890 3770 8930
rect 3730 8790 3770 8830
rect 3730 8690 3770 8730
rect 4060 8990 4100 9030
rect 4060 8890 4100 8930
rect 4060 8790 4100 8830
rect 4060 8690 4100 8730
rect 4320 8990 4360 9030
rect 4320 8890 4360 8930
rect 4320 8790 4360 8830
rect 4320 8690 4360 8730
rect 5100 8990 5140 9030
rect 5100 8890 5140 8930
rect 5100 8790 5140 8830
rect 5100 8690 5140 8730
rect -420 6800 -380 6840
rect -420 6700 -380 6740
rect 1060 6800 1100 6840
rect 1060 6700 1100 6740
rect 1480 6800 1520 6840
rect 1480 6700 1520 6740
rect 2960 6800 3000 6840
rect 2960 6700 3000 6740
rect 11139 6811 11399 6845
rect -430 6200 -390 6240
rect -430 6100 -390 6140
rect -430 6000 -390 6040
rect -430 5900 -390 5940
rect -430 5800 -390 5840
rect -430 5700 -390 5740
rect 2970 6200 3010 6240
rect 2970 6100 3010 6140
rect 2970 6000 3010 6040
rect 2970 5900 3010 5940
rect 3430 6000 3470 6040
rect 3430 5900 3470 5940
rect 4040 6000 4080 6040
rect 4040 5900 4080 5940
rect 2970 5800 3010 5840
rect 2970 5700 3010 5740
rect 11043 5659 11077 6749
rect 11461 5659 11495 6749
rect 11139 5563 11399 5597
rect -1530 4640 -1490 4680
rect -1530 4540 -1490 4580
rect 1030 4640 1070 4680
rect 1030 4540 1070 4580
rect 1510 4640 1550 4680
rect 1510 4540 1550 4580
rect 4070 4640 4110 4680
rect 8520 4720 8560 4760
rect 8520 4620 8560 4660
rect 9500 4720 9540 4760
rect 9500 4620 9540 4660
rect 9660 4720 9700 4760
rect 9660 4620 9700 4660
rect 10640 4720 10680 4760
rect 10640 4620 10680 4660
rect 4070 4540 4110 4580
rect 11139 4347 11399 4381
rect 7450 4070 7490 4110
rect 7450 3970 7490 4010
rect 7450 3870 7490 3910
rect 7450 3770 7490 3810
rect 7450 3670 7490 3710
rect 9650 4070 9690 4110
rect 9650 3970 9690 4010
rect 9650 3870 9690 3910
rect 9650 3770 9690 3810
rect 9650 3670 9690 3710
rect 11043 3139 11077 4285
rect 11461 3139 11495 4285
rect 11139 3043 11399 3077
rect -474 1338 -440 1372
rect -384 1338 -350 1372
rect -294 1338 -260 1372
rect -204 1338 -170 1372
rect -114 1338 -80 1372
rect -24 1338 10 1372
rect 66 1338 100 1372
rect 156 1338 190 1372
rect 246 1338 280 1372
rect -532 1262 -498 1296
rect 358 1281 392 1315
rect -532 1172 -498 1206
rect -532 1082 -498 1116
rect -532 992 -498 1026
rect -532 902 -498 936
rect -532 812 -498 846
rect -532 722 -498 756
rect -532 632 -498 666
rect -532 542 -498 576
rect 358 1191 392 1225
rect 358 1101 392 1135
rect 358 1011 392 1045
rect 358 921 392 955
rect 358 831 392 865
rect 358 741 392 775
rect 358 651 392 685
rect 358 561 392 595
rect -440 448 -406 482
rect -350 448 -316 482
rect -260 448 -226 482
rect -170 448 -136 482
rect -80 448 -46 482
rect 10 448 44 482
rect 100 448 134 482
rect 190 448 224 482
rect 280 448 314 482
rect 886 1338 920 1372
rect 976 1338 1010 1372
rect 1066 1338 1100 1372
rect 1156 1338 1190 1372
rect 1246 1338 1280 1372
rect 1336 1338 1370 1372
rect 1426 1338 1460 1372
rect 1516 1338 1550 1372
rect 1606 1338 1640 1372
rect 828 1262 862 1296
rect 1718 1281 1752 1315
rect 828 1172 862 1206
rect 828 1082 862 1116
rect 828 992 862 1026
rect 828 902 862 936
rect 828 812 862 846
rect 828 722 862 756
rect 828 632 862 666
rect 828 542 862 576
rect 1718 1191 1752 1225
rect 1718 1101 1752 1135
rect 1718 1011 1752 1045
rect 1718 921 1752 955
rect 1718 831 1752 865
rect 1718 741 1752 775
rect 1718 651 1752 685
rect 1718 561 1752 595
rect 920 448 954 482
rect 1010 448 1044 482
rect 1100 448 1134 482
rect 1190 448 1224 482
rect 1280 448 1314 482
rect 1370 448 1404 482
rect 1460 448 1494 482
rect 1550 448 1584 482
rect 1640 448 1674 482
rect 2246 1338 2280 1372
rect 2336 1338 2370 1372
rect 2426 1338 2460 1372
rect 2516 1338 2550 1372
rect 2606 1338 2640 1372
rect 2696 1338 2730 1372
rect 2786 1338 2820 1372
rect 2876 1338 2910 1372
rect 2966 1338 3000 1372
rect 2188 1262 2222 1296
rect 3078 1281 3112 1315
rect 2188 1172 2222 1206
rect 2188 1082 2222 1116
rect 2188 992 2222 1026
rect 2188 902 2222 936
rect 2188 812 2222 846
rect 2188 722 2222 756
rect 2188 632 2222 666
rect 2188 542 2222 576
rect 3078 1191 3112 1225
rect 3078 1101 3112 1135
rect 3078 1011 3112 1045
rect 3078 921 3112 955
rect 3078 831 3112 865
rect 3078 741 3112 775
rect 3078 651 3112 685
rect 3078 561 3112 595
rect 2280 448 2314 482
rect 2370 448 2404 482
rect 2460 448 2494 482
rect 2550 448 2584 482
rect 2640 448 2674 482
rect 2730 448 2764 482
rect 2820 448 2854 482
rect 2910 448 2944 482
rect 3000 448 3034 482
rect -1731 149 -1139 183
rect -2844 -382 -2252 -348
rect -3631 -781 -3371 -747
rect -3727 -2171 -3693 -843
rect -3309 -2171 -3275 -843
rect -3631 -2267 -3371 -2233
rect -2940 -2174 -2906 -444
rect -2190 -2174 -2156 -444
rect -2844 -2270 -2252 -2236
rect -1827 -2171 -1793 87
rect -1077 -2171 -1043 87
rect -474 -22 -440 12
rect -384 -22 -350 12
rect -294 -22 -260 12
rect -204 -22 -170 12
rect -114 -22 -80 12
rect -24 -22 10 12
rect 66 -22 100 12
rect 156 -22 190 12
rect 246 -22 280 12
rect -532 -98 -498 -64
rect 358 -79 392 -45
rect -532 -188 -498 -154
rect -532 -278 -498 -244
rect -532 -368 -498 -334
rect -532 -458 -498 -424
rect -532 -548 -498 -514
rect -532 -638 -498 -604
rect -532 -728 -498 -694
rect -532 -818 -498 -784
rect 358 -169 392 -135
rect 358 -259 392 -225
rect 358 -349 392 -315
rect 358 -439 392 -405
rect 358 -529 392 -495
rect 358 -619 392 -585
rect 358 -709 392 -675
rect 358 -799 392 -765
rect -440 -912 -406 -878
rect -350 -912 -316 -878
rect -260 -912 -226 -878
rect -170 -912 -136 -878
rect -80 -912 -46 -878
rect 10 -912 44 -878
rect 100 -912 134 -878
rect 190 -912 224 -878
rect 280 -912 314 -878
rect 886 -22 920 12
rect 976 -22 1010 12
rect 1066 -22 1100 12
rect 1156 -22 1190 12
rect 1246 -22 1280 12
rect 1336 -22 1370 12
rect 1426 -22 1460 12
rect 1516 -22 1550 12
rect 1606 -22 1640 12
rect 828 -98 862 -64
rect 1718 -79 1752 -45
rect 828 -188 862 -154
rect 828 -278 862 -244
rect 828 -368 862 -334
rect 828 -458 862 -424
rect 828 -548 862 -514
rect 828 -638 862 -604
rect 828 -728 862 -694
rect 828 -818 862 -784
rect 1718 -169 1752 -135
rect 1718 -259 1752 -225
rect 1718 -349 1752 -315
rect 1718 -439 1752 -405
rect 1718 -529 1752 -495
rect 1718 -619 1752 -585
rect 1718 -709 1752 -675
rect 1718 -799 1752 -765
rect 920 -912 954 -878
rect 1010 -912 1044 -878
rect 1100 -912 1134 -878
rect 1190 -912 1224 -878
rect 1280 -912 1314 -878
rect 1370 -912 1404 -878
rect 1460 -912 1494 -878
rect 1550 -912 1584 -878
rect 1640 -912 1674 -878
rect 2246 -22 2280 12
rect 2336 -22 2370 12
rect 2426 -22 2460 12
rect 2516 -22 2550 12
rect 2606 -22 2640 12
rect 2696 -22 2730 12
rect 2786 -22 2820 12
rect 2876 -22 2910 12
rect 2966 -22 3000 12
rect 2188 -98 2222 -64
rect 3078 -79 3112 -45
rect 2188 -188 2222 -154
rect 2188 -278 2222 -244
rect 2188 -368 2222 -334
rect 2188 -458 2222 -424
rect 2188 -548 2222 -514
rect 2188 -638 2222 -604
rect 2188 -728 2222 -694
rect 2188 -818 2222 -784
rect 3078 -169 3112 -135
rect 3078 -259 3112 -225
rect 3078 -349 3112 -315
rect 3078 -439 3112 -405
rect 3078 -529 3112 -495
rect 3078 -619 3112 -585
rect 3078 -709 3112 -675
rect 3078 -799 3112 -765
rect 2280 -912 2314 -878
rect 2370 -912 2404 -878
rect 2460 -912 2494 -878
rect 2550 -912 2584 -878
rect 2640 -912 2674 -878
rect 2730 -912 2764 -878
rect 2820 -912 2854 -878
rect 2910 -912 2944 -878
rect 3000 -912 3034 -878
rect 3589 149 4181 183
rect -1731 -2267 -1139 -2233
rect -474 -1382 -440 -1348
rect -384 -1382 -350 -1348
rect -294 -1382 -260 -1348
rect -204 -1382 -170 -1348
rect -114 -1382 -80 -1348
rect -24 -1382 10 -1348
rect 66 -1382 100 -1348
rect 156 -1382 190 -1348
rect 246 -1382 280 -1348
rect -532 -1458 -498 -1424
rect 358 -1439 392 -1405
rect -532 -1548 -498 -1514
rect -532 -1638 -498 -1604
rect -532 -1728 -498 -1694
rect -532 -1818 -498 -1784
rect -532 -1908 -498 -1874
rect -532 -1998 -498 -1964
rect -532 -2088 -498 -2054
rect -532 -2178 -498 -2144
rect 358 -1529 392 -1495
rect 358 -1619 392 -1585
rect 358 -1709 392 -1675
rect 358 -1799 392 -1765
rect 358 -1889 392 -1855
rect 358 -1979 392 -1945
rect 358 -2069 392 -2035
rect 358 -2159 392 -2125
rect -440 -2272 -406 -2238
rect -350 -2272 -316 -2238
rect -260 -2272 -226 -2238
rect -170 -2272 -136 -2238
rect -80 -2272 -46 -2238
rect 10 -2272 44 -2238
rect 100 -2272 134 -2238
rect 190 -2272 224 -2238
rect 280 -2272 314 -2238
rect 886 -1382 920 -1348
rect 976 -1382 1010 -1348
rect 1066 -1382 1100 -1348
rect 1156 -1382 1190 -1348
rect 1246 -1382 1280 -1348
rect 1336 -1382 1370 -1348
rect 1426 -1382 1460 -1348
rect 1516 -1382 1550 -1348
rect 1606 -1382 1640 -1348
rect 828 -1458 862 -1424
rect 1718 -1439 1752 -1405
rect 828 -1548 862 -1514
rect 828 -1638 862 -1604
rect 828 -1728 862 -1694
rect 828 -1818 862 -1784
rect 828 -1908 862 -1874
rect 828 -1998 862 -1964
rect 828 -2088 862 -2054
rect 828 -2178 862 -2144
rect 1718 -1529 1752 -1495
rect 1718 -1619 1752 -1585
rect 1718 -1709 1752 -1675
rect 1718 -1799 1752 -1765
rect 1718 -1889 1752 -1855
rect 1718 -1979 1752 -1945
rect 1718 -2069 1752 -2035
rect 1718 -2159 1752 -2125
rect 920 -2272 954 -2238
rect 1010 -2272 1044 -2238
rect 1100 -2272 1134 -2238
rect 1190 -2272 1224 -2238
rect 1280 -2272 1314 -2238
rect 1370 -2272 1404 -2238
rect 1460 -2272 1494 -2238
rect 1550 -2272 1584 -2238
rect 1640 -2272 1674 -2238
rect 2246 -1382 2280 -1348
rect 2336 -1382 2370 -1348
rect 2426 -1382 2460 -1348
rect 2516 -1382 2550 -1348
rect 2606 -1382 2640 -1348
rect 2696 -1382 2730 -1348
rect 2786 -1382 2820 -1348
rect 2876 -1382 2910 -1348
rect 2966 -1382 3000 -1348
rect 2188 -1458 2222 -1424
rect 3078 -1439 3112 -1405
rect 2188 -1548 2222 -1514
rect 2188 -1638 2222 -1604
rect 2188 -1728 2222 -1694
rect 2188 -1818 2222 -1784
rect 2188 -1908 2222 -1874
rect 2188 -1998 2222 -1964
rect 2188 -2088 2222 -2054
rect 2188 -2178 2222 -2144
rect 3078 -1529 3112 -1495
rect 3078 -1619 3112 -1585
rect 3078 -1709 3112 -1675
rect 3078 -1799 3112 -1765
rect 3078 -1889 3112 -1855
rect 3078 -1979 3112 -1945
rect 3078 -2069 3112 -2035
rect 3078 -2159 3112 -2125
rect 2280 -2272 2314 -2238
rect 2370 -2272 2404 -2238
rect 2460 -2272 2494 -2238
rect 2550 -2272 2584 -2238
rect 2640 -2272 2674 -2238
rect 2730 -2272 2764 -2238
rect 2820 -2272 2854 -2238
rect 2910 -2272 2944 -2238
rect 3000 -2272 3034 -2238
rect 3493 -2171 3527 87
rect 4243 -2171 4277 87
rect 5489 -781 5749 -747
rect 3589 -2267 4181 -2233
rect 4702 -988 4962 -954
rect 4606 -2168 4640 -1050
rect 5024 -2168 5058 -1050
rect 4702 -2264 4962 -2230
rect 5393 -2171 5427 -843
rect 5811 -2171 5845 -843
rect 5489 -2267 5749 -2233
rect 2959 -2949 5381 -2915
rect 2863 -3271 2897 -3011
rect 5443 -3271 5477 -3011
rect 2959 -3367 5381 -3333
<< poly >>
rect 11290 14350 11320 14380
rect 11810 14350 11840 14380
rect 12330 14350 12360 14380
rect 12930 14350 12960 14380
rect 11290 14120 11320 14150
rect 11810 14120 11840 14150
rect 12330 14120 12360 14150
rect 12930 14120 12960 14150
rect 11276 14102 11334 14120
rect 11276 14068 11288 14102
rect 11322 14068 11334 14102
rect 11276 14050 11334 14068
rect 11796 14102 11854 14120
rect 11796 14068 11808 14102
rect 11842 14068 11854 14102
rect 11796 14050 11854 14068
rect 12316 14102 12374 14120
rect 12316 14068 12328 14102
rect 12362 14068 12374 14102
rect 12316 14050 12374 14068
rect 12884 14102 12960 14120
rect 12884 14068 12896 14102
rect 12930 14068 12960 14102
rect 12884 14050 12960 14068
rect 11290 13970 11320 14000
rect 11810 13970 11840 14000
rect 12330 13970 12360 14000
rect 390 13310 470 13330
rect 390 13270 410 13310
rect 450 13270 470 13310
rect 390 13250 470 13270
rect 1340 13290 1420 13310
rect 1340 13250 1360 13290
rect 1400 13250 1420 13290
rect 2410 13300 2490 13320
rect 2410 13260 2430 13300
rect 2470 13260 2490 13300
rect 2410 13250 2490 13260
rect 3970 13300 4060 13320
rect 3970 13260 3990 13300
rect 4030 13260 4060 13300
rect 3970 13250 4060 13260
rect 6584 13310 6650 13330
rect 7150 13310 7180 13340
rect 7260 13310 7290 13340
rect 7370 13310 7400 13340
rect 7480 13310 7510 13340
rect 7810 13310 7840 13340
rect 7920 13310 7950 13340
rect 8030 13310 8060 13340
rect 8450 13310 8480 13340
rect 8560 13310 8590 13340
rect 8670 13310 8700 13340
rect 8780 13310 8810 13340
rect 9110 13310 9140 13340
rect 9220 13310 9250 13340
rect 9330 13310 9360 13340
rect 9750 13310 9780 13340
rect 9860 13310 9890 13340
rect 9970 13310 10000 13340
rect 10080 13310 10110 13340
rect 10410 13310 10440 13340
rect 10520 13310 10550 13340
rect 10630 13310 10660 13340
rect 6584 13270 6594 13310
rect 6634 13270 6650 13310
rect 6584 13250 6650 13270
rect 520 13220 550 13250
rect 630 13220 660 13250
rect 740 13220 770 13250
rect 850 13220 880 13250
rect 1100 13220 1130 13250
rect 1210 13220 1240 13250
rect 1340 13230 1420 13250
rect 520 13090 550 13120
rect 630 13100 660 13120
rect 740 13100 770 13120
rect 850 13100 880 13120
rect 1100 13100 1130 13120
rect 630 13090 1130 13100
rect 500 13070 580 13090
rect 630 13070 1160 13090
rect 500 13030 520 13070
rect 560 13030 580 13070
rect 500 13010 580 13030
rect 680 12900 710 13070
rect 1080 13030 1100 13070
rect 1140 13030 1160 13070
rect 1080 13010 1160 13030
rect 1210 12990 1240 13120
rect 1340 12990 1370 13230
rect 1550 13220 1580 13250
rect 1660 13220 1690 13250
rect 1770 13220 1800 13250
rect 1880 13220 1910 13250
rect 2210 13220 2240 13250
rect 2320 13220 2350 13250
rect 2430 13220 2460 13250
rect 2540 13220 2570 13250
rect 2890 13220 2920 13250
rect 3000 13220 3030 13250
rect 3110 13220 3140 13250
rect 3220 13220 3250 13250
rect 3470 13220 3500 13250
rect 3580 13220 3610 13250
rect 4030 13220 4060 13250
rect 4390 13220 4420 13250
rect 4640 13220 4670 13250
rect 4750 13220 4780 13250
rect 4860 13220 4890 13250
rect 4970 13220 5000 13250
rect 5300 13220 5330 13250
rect 5410 13220 5440 13250
rect 5520 13220 5550 13250
rect 5850 13220 5880 13250
rect 5960 13220 5990 13250
rect 6070 13220 6100 13250
rect 6180 13220 6210 13250
rect 6510 13220 6540 13250
rect 6620 13220 6650 13250
rect 6730 13220 6760 13250
rect 7150 13180 7180 13210
rect 7260 13190 7290 13210
rect 7370 13190 7400 13210
rect 7480 13190 7510 13210
rect 7810 13190 7840 13210
rect 7130 13160 7210 13180
rect 7130 13120 7150 13160
rect 7190 13120 7210 13160
rect 1420 13070 1500 13090
rect 1420 13030 1440 13070
rect 1480 13030 1500 13070
rect 1420 13010 1500 13030
rect 1550 13010 1580 13120
rect 1660 13090 1690 13120
rect 1770 13090 1800 13120
rect 1880 13090 1910 13120
rect 1660 13070 2080 13090
rect 1660 13060 2020 13070
rect 1210 12960 1370 12990
rect 1550 12990 1700 13010
rect 1550 12980 1640 12990
rect 1100 12900 1130 12930
rect 1210 12900 1240 12960
rect 370 12870 450 12890
rect 370 12830 390 12870
rect 430 12830 450 12870
rect 370 12810 450 12830
rect 680 12770 710 12800
rect 1100 12770 1130 12800
rect 1210 12770 1240 12800
rect 1340 12790 1370 12960
rect 1620 12950 1640 12980
rect 1680 12950 1700 12990
rect 1620 12930 1700 12950
rect 1770 12900 1800 13060
rect 2000 13030 2020 13060
rect 2060 13030 2080 13070
rect 2000 13020 2080 13030
rect 2020 12960 2100 12970
rect 1880 12950 2100 12960
rect 1880 12930 2040 12950
rect 1880 12900 1910 12930
rect 2020 12910 2040 12930
rect 2080 12910 2100 12950
rect 2020 12890 2100 12910
rect 2210 12900 2240 13120
rect 2320 12900 2350 13120
rect 2430 12900 2460 13120
rect 2540 13090 2570 13120
rect 2890 13090 2920 13120
rect 3000 13100 3030 13120
rect 3110 13100 3140 13120
rect 3220 13100 3250 13120
rect 3470 13100 3500 13120
rect 3000 13090 3500 13100
rect 2520 13070 2750 13090
rect 2520 13030 2540 13070
rect 2580 13060 2750 13070
rect 2580 13030 2600 13060
rect 2520 13020 2600 13030
rect 2720 12970 2750 13060
rect 2870 13070 2950 13090
rect 3000 13070 3530 13090
rect 2870 13030 2890 13070
rect 2930 13030 2950 13070
rect 2870 13020 2950 13030
rect 3050 12970 3080 13070
rect 3450 13030 3470 13070
rect 3510 13030 3530 13070
rect 3450 13010 3530 13030
rect 2720 12940 3080 12970
rect 3050 12900 3080 12940
rect 3580 12970 3610 13120
rect 3660 13070 3740 13090
rect 3660 13030 3680 13070
rect 3720 13060 3740 13070
rect 3900 13070 3980 13090
rect 3900 13060 3920 13070
rect 3720 13030 3920 13060
rect 3960 13030 3980 13070
rect 3660 13020 3740 13030
rect 3900 13010 3980 13030
rect 3580 12950 3800 12970
rect 4030 12950 4060 13120
rect 4240 13060 4320 13080
rect 4240 13020 4260 13060
rect 4300 13020 4320 13060
rect 4240 13000 4320 13020
rect 4390 13020 4420 13120
rect 4510 13020 4590 13040
rect 4390 12990 4530 13020
rect 4390 12950 4420 12990
rect 4510 12980 4530 12990
rect 4570 12980 4590 13020
rect 4640 13010 4670 13120
rect 4750 13090 4780 13120
rect 4860 13090 4890 13120
rect 4970 13090 5000 13120
rect 4750 13070 5220 13090
rect 4750 13060 5160 13070
rect 4640 12990 4790 13010
rect 4640 12980 4730 12990
rect 4510 12960 4590 12980
rect 3580 12940 3740 12950
rect 3470 12900 3500 12930
rect 3580 12900 3610 12940
rect 3720 12910 3740 12940
rect 3780 12910 3800 12950
rect 3720 12890 3800 12910
rect 3920 12920 4060 12950
rect 3920 12900 3950 12920
rect 4030 12900 4060 12920
rect 4280 12920 4420 12950
rect 4710 12950 4730 12980
rect 4770 12950 4790 12990
rect 4710 12930 4790 12950
rect 4280 12900 4310 12920
rect 4390 12900 4420 12920
rect 4860 12900 4890 13060
rect 5140 13030 5160 13060
rect 5200 13030 5220 13070
rect 5140 13020 5220 13030
rect 5110 12960 5190 12970
rect 4970 12950 5190 12960
rect 4970 12930 5130 12950
rect 4970 12900 5000 12930
rect 5110 12910 5130 12930
rect 5170 12910 5190 12950
rect 5110 12890 5190 12910
rect 5300 12900 5330 13120
rect 5410 12970 5440 13120
rect 5520 13090 5550 13120
rect 5850 13090 5880 13120
rect 5960 13100 5990 13120
rect 6070 13100 6100 13120
rect 6180 13100 6210 13120
rect 6510 13100 6540 13120
rect 5500 13070 5710 13090
rect 5500 13030 5520 13070
rect 5560 13060 5710 13070
rect 5560 13030 5580 13060
rect 5500 13020 5580 13030
rect 5680 12970 5710 13060
rect 5830 13070 5910 13090
rect 5830 13030 5850 13070
rect 5890 13030 5910 13070
rect 5830 13020 5910 13030
rect 5960 13070 6540 13100
rect 5960 12970 5990 13070
rect 6410 13030 6430 13070
rect 6470 13030 6490 13070
rect 6410 13010 6490 13030
rect 6620 13010 6650 13120
rect 5410 12940 5570 12970
rect 5680 12940 5990 12970
rect 6240 12990 6320 13010
rect 6240 12950 6260 12990
rect 6300 12950 6320 12990
rect 6540 12980 6650 13010
rect 6730 13040 6760 13120
rect 7130 13100 7210 13120
rect 7260 13160 7840 13190
rect 6880 13050 6960 13070
rect 6880 13040 6900 13050
rect 6730 13010 6900 13040
rect 6940 13010 6960 13050
rect 6540 12950 6570 12980
rect 5410 12900 5440 12940
rect 5540 12890 5570 12940
rect 5920 12900 5950 12940
rect 6240 12930 6320 12950
rect 6260 12900 6290 12930
rect 6370 12920 6570 12950
rect 6370 12900 6400 12920
rect 6620 12900 6650 12930
rect 6730 12900 6760 13010
rect 6880 12990 6960 13010
rect 7260 12960 7290 13160
rect 7710 13120 7730 13160
rect 7770 13120 7790 13160
rect 7710 13100 7790 13120
rect 7920 13040 7950 13210
rect 7670 13010 7950 13040
rect 8030 13040 8060 13210
rect 8450 13180 8480 13210
rect 8560 13190 8590 13210
rect 8670 13190 8700 13210
rect 8780 13190 8810 13210
rect 9110 13190 9140 13210
rect 8430 13160 8510 13180
rect 8430 13120 8450 13160
rect 8490 13120 8510 13160
rect 8430 13100 8510 13120
rect 8560 13160 9140 13190
rect 8180 13050 8260 13070
rect 8180 13040 8200 13050
rect 8030 13010 8200 13040
rect 8240 13010 8260 13050
rect 7220 12930 7290 12960
rect 7540 12990 7620 13010
rect 7540 12950 7560 12990
rect 7600 12950 7620 12990
rect 7540 12930 7620 12950
rect 7220 12900 7250 12930
rect 7560 12900 7590 12930
rect 7670 12900 7700 13010
rect 7920 12900 7950 12930
rect 8030 12900 8060 13010
rect 8180 12990 8260 13010
rect 8560 12960 8590 13160
rect 9010 13120 9030 13160
rect 9070 13120 9090 13160
rect 9010 13100 9090 13120
rect 9220 13040 9250 13210
rect 8970 13010 9250 13040
rect 9330 13040 9360 13210
rect 9750 13180 9780 13210
rect 9860 13190 9890 13210
rect 9970 13190 10000 13210
rect 10080 13190 10110 13210
rect 10410 13190 10440 13210
rect 9730 13160 9810 13180
rect 9730 13120 9750 13160
rect 9790 13120 9810 13160
rect 9730 13100 9810 13120
rect 9860 13160 10440 13190
rect 9480 13050 9560 13070
rect 9480 13040 9500 13050
rect 9330 13010 9500 13040
rect 9540 13010 9560 13050
rect 8520 12930 8590 12960
rect 8840 12990 8920 13010
rect 8840 12950 8860 12990
rect 8900 12950 8920 12990
rect 8840 12930 8920 12950
rect 8520 12900 8550 12930
rect 8860 12900 8890 12930
rect 8970 12900 9000 13010
rect 9220 12900 9250 12930
rect 9330 12900 9360 13010
rect 9480 12990 9560 13010
rect 9860 12960 9890 13160
rect 10310 13120 10330 13160
rect 10370 13120 10390 13160
rect 10310 13100 10390 13120
rect 10520 13040 10550 13210
rect 10270 13010 10550 13040
rect 10630 13040 10660 13210
rect 11290 13640 11320 13670
rect 11810 13640 11840 13670
rect 12330 13640 12360 13670
rect 11290 13622 11348 13640
rect 11290 13588 11302 13622
rect 11336 13588 11348 13622
rect 11290 13570 11348 13588
rect 11810 13622 11868 13640
rect 11810 13588 11822 13622
rect 11856 13588 11868 13622
rect 11810 13570 11868 13588
rect 12330 13622 12388 13640
rect 12330 13588 12342 13622
rect 12376 13588 12388 13622
rect 12330 13570 12388 13588
rect 11288 13490 11320 13520
rect 11808 13490 11840 13520
rect 12328 13490 12360 13520
rect 11288 13260 11320 13290
rect 11808 13260 11840 13290
rect 12328 13260 12360 13290
rect 11262 13242 11320 13260
rect 11262 13208 11274 13242
rect 11308 13208 11320 13242
rect 11262 13190 11320 13208
rect 11782 13242 11840 13260
rect 11782 13208 11794 13242
rect 11828 13208 11840 13242
rect 11782 13190 11840 13208
rect 12302 13242 12360 13260
rect 12302 13208 12314 13242
rect 12348 13208 12360 13242
rect 12302 13190 12360 13208
rect 10762 13042 10820 13070
rect 10762 13040 10774 13042
rect 10630 13010 10774 13040
rect 9820 12930 9890 12960
rect 10140 12990 10220 13010
rect 10140 12950 10160 12990
rect 10200 12950 10220 12990
rect 10140 12930 10220 12950
rect 9820 12900 9850 12930
rect 10160 12900 10190 12930
rect 10270 12900 10300 13010
rect 10520 12900 10550 12930
rect 10630 12900 10660 13010
rect 10762 13008 10774 13010
rect 10808 13008 10820 13042
rect 10762 12990 10820 13008
rect 5540 12870 5780 12890
rect 5540 12860 5720 12870
rect 5700 12830 5720 12860
rect 5760 12830 5780 12870
rect 5700 12810 5780 12830
rect 1340 12770 1420 12790
rect 1770 12770 1800 12800
rect 1880 12770 1910 12800
rect 2210 12770 2240 12800
rect 2320 12770 2350 12800
rect 2430 12770 2460 12800
rect 3050 12770 3080 12800
rect 3470 12770 3500 12800
rect 3580 12770 3610 12800
rect 3920 12770 3950 12800
rect 4030 12770 4060 12800
rect 4280 12770 4310 12800
rect 4390 12770 4420 12800
rect 4860 12770 4890 12800
rect 4970 12770 5000 12800
rect 1030 12750 1130 12770
rect 1030 12710 1050 12750
rect 1090 12710 1130 12750
rect 1340 12730 1360 12770
rect 1400 12730 1420 12770
rect 1340 12710 1420 12730
rect 2150 12750 2240 12770
rect 2150 12710 2170 12750
rect 2210 12710 2240 12750
rect 1030 12690 1130 12710
rect 2150 12690 2240 12710
rect 2290 12750 2350 12770
rect 2290 12710 2300 12750
rect 2340 12710 2350 12750
rect 2290 12690 2350 12710
rect 3410 12750 3500 12770
rect 5300 12760 5330 12800
rect 5410 12770 5440 12800
rect 5920 12770 5950 12800
rect 6260 12770 6290 12800
rect 6370 12770 6400 12800
rect 6620 12780 6650 12800
rect 6730 12780 6760 12800
rect 3410 12710 3430 12750
rect 3470 12710 3500 12750
rect 3410 12690 3500 12710
rect 5170 12740 5330 12760
rect 6620 12750 6760 12780
rect 7220 12770 7250 12800
rect 7560 12770 7590 12800
rect 7670 12770 7700 12800
rect 7920 12780 7950 12800
rect 8030 12780 8060 12800
rect 7670 12750 7780 12770
rect 7920 12750 8060 12780
rect 8520 12770 8550 12800
rect 8860 12770 8890 12800
rect 8970 12770 9000 12800
rect 9220 12780 9250 12800
rect 9330 12780 9360 12800
rect 8970 12750 9080 12770
rect 9220 12750 9360 12780
rect 9820 12770 9850 12800
rect 10160 12770 10190 12800
rect 10270 12770 10300 12800
rect 10520 12780 10550 12800
rect 10630 12780 10660 12800
rect 10270 12750 10380 12770
rect 10520 12750 10660 12780
rect 5170 12700 5190 12740
rect 5230 12730 5330 12740
rect 5230 12700 5250 12730
rect 5170 12690 5250 12700
rect 7670 12710 7720 12750
rect 7760 12710 7780 12750
rect 7670 12690 7780 12710
rect 8970 12710 9020 12750
rect 9060 12710 9080 12750
rect 8970 12690 9080 12710
rect 10270 12710 10320 12750
rect 10360 12710 10380 12750
rect 10270 12690 10380 12710
rect 11262 12852 11320 12870
rect 11262 12818 11274 12852
rect 11308 12818 11320 12852
rect 11262 12800 11320 12818
rect 11782 12852 11840 12870
rect 11782 12818 11794 12852
rect 11828 12818 11840 12852
rect 11782 12800 11840 12818
rect 12302 12852 12360 12870
rect 12302 12818 12314 12852
rect 12348 12818 12360 12852
rect 12302 12800 12360 12818
rect 11288 12770 11320 12800
rect 11808 12770 11840 12800
rect 12328 12770 12360 12800
rect 11288 12340 11320 12370
rect 11808 12340 11840 12370
rect 12328 12340 12360 12370
rect 11290 12272 11348 12290
rect 11290 12238 11302 12272
rect 11336 12238 11348 12272
rect 11290 12220 11348 12238
rect 11810 12272 11868 12290
rect 11810 12238 11822 12272
rect 11856 12238 11868 12272
rect 11810 12220 11868 12238
rect 12330 12272 12388 12290
rect 12330 12238 12342 12272
rect 12376 12238 12388 12272
rect 12330 12220 12388 12238
rect 11290 12190 11320 12220
rect 11810 12190 11840 12220
rect 12330 12190 12360 12220
rect 11290 11560 11320 11590
rect 11810 11560 11840 11590
rect 12330 11560 12360 11590
rect 11400 11390 11480 11410
rect 11400 11350 11420 11390
rect 11460 11350 11480 11390
rect 11400 11330 11480 11350
rect 11920 11390 12000 11410
rect 11920 11350 11940 11390
rect 11980 11350 12000 11390
rect 11920 11330 12000 11350
rect 12440 11390 12520 11410
rect 12440 11350 12460 11390
rect 12500 11350 12520 11390
rect 12440 11330 12520 11350
rect 12970 11390 13030 11410
rect 12970 11350 12980 11390
rect 13020 11350 13030 11390
rect 12970 11330 13030 11350
rect 11290 11300 11590 11330
rect 11810 11300 12110 11330
rect 12330 11300 12630 11330
rect 12850 11300 13150 11330
rect 11290 10870 11590 10900
rect 11810 10870 12110 10900
rect 12330 10870 12630 10900
rect 12850 10870 13150 10900
rect 1860 10320 2270 10350
rect 1340 10240 1370 10270
rect 1450 10240 1480 10270
rect 1860 10240 1890 10320
rect 1970 10240 2000 10270
rect 2240 10240 2270 10320
rect 3390 10330 3470 10350
rect 3390 10290 3410 10330
rect 3450 10290 3470 10330
rect 3390 10270 3470 10290
rect 2350 10240 2380 10270
rect 2760 10240 2790 10270
rect 2870 10240 2900 10270
rect 3280 10240 3310 10270
rect 3390 10240 3420 10270
rect 3720 10240 3750 10270
rect 4050 10240 4080 10270
rect 4490 10240 4520 10270
rect 4880 10240 4910 10270
rect 5270 10240 5300 10270
rect 5560 10240 5590 10270
rect 1340 9970 1370 10040
rect 1140 9950 1370 9970
rect 1140 9910 1160 9950
rect 1200 9940 1370 9950
rect 1200 9910 1220 9940
rect 1140 9890 1220 9910
rect 1340 9820 1370 9940
rect 1450 10010 1480 10040
rect 1450 9990 1550 10010
rect 1860 10000 1890 10040
rect 1450 9950 1490 9990
rect 1530 9950 1550 9990
rect 1450 9930 1550 9950
rect 1640 9970 1890 10000
rect 1450 9820 1480 9930
rect 1640 9510 1670 9970
rect 1860 9820 1890 9970
rect 1970 9930 2000 10040
rect 1970 9910 2070 9930
rect 1970 9870 2010 9910
rect 2050 9870 2070 9910
rect 1970 9850 2070 9870
rect 1970 9820 2000 9850
rect 2240 9820 2270 10040
rect 2350 10010 2380 10040
rect 2350 9990 2450 10010
rect 2760 10000 2790 10040
rect 2350 9950 2390 9990
rect 2430 9950 2450 9990
rect 2350 9930 2450 9950
rect 2540 9970 2790 10000
rect 2350 9820 2380 9930
rect 1590 9490 1670 9510
rect 1590 9450 1610 9490
rect 1650 9450 1670 9490
rect 1590 9430 1670 9450
rect 2540 9510 2570 9970
rect 2760 9820 2790 9970
rect 2870 10000 2900 10040
rect 2870 9980 3120 10000
rect 2870 9970 3060 9980
rect 2870 9820 2900 9970
rect 3040 9940 3060 9970
rect 3100 9940 3120 9980
rect 3040 9920 3120 9940
rect 3280 9820 3310 10040
rect 3390 9820 3420 10040
rect 3470 9940 3550 9960
rect 3720 9940 3750 10040
rect 3470 9900 3490 9940
rect 3530 9910 3750 9940
rect 3530 9900 3550 9910
rect 3470 9880 3550 9900
rect 3720 9820 3750 9910
rect 3800 9940 3880 9960
rect 4050 9940 4080 10040
rect 4260 9970 4340 9990
rect 3800 9900 3820 9940
rect 3860 9910 4080 9940
rect 3860 9900 3880 9910
rect 3800 9880 3880 9900
rect 4050 9820 4080 9910
rect 4130 9940 4210 9960
rect 4130 9900 4150 9940
rect 4190 9900 4210 9940
rect 4260 9930 4280 9970
rect 4320 9940 4340 9970
rect 4490 9940 4520 10040
rect 4880 9960 4910 10040
rect 5270 10010 5300 10040
rect 5560 10010 5590 10040
rect 4320 9930 4520 9940
rect 4260 9910 4520 9930
rect 4130 9880 4210 9900
rect 4490 9820 4520 9910
rect 4830 9940 4910 9960
rect 4830 9900 4850 9940
rect 4890 9900 4910 9940
rect 5220 9990 5980 10010
rect 5220 9950 5240 9990
rect 5280 9980 5980 9990
rect 5280 9950 5300 9980
rect 5220 9930 5300 9950
rect 4830 9880 4910 9900
rect 4880 9820 4910 9880
rect 5270 9820 5300 9930
rect 5350 9910 5430 9930
rect 5350 9870 5370 9910
rect 5410 9880 5430 9910
rect 5700 9910 5780 9930
rect 5700 9880 5720 9910
rect 5410 9870 5720 9880
rect 5760 9870 5780 9910
rect 5350 9850 5780 9870
rect 5560 9820 5590 9850
rect 5950 9820 5980 9980
rect 7550 9880 7630 9900
rect 7550 9840 7570 9880
rect 7610 9850 7630 9880
rect 10390 9880 10470 9900
rect 10390 9850 10410 9880
rect 7610 9840 7760 9850
rect 7550 9820 7760 9840
rect 2490 9490 2570 9510
rect 2490 9450 2510 9490
rect 2550 9450 2570 9490
rect 2490 9430 2570 9450
rect 7640 9790 7760 9820
rect 7860 9810 8640 9850
rect 7860 9790 7980 9810
rect 8080 9790 8200 9810
rect 8300 9790 8420 9810
rect 8520 9790 8640 9810
rect 8740 9790 8860 9820
rect 9160 9790 9280 9820
rect 9380 9810 10160 9850
rect 9380 9790 9500 9810
rect 9600 9790 9720 9810
rect 9820 9790 9940 9810
rect 10040 9790 10160 9810
rect 10260 9840 10410 9850
rect 10450 9840 10470 9880
rect 10260 9820 10470 9840
rect 10260 9790 10380 9820
rect 1340 9390 1370 9420
rect 1450 9390 1480 9420
rect 1860 9390 1890 9420
rect 1970 9390 2000 9420
rect 2240 9390 2270 9420
rect 2350 9390 2380 9420
rect 2760 9390 2790 9420
rect 2870 9390 2900 9420
rect 3280 9390 3310 9420
rect 3390 9390 3420 9420
rect 3720 9390 3750 9420
rect 4050 9390 4080 9420
rect 4490 9390 4520 9420
rect 4880 9390 4910 9420
rect 5270 9390 5300 9420
rect 5560 9390 5590 9420
rect 5950 9390 5980 9420
rect 3260 9370 3340 9390
rect 3260 9330 3280 9370
rect 3320 9330 3340 9370
rect 7640 9360 7760 9390
rect 7860 9370 7980 9390
rect 8080 9370 8200 9390
rect 8300 9370 8420 9390
rect 8520 9370 8640 9390
rect 7860 9340 8640 9370
rect 8740 9370 8860 9390
rect 9160 9370 9280 9390
rect 8740 9340 9280 9370
rect 9380 9360 9500 9390
rect 9600 9360 9720 9390
rect 9820 9360 9940 9390
rect 10040 9360 10160 9390
rect 10260 9360 10380 9390
rect 7860 9330 8230 9340
rect 3260 9320 3340 9330
rect 8210 9300 8230 9330
rect 8270 9330 8640 9340
rect 8270 9300 8290 9330
rect 8210 9280 8290 9300
rect 8970 9300 8990 9340
rect 9030 9300 9050 9340
rect 8970 9280 9050 9300
rect 9380 9330 10160 9360
rect 9380 9310 9460 9330
rect 9380 9270 9400 9310
rect 9440 9270 9460 9310
rect 9380 9250 9460 9270
rect 10080 9310 10160 9330
rect 10080 9270 10100 9310
rect 10140 9270 10160 9310
rect 10080 9250 10160 9270
rect 1710 9150 1790 9170
rect 1710 9110 1730 9150
rect 1770 9110 1790 9150
rect 1710 9090 1790 9110
rect 4830 9150 4910 9160
rect 4830 9110 4850 9150
rect 4890 9110 4910 9150
rect 4830 9090 4910 9110
rect 1340 9060 1370 9090
rect 1450 9060 1480 9090
rect 1860 9060 1890 9090
rect 1970 9060 2000 9090
rect 2240 9060 2270 9090
rect 2350 9060 2380 9090
rect 2760 9060 2790 9090
rect 2870 9060 2900 9090
rect 3270 9060 3300 9090
rect 3600 9060 3630 9090
rect 3930 9060 3960 9090
rect 4490 9060 4520 9090
rect 4880 9060 4910 9090
rect 5270 9060 5300 9090
rect 5560 9060 5590 9090
rect 1590 9030 1670 9050
rect 1590 8990 1610 9030
rect 1650 8990 1670 9030
rect 1590 8970 1670 8990
rect 1140 8570 1220 8590
rect 1140 8530 1160 8570
rect 1200 8540 1220 8570
rect 1340 8540 1370 8660
rect 1200 8530 1370 8540
rect 1140 8510 1370 8530
rect 1340 8440 1370 8510
rect 1450 8550 1480 8660
rect 1450 8530 1550 8550
rect 1450 8490 1490 8530
rect 1530 8490 1550 8530
rect 1450 8470 1550 8490
rect 1640 8510 1670 8970
rect 2490 9030 2570 9050
rect 2490 8990 2510 9030
rect 2550 8990 2570 9030
rect 2490 8970 2570 8990
rect 1860 8510 1890 8660
rect 1640 8480 1890 8510
rect 1450 8440 1480 8470
rect 1860 8440 1890 8480
rect 1970 8630 2000 8660
rect 1970 8610 2070 8630
rect 1970 8570 2010 8610
rect 2050 8570 2070 8610
rect 1970 8550 2070 8570
rect 1970 8440 2000 8550
rect 2240 8440 2270 8660
rect 2350 8550 2380 8660
rect 2350 8530 2450 8550
rect 2350 8490 2390 8530
rect 2430 8490 2450 8530
rect 2350 8470 2450 8490
rect 2540 8510 2570 8970
rect 9820 8810 9900 8830
rect 7790 8770 7870 8790
rect 7790 8740 7810 8770
rect 7660 8730 7810 8740
rect 7850 8740 7870 8770
rect 8330 8780 8410 8800
rect 8330 8740 8350 8780
rect 8390 8740 8410 8780
rect 9410 8780 9490 8800
rect 9410 8740 9430 8780
rect 9470 8740 9490 8780
rect 9820 8770 9840 8810
rect 9880 8770 9900 8810
rect 9820 8750 9900 8770
rect 10080 8810 10160 8830
rect 10080 8770 10100 8810
rect 10140 8770 10160 8810
rect 10080 8750 10160 8770
rect 7850 8730 8000 8740
rect 7440 8690 7560 8720
rect 7660 8710 8000 8730
rect 7660 8690 7780 8710
rect 7880 8690 8000 8710
rect 8100 8710 8640 8740
rect 8100 8690 8220 8710
rect 8520 8690 8640 8710
rect 8740 8710 9080 8740
rect 8740 8690 8860 8710
rect 8960 8690 9080 8710
rect 9180 8710 9720 8740
rect 9180 8690 9300 8710
rect 9600 8690 9720 8710
rect 9820 8720 10160 8750
rect 9820 8690 9940 8720
rect 10040 8690 10160 8720
rect 10260 8690 10380 8720
rect 2760 8510 2790 8660
rect 2540 8480 2790 8510
rect 2350 8440 2380 8470
rect 2760 8440 2790 8480
rect 2870 8600 2900 8660
rect 2870 8580 3220 8600
rect 2870 8570 3080 8580
rect 2870 8440 2900 8570
rect 3060 8540 3080 8570
rect 3120 8540 3160 8580
rect 3200 8540 3220 8580
rect 3060 8520 3220 8540
rect 3270 8570 3300 8660
rect 3470 8580 3550 8600
rect 3470 8570 3490 8580
rect 3270 8540 3490 8570
rect 3530 8540 3550 8580
rect 3270 8440 3300 8540
rect 3470 8520 3550 8540
rect 3600 8570 3630 8660
rect 3800 8580 3880 8600
rect 3800 8570 3820 8580
rect 3600 8540 3820 8570
rect 3860 8540 3880 8580
rect 3600 8440 3630 8540
rect 3800 8520 3880 8540
rect 3930 8570 3960 8660
rect 4090 8580 4170 8600
rect 4090 8570 4110 8580
rect 3930 8540 4110 8570
rect 4150 8540 4170 8580
rect 3930 8440 3960 8540
rect 4090 8520 4170 8540
rect 4240 8570 4320 8590
rect 4240 8530 4260 8570
rect 4300 8540 4320 8570
rect 4490 8540 4520 8660
rect 4880 8630 4910 8660
rect 5270 8620 5300 8660
rect 5560 8620 5590 8660
rect 4960 8600 5980 8620
rect 4960 8560 4980 8600
rect 5020 8590 5980 8600
rect 5020 8560 5040 8590
rect 4960 8540 5040 8560
rect 4300 8530 4520 8540
rect 4240 8510 4520 8530
rect 4490 8440 4520 8510
rect 4880 8440 4910 8470
rect 5270 8440 5300 8590
rect 5350 8520 5430 8530
rect 5350 8480 5370 8520
rect 5410 8490 5430 8520
rect 5410 8480 5590 8490
rect 5350 8460 5590 8480
rect 5560 8440 5590 8460
rect 5950 8440 5980 8590
rect 7440 8260 7560 8290
rect 7350 8240 7560 8260
rect 1340 8210 1370 8240
rect 1450 8210 1480 8240
rect 1860 8160 1890 8240
rect 1970 8210 2000 8240
rect 2240 8160 2270 8240
rect 2350 8210 2380 8240
rect 2760 8210 2790 8240
rect 2870 8210 2900 8240
rect 3270 8210 3300 8240
rect 3600 8210 3630 8240
rect 3930 8210 3960 8240
rect 4490 8210 4520 8240
rect 4880 8210 4910 8240
rect 5270 8210 5300 8240
rect 5560 8210 5590 8240
rect 5950 8210 5980 8240
rect 1860 8130 2270 8160
rect 4880 8190 4990 8210
rect 4880 8150 4930 8190
rect 4970 8150 4990 8190
rect 4880 8130 4990 8150
rect 5540 8190 5620 8210
rect 5540 8150 5560 8190
rect 5600 8150 5620 8190
rect 7350 8200 7370 8240
rect 7410 8230 7560 8240
rect 7660 8270 7780 8290
rect 7880 8270 8000 8290
rect 7660 8230 8000 8270
rect 8100 8260 8220 8290
rect 8520 8260 8640 8290
rect 8740 8270 8860 8290
rect 8960 8270 9080 8290
rect 7410 8200 7430 8230
rect 7350 8180 7430 8200
rect 7880 8210 8000 8230
rect 8740 8230 9080 8270
rect 9180 8260 9300 8290
rect 9600 8260 9720 8290
rect 9820 8270 9940 8290
rect 10040 8270 10160 8290
rect 9820 8230 10160 8270
rect 10260 8260 10380 8290
rect 10260 8240 10470 8260
rect 10260 8230 10410 8240
rect 8740 8210 8860 8230
rect 7880 8180 8860 8210
rect 10390 8200 10410 8230
rect 10450 8200 10470 8240
rect 10390 8180 10470 8200
rect 5540 8130 5620 8150
rect -360 6960 -280 6980
rect -360 6920 -340 6960
rect -300 6930 -280 6960
rect 960 6960 1040 6980
rect 960 6930 980 6960
rect -300 6920 -250 6930
rect -360 6900 -250 6920
rect 930 6920 980 6930
rect 1020 6920 1040 6960
rect 930 6900 1040 6920
rect 1540 6960 1620 6980
rect 1540 6920 1560 6960
rect 1600 6930 1620 6960
rect 2860 6960 2940 6980
rect 2860 6930 2880 6960
rect 1600 6920 1650 6930
rect 1540 6900 1650 6920
rect 2830 6920 2880 6930
rect 2920 6920 2940 6960
rect 2830 6900 2940 6920
rect -280 6870 -250 6900
rect -170 6870 -140 6900
rect -60 6870 -30 6900
rect 50 6870 80 6900
rect 160 6870 190 6900
rect 270 6870 300 6900
rect 380 6870 410 6900
rect 490 6870 520 6900
rect 600 6870 630 6900
rect 710 6870 740 6900
rect 820 6870 850 6900
rect 930 6870 960 6900
rect 1620 6870 1650 6900
rect 1730 6870 1760 6900
rect 1840 6870 1870 6900
rect 1950 6870 1980 6900
rect 2060 6870 2090 6900
rect 2170 6870 2200 6900
rect 2280 6870 2310 6900
rect 2390 6870 2420 6900
rect 2500 6870 2530 6900
rect 2610 6870 2640 6900
rect 2720 6870 2750 6900
rect 2830 6870 2860 6900
rect -280 6640 -250 6670
rect -170 6640 -140 6670
rect -60 6640 -30 6670
rect 50 6640 80 6670
rect 160 6640 190 6670
rect 270 6640 300 6670
rect 380 6640 410 6670
rect 490 6640 520 6670
rect 600 6640 630 6670
rect 710 6640 740 6670
rect 820 6640 850 6670
rect 930 6640 960 6670
rect 1620 6640 1650 6670
rect 1730 6640 1760 6670
rect 1840 6640 1870 6670
rect 1950 6640 1980 6670
rect 2060 6640 2090 6670
rect 2170 6640 2200 6670
rect 2280 6640 2310 6670
rect 2390 6640 2420 6670
rect 2500 6640 2530 6670
rect 2610 6640 2640 6670
rect 2720 6640 2750 6670
rect 2830 6640 2860 6670
rect -184 6622 -126 6640
rect -184 6588 -172 6622
rect -138 6588 -126 6622
rect -184 6570 -126 6588
rect -74 6622 -16 6640
rect -74 6588 -62 6622
rect -28 6588 -16 6622
rect -74 6570 -16 6588
rect 36 6622 94 6640
rect 36 6588 48 6622
rect 82 6588 94 6622
rect 36 6570 94 6588
rect 146 6622 204 6640
rect 146 6588 158 6622
rect 192 6588 204 6622
rect 146 6570 204 6588
rect 256 6622 314 6640
rect 256 6588 268 6622
rect 302 6588 314 6622
rect 256 6570 314 6588
rect 366 6622 424 6640
rect 366 6588 378 6622
rect 412 6588 424 6622
rect 366 6570 424 6588
rect 476 6622 534 6640
rect 476 6588 488 6622
rect 522 6588 534 6622
rect 476 6570 534 6588
rect 586 6622 644 6640
rect 586 6588 598 6622
rect 632 6588 644 6622
rect 586 6570 644 6588
rect 696 6622 754 6640
rect 696 6588 708 6622
rect 742 6588 754 6622
rect 696 6570 754 6588
rect 806 6622 864 6640
rect 806 6588 818 6622
rect 852 6588 864 6622
rect 806 6570 864 6588
rect 1716 6622 1774 6640
rect 1716 6588 1728 6622
rect 1762 6588 1774 6622
rect 1716 6570 1774 6588
rect 1826 6622 1884 6640
rect 1826 6588 1838 6622
rect 1872 6588 1884 6622
rect 1826 6570 1884 6588
rect 1936 6622 1994 6640
rect 1936 6588 1948 6622
rect 1982 6588 1994 6622
rect 1936 6570 1994 6588
rect 2046 6622 2104 6640
rect 2046 6588 2058 6622
rect 2092 6588 2104 6622
rect 2046 6570 2104 6588
rect 2156 6622 2214 6640
rect 2156 6588 2168 6622
rect 2202 6588 2214 6622
rect 2156 6570 2214 6588
rect 2266 6622 2324 6640
rect 2266 6588 2278 6622
rect 2312 6588 2324 6622
rect 2266 6570 2324 6588
rect 2376 6622 2434 6640
rect 2376 6588 2388 6622
rect 2422 6588 2434 6622
rect 2376 6570 2434 6588
rect 2486 6622 2544 6640
rect 2486 6588 2498 6622
rect 2532 6588 2544 6622
rect 2486 6570 2544 6588
rect 2596 6622 2654 6640
rect 2596 6588 2608 6622
rect 2642 6588 2654 6622
rect 2596 6570 2654 6588
rect 2706 6622 2764 6640
rect 2706 6588 2718 6622
rect 2752 6588 2764 6622
rect 2706 6570 2764 6588
rect -370 6360 -290 6380
rect -370 6320 -350 6360
rect -310 6330 -290 6360
rect 2870 6360 2950 6380
rect 2870 6330 2890 6360
rect -310 6320 -190 6330
rect -370 6300 -190 6320
rect 2770 6320 2890 6330
rect 2930 6320 2950 6360
rect 2770 6300 2950 6320
rect 7254 6340 7684 6356
rect 7254 6306 7270 6340
rect 7304 6306 7684 6340
rect -290 6270 -190 6300
rect -110 6270 -10 6300
rect 70 6270 170 6300
rect 250 6270 350 6300
rect 430 6270 530 6300
rect 610 6270 710 6300
rect 790 6270 890 6300
rect 970 6270 1070 6300
rect 1150 6270 1250 6300
rect 1330 6270 1430 6300
rect 1510 6270 1610 6300
rect 1690 6270 1790 6300
rect 1870 6270 1970 6300
rect 2050 6270 2150 6300
rect 2230 6270 2330 6300
rect 2410 6270 2510 6300
rect 2590 6270 2690 6300
rect 2770 6270 2870 6300
rect 7254 6290 7684 6306
rect 8164 6340 8594 6356
rect 8164 6306 8544 6340
rect 8578 6306 8594 6340
rect 8164 6290 8594 6306
rect 3510 6160 3570 6180
rect 3510 6120 3520 6160
rect 3560 6120 3570 6160
rect 3950 6160 4010 6180
rect 3950 6120 3960 6160
rect 4000 6120 4010 6160
rect 3510 6090 3610 6120
rect 3580 6070 3610 6090
rect 3690 6070 3720 6100
rect 3800 6070 3830 6100
rect 3910 6090 4010 6120
rect 8210 6150 8290 6170
rect 8210 6110 8230 6150
rect 8270 6110 8290 6150
rect 8610 6150 8690 6170
rect 8610 6110 8630 6150
rect 8670 6110 8690 6150
rect 3910 6070 3940 6090
rect 7500 6060 7600 6090
rect 7700 6080 9200 6110
rect 7700 6060 7800 6080
rect 7900 6060 8000 6080
rect 8100 6060 8200 6080
rect 8300 6060 8400 6080
rect 8500 6060 8600 6080
rect 8700 6060 8800 6080
rect 8900 6060 9000 6080
rect 9100 6060 9200 6080
rect 9300 6060 9400 6090
rect 3580 5840 3610 5870
rect 3690 5850 3720 5870
rect 3800 5850 3830 5870
rect 3690 5820 3830 5850
rect 3910 5840 3940 5870
rect 3720 5780 3740 5820
rect 3780 5780 3800 5820
rect 7500 5780 7600 5810
rect 7700 5780 7800 5810
rect 7900 5780 8000 5810
rect 8100 5780 8200 5810
rect 8300 5780 8400 5810
rect 8500 5780 8600 5810
rect 8700 5780 8800 5810
rect 8900 5780 9000 5810
rect 9100 5780 9200 5810
rect 9300 5780 9400 5810
rect 3720 5760 3800 5780
rect 7410 5760 7600 5780
rect 7410 5720 7430 5760
rect 7470 5750 7600 5760
rect 9300 5760 9490 5780
rect 9300 5750 9430 5760
rect 7470 5720 7490 5750
rect 7410 5700 7490 5720
rect 9410 5720 9430 5750
rect 9470 5720 9490 5760
rect 9410 5700 9490 5720
rect -290 5640 -190 5670
rect -110 5640 -10 5670
rect 70 5640 170 5670
rect 250 5640 350 5670
rect 430 5640 530 5670
rect 610 5640 710 5670
rect 790 5640 890 5670
rect 970 5640 1070 5670
rect 1150 5640 1250 5670
rect 1330 5640 1430 5670
rect 1510 5640 1610 5670
rect 1690 5640 1790 5670
rect 1870 5640 1970 5670
rect 2050 5640 2150 5670
rect 2230 5640 2330 5670
rect 2410 5640 2510 5670
rect -90 5620 -20 5640
rect -90 5580 -80 5620
rect -40 5580 -20 5620
rect -90 5560 -20 5580
rect 80 5620 160 5640
rect 80 5580 100 5620
rect 140 5580 160 5620
rect 80 5560 160 5580
rect 260 5620 340 5640
rect 260 5580 280 5620
rect 320 5580 340 5620
rect 260 5560 340 5580
rect 440 5620 520 5640
rect 440 5580 460 5620
rect 500 5580 520 5620
rect 440 5560 520 5580
rect 620 5620 700 5640
rect 620 5580 640 5620
rect 680 5580 700 5620
rect 620 5560 700 5580
rect 800 5620 880 5640
rect 800 5580 820 5620
rect 860 5580 880 5620
rect 800 5560 880 5580
rect 980 5620 1060 5640
rect 980 5580 1000 5620
rect 1040 5580 1060 5620
rect 980 5560 1060 5580
rect 1160 5620 1230 5640
rect 1160 5580 1180 5620
rect 1220 5580 1230 5620
rect 1160 5560 1230 5580
rect 1350 5620 1420 5640
rect 1350 5580 1360 5620
rect 1400 5580 1420 5620
rect 1350 5560 1420 5580
rect 1520 5620 1600 5640
rect 1520 5580 1540 5620
rect 1580 5580 1600 5620
rect 1520 5560 1600 5580
rect 1700 5620 1780 5640
rect 1700 5580 1720 5620
rect 1760 5580 1780 5620
rect 1700 5560 1780 5580
rect 1880 5620 1960 5640
rect 1880 5580 1900 5620
rect 1940 5580 1960 5620
rect 1880 5560 1960 5580
rect 2060 5620 2140 5640
rect 2060 5580 2080 5620
rect 2120 5580 2140 5620
rect 2060 5560 2140 5580
rect 2240 5620 2320 5640
rect 2240 5580 2260 5620
rect 2300 5580 2320 5620
rect 2240 5560 2320 5580
rect 2420 5620 2500 5640
rect 2590 5630 2690 5670
rect 2770 5640 2870 5670
rect 2420 5580 2440 5620
rect 2480 5580 2500 5620
rect 2420 5560 2500 5580
rect 2600 5620 2670 5630
rect 2600 5580 2620 5620
rect 2660 5580 2670 5620
rect 2600 5560 2670 5580
rect 7520 5470 7610 5490
rect 7520 5420 7540 5470
rect 7590 5420 7610 5470
rect 7520 5400 7610 5420
rect 8170 5470 8260 5490
rect 8170 5420 8190 5470
rect 8240 5420 8260 5470
rect 8170 5400 8260 5420
rect 8660 5460 8740 5480
rect 8660 5420 8680 5460
rect 8720 5420 8740 5460
rect 8660 5400 8740 5420
rect 9320 5460 9400 5480
rect 9320 5420 9340 5460
rect 9380 5420 9400 5460
rect 9320 5400 9400 5420
rect 9800 5460 9880 5480
rect 9800 5420 9820 5460
rect 9860 5420 9880 5460
rect 9800 5400 9880 5420
rect 10460 5460 10540 5480
rect 10460 5420 10480 5460
rect 10520 5420 10540 5460
rect 10460 5400 10540 5420
rect 7550 5370 7580 5400
rect 7680 5370 7710 5400
rect 7810 5370 7840 5400
rect 7940 5370 7970 5400
rect 8070 5370 8100 5400
rect 8200 5370 8230 5400
rect 8690 5370 8720 5400
rect 8820 5370 8850 5400
rect 8950 5370 8980 5400
rect 9080 5370 9110 5400
rect 9210 5370 9240 5400
rect 9340 5370 9370 5400
rect 9830 5370 9860 5400
rect 9960 5370 9990 5400
rect 10090 5370 10120 5400
rect 10220 5370 10250 5400
rect 10350 5370 10380 5400
rect 10480 5370 10510 5400
rect 7550 5240 7580 5270
rect 7680 5250 7710 5270
rect 7810 5250 7840 5270
rect 7940 5250 7970 5270
rect 8070 5250 8100 5270
rect 7680 5220 8100 5250
rect 8200 5240 8230 5270
rect 8690 5240 8720 5270
rect 8820 5250 8850 5270
rect 8950 5250 8980 5270
rect 8820 5240 8980 5250
rect 8770 5220 8980 5240
rect 9080 5250 9110 5270
rect 9210 5250 9240 5270
rect 9080 5240 9240 5250
rect 9340 5240 9370 5270
rect 9830 5240 9860 5270
rect 9080 5220 9290 5240
rect 7720 5180 7740 5220
rect 7780 5180 7800 5220
rect 7720 5160 7800 5180
rect 8770 5180 8790 5220
rect 8830 5180 8850 5220
rect 8770 5160 8850 5180
rect 9210 5180 9230 5220
rect 9270 5180 9290 5220
rect 9210 5160 9290 5180
rect 9960 5190 9990 5270
rect 10090 5190 10120 5270
rect 10220 5190 10250 5270
rect 10350 5190 10380 5270
rect 10480 5240 10510 5270
rect 10750 5220 10830 5240
rect 10750 5190 10770 5220
rect 9960 5180 10770 5190
rect 10810 5180 10830 5220
rect 9960 5160 10830 5180
rect 9960 5120 9990 5160
rect 9910 5100 9990 5120
rect 9910 5060 9930 5100
rect 9970 5060 9990 5100
rect 9910 5040 9990 5060
rect 7630 4880 7710 4900
rect 7630 4840 7650 4880
rect 7690 4840 7710 4880
rect 8070 4880 8150 4900
rect 8070 4840 8090 4880
rect 8130 4840 8150 4880
rect 8860 4890 8940 4910
rect 8860 4850 8880 4890
rect 8920 4850 8940 4890
rect 8860 4840 8940 4850
rect 9910 4880 10830 4900
rect 9910 4840 9930 4880
rect 9970 4870 10770 4880
rect 9970 4840 9990 4870
rect 7630 4820 7840 4840
rect -1460 4800 -1400 4820
rect -1460 4760 -1450 4800
rect -1410 4770 -1400 4800
rect 940 4800 1000 4820
rect 940 4770 950 4800
rect -1410 4760 -1350 4770
rect -1460 4740 -1350 4760
rect 890 4760 950 4770
rect 990 4760 1000 4800
rect 890 4740 1000 4760
rect 1580 4800 1640 4820
rect 1580 4760 1590 4800
rect 1630 4770 1640 4800
rect 3980 4800 4040 4820
rect 3980 4770 3990 4800
rect 1630 4760 1690 4770
rect 1580 4740 1690 4760
rect 3930 4760 3990 4770
rect 4030 4760 4040 4800
rect 7550 4790 7580 4820
rect 7680 4810 7840 4820
rect 7680 4790 7710 4810
rect 7810 4790 7840 4810
rect 7940 4820 8150 4840
rect 7940 4810 8100 4820
rect 7940 4790 7970 4810
rect 8070 4790 8100 4810
rect 8200 4790 8230 4820
rect 8690 4790 8720 4820
rect 8820 4810 9240 4840
rect 9910 4820 9990 4840
rect 8820 4790 8850 4810
rect 8950 4790 8980 4810
rect 9080 4790 9110 4810
rect 9210 4790 9240 4810
rect 9340 4790 9370 4820
rect 9830 4790 9860 4820
rect 9960 4790 9990 4820
rect 10090 4790 10120 4870
rect 10220 4790 10250 4870
rect 10350 4790 10380 4870
rect 10750 4840 10770 4870
rect 10810 4840 10830 4880
rect 10750 4820 10830 4840
rect 10480 4790 10510 4820
rect 3930 4740 4040 4760
rect -1390 4710 -1350 4740
rect -1270 4710 -1230 4740
rect -1150 4710 -1110 4740
rect -1030 4710 -990 4740
rect -910 4710 -870 4740
rect -790 4710 -750 4740
rect -670 4710 -630 4740
rect -550 4710 -510 4740
rect -430 4710 -390 4740
rect -310 4710 -270 4740
rect -190 4710 -150 4740
rect -70 4710 -30 4740
rect 50 4710 90 4740
rect 170 4710 210 4740
rect 290 4710 330 4740
rect 410 4710 450 4740
rect 530 4710 570 4740
rect 650 4710 690 4740
rect 770 4710 810 4740
rect 890 4710 930 4740
rect 1650 4710 1690 4740
rect 1770 4710 1810 4740
rect 1890 4710 1930 4740
rect 2010 4710 2050 4740
rect 2130 4710 2170 4740
rect 2250 4710 2290 4740
rect 2370 4710 2410 4740
rect 2490 4710 2530 4740
rect 2610 4710 2650 4740
rect 2730 4710 2770 4740
rect 2850 4710 2890 4740
rect 2970 4710 3010 4740
rect 3090 4710 3130 4740
rect 3210 4710 3250 4740
rect 3330 4710 3370 4740
rect 3450 4710 3490 4740
rect 3570 4710 3610 4740
rect 3690 4710 3730 4740
rect 3810 4710 3850 4740
rect 3930 4710 3970 4740
rect 7550 4560 7580 4590
rect 7680 4560 7710 4590
rect 7810 4560 7840 4590
rect 7940 4560 7970 4590
rect 8070 4560 8100 4590
rect 8200 4560 8230 4590
rect 8690 4560 8720 4590
rect 8820 4560 8850 4590
rect 8950 4560 8980 4590
rect 9080 4560 9110 4590
rect 9210 4560 9240 4590
rect 9340 4560 9370 4590
rect 9830 4560 9860 4590
rect 9960 4560 9990 4590
rect 10090 4560 10120 4590
rect 10220 4560 10250 4590
rect 10350 4560 10380 4590
rect 10480 4560 10510 4590
rect 7520 4540 7600 4560
rect -1390 4480 -1350 4510
rect -1270 4470 -1230 4510
rect -1150 4490 -1110 4510
rect -1030 4490 -990 4510
rect -910 4490 -870 4510
rect -790 4490 -750 4510
rect -1280 4450 -1220 4470
rect -1150 4460 -750 4490
rect -670 4490 -630 4510
rect -550 4490 -510 4510
rect -670 4460 -510 4490
rect -430 4490 -390 4510
rect -310 4490 -270 4510
rect -190 4490 -150 4510
rect -70 4490 -30 4510
rect -430 4460 -30 4490
rect 50 4490 90 4510
rect 170 4490 210 4510
rect 50 4460 210 4490
rect 290 4490 330 4510
rect 410 4490 450 4510
rect 530 4490 570 4510
rect 650 4490 690 4510
rect 290 4460 690 4490
rect 770 4480 810 4510
rect 890 4480 930 4510
rect 1650 4480 1690 4510
rect 1770 4480 1810 4510
rect 1890 4490 1930 4510
rect 2010 4490 2050 4510
rect 2130 4490 2170 4510
rect 2250 4490 2290 4510
rect 760 4460 820 4480
rect -1280 4410 -1270 4450
rect -1230 4410 -1220 4450
rect -1280 4390 -1220 4410
rect -1110 4420 -1090 4460
rect -1050 4420 -1030 4460
rect -1110 4400 -1030 4420
rect -620 4420 -610 4460
rect -570 4420 -560 4460
rect -620 4400 -560 4420
rect -390 4420 -370 4460
rect -330 4420 -310 4460
rect -390 4400 -310 4420
rect 100 4420 110 4460
rect 150 4420 160 4460
rect 100 4400 160 4420
rect 330 4420 350 4460
rect 390 4420 410 4460
rect 330 4400 410 4420
rect 760 4420 770 4460
rect 810 4420 820 4460
rect 760 4400 820 4420
rect 1760 4460 1820 4480
rect 1890 4460 2290 4490
rect 2370 4490 2410 4510
rect 2490 4490 2530 4510
rect 2370 4460 2530 4490
rect 2610 4490 2650 4510
rect 2730 4490 2770 4510
rect 2850 4490 2890 4510
rect 2970 4490 3010 4510
rect 2610 4460 3010 4490
rect 3090 4490 3130 4510
rect 3210 4490 3250 4510
rect 3090 4460 3250 4490
rect 3330 4490 3370 4510
rect 3450 4490 3490 4510
rect 3570 4490 3610 4510
rect 3690 4490 3730 4510
rect 3330 4460 3730 4490
rect 3810 4470 3850 4510
rect 3930 4480 3970 4510
rect 7520 4500 7540 4540
rect 7580 4500 7600 4540
rect 7520 4480 7600 4500
rect 8180 4540 8260 4560
rect 8180 4500 8200 4540
rect 8240 4500 8260 4540
rect 8180 4480 8260 4500
rect 8660 4540 8740 4560
rect 8660 4500 8680 4540
rect 8720 4500 8740 4540
rect 8660 4480 8740 4500
rect 9320 4540 9400 4560
rect 9320 4500 9340 4540
rect 9380 4500 9400 4540
rect 9320 4480 9400 4500
rect 9800 4540 9880 4560
rect 9800 4500 9820 4540
rect 9860 4500 9880 4540
rect 9800 4480 9880 4500
rect 10460 4540 10540 4560
rect 10460 4500 10480 4540
rect 10520 4500 10540 4540
rect 10460 4480 10540 4500
rect 1760 4420 1770 4460
rect 1810 4420 1820 4460
rect 1760 4400 1820 4420
rect 2170 4420 2190 4460
rect 2230 4420 2250 4460
rect 2170 4400 2250 4420
rect 2420 4420 2430 4460
rect 2470 4420 2480 4460
rect 2420 4400 2480 4420
rect 2890 4420 2910 4460
rect 2950 4420 2970 4460
rect 2890 4400 2970 4420
rect 3140 4420 3150 4460
rect 3190 4420 3200 4460
rect 3140 4400 3200 4420
rect 3610 4420 3630 4460
rect 3670 4420 3690 4460
rect 3610 4400 3690 4420
rect 3800 4450 3860 4470
rect 3800 4410 3810 4450
rect 3850 4410 3860 4450
rect 3800 4390 3860 4410
rect 7530 4230 7610 4250
rect 7530 4190 7550 4230
rect 7590 4200 7610 4230
rect 9530 4230 9610 4250
rect 9530 4200 9550 4230
rect 7590 4190 7720 4200
rect 7530 4170 7720 4190
rect 9420 4190 9550 4200
rect 9590 4190 9610 4230
rect 9420 4170 9610 4190
rect 7620 4140 7720 4170
rect 7820 4140 7920 4170
rect 8020 4140 8120 4170
rect 8220 4140 8320 4170
rect 8420 4140 8520 4170
rect 8620 4140 8720 4170
rect 8820 4140 8920 4170
rect 9020 4140 9120 4170
rect 9220 4140 9320 4170
rect 9420 4140 9520 4170
rect -458 3852 -390 3870
rect -458 3818 -446 3852
rect -412 3818 -390 3852
rect -458 3800 -390 3818
rect -550 3770 -510 3800
rect -430 3770 -390 3800
rect -310 3852 -242 3870
rect -310 3818 -288 3852
rect -254 3818 -242 3852
rect -310 3800 -242 3818
rect 24 3852 90 3870
rect 24 3818 36 3852
rect 70 3818 90 3852
rect 24 3800 90 3818
rect -310 3770 -270 3800
rect -190 3770 -150 3800
rect -70 3770 -30 3800
rect 50 3770 90 3800
rect 170 3852 236 3870
rect 170 3818 190 3852
rect 224 3818 236 3852
rect 170 3800 236 3818
rect 502 3852 570 3870
rect 502 3818 514 3852
rect 548 3818 570 3852
rect 2010 3852 2078 3870
rect 502 3800 570 3818
rect 170 3770 210 3800
rect 290 3770 330 3800
rect 410 3770 450 3800
rect 530 3770 570 3800
rect -550 3640 -510 3670
rect -430 3640 -390 3670
rect -310 3640 -270 3670
rect -190 3640 -150 3670
rect -70 3640 -30 3670
rect 50 3640 90 3670
rect 170 3640 210 3670
rect 290 3640 330 3670
rect 410 3640 450 3670
rect 530 3640 570 3670
rect -559 3622 -501 3640
rect -559 3588 -547 3622
rect -513 3588 -501 3622
rect -559 3570 -501 3588
rect -199 3622 -141 3640
rect -199 3588 -187 3622
rect -153 3588 -141 3622
rect -199 3570 -141 3588
rect -79 3622 -21 3640
rect -79 3588 -67 3622
rect -33 3588 -21 3622
rect -79 3570 -21 3588
rect 281 3622 339 3640
rect 281 3588 293 3622
rect 327 3588 339 3622
rect 281 3570 339 3588
rect 401 3622 459 3640
rect 401 3588 413 3622
rect 447 3588 459 3622
rect 401 3570 459 3588
rect 2010 3818 2032 3852
rect 2066 3818 2078 3852
rect 2010 3800 2078 3818
rect 2344 3852 2410 3870
rect 2344 3818 2356 3852
rect 2390 3818 2410 3852
rect 2344 3800 2410 3818
rect 2010 3770 2050 3800
rect 2130 3770 2170 3800
rect 2250 3770 2290 3800
rect 2370 3770 2410 3800
rect 2490 3852 2556 3870
rect 2490 3818 2510 3852
rect 2544 3818 2556 3852
rect 2490 3800 2556 3818
rect 2822 3852 2890 3870
rect 2822 3818 2834 3852
rect 2868 3818 2890 3852
rect 2822 3800 2890 3818
rect 2490 3770 2530 3800
rect 2610 3770 2650 3800
rect 2730 3770 2770 3800
rect 2850 3770 2890 3800
rect 2970 3852 3038 3870
rect 2970 3818 2992 3852
rect 3026 3818 3038 3852
rect 2970 3800 3038 3818
rect 2970 3770 3010 3800
rect 3090 3770 3130 3800
rect 2010 3640 2050 3670
rect 2130 3640 2170 3670
rect 2250 3640 2290 3670
rect 2370 3640 2410 3670
rect 2490 3640 2530 3670
rect 2610 3640 2650 3670
rect 2730 3640 2770 3670
rect 2850 3640 2890 3670
rect 2970 3640 3010 3670
rect 3090 3640 3130 3670
rect 2121 3622 2179 3640
rect 2121 3588 2133 3622
rect 2167 3588 2179 3622
rect 2121 3570 2179 3588
rect 2241 3622 2299 3640
rect 2241 3588 2253 3622
rect 2287 3588 2299 3622
rect 2241 3570 2299 3588
rect 2601 3622 2659 3640
rect 2601 3588 2613 3622
rect 2647 3588 2659 3622
rect 2601 3570 2659 3588
rect 2721 3622 2779 3640
rect 2721 3588 2733 3622
rect 2767 3588 2779 3622
rect 2721 3570 2779 3588
rect 3081 3622 3139 3640
rect 3081 3588 3093 3622
rect 3127 3588 3139 3622
rect 7620 3610 7720 3640
rect 7820 3620 7920 3640
rect 8020 3620 8120 3640
rect 8220 3620 8320 3640
rect 8420 3620 8520 3640
rect 8620 3620 8720 3640
rect 8820 3620 8920 3640
rect 9020 3620 9120 3640
rect 9220 3620 9320 3640
rect 7820 3590 9320 3620
rect 9420 3610 9520 3640
rect 3081 3570 3139 3588
rect 8330 3550 8350 3590
rect 8390 3550 8410 3590
rect 8330 3530 8410 3550
rect 8730 3550 8750 3590
rect 8790 3550 8810 3590
rect 8730 3530 8810 3550
rect -1070 3250 -990 3270
rect -1070 3210 -1050 3250
rect -1010 3210 -990 3250
rect -1070 3190 -990 3210
rect -830 3250 -750 3270
rect -830 3210 -810 3250
rect -770 3210 -750 3250
rect -830 3190 -750 3210
rect -590 3250 -510 3270
rect -590 3210 -570 3250
rect -530 3210 -510 3250
rect -590 3190 -510 3210
rect -350 3250 -270 3270
rect -350 3210 -330 3250
rect -290 3210 -270 3250
rect -350 3190 -270 3210
rect 290 3250 370 3270
rect 290 3210 310 3250
rect 350 3210 370 3250
rect 290 3190 370 3210
rect 530 3250 610 3270
rect 530 3210 550 3250
rect 590 3210 610 3250
rect 530 3190 610 3210
rect 770 3250 850 3270
rect 770 3210 790 3250
rect 830 3210 850 3250
rect 770 3190 850 3210
rect 1730 3250 1810 3270
rect 1730 3210 1750 3250
rect 1790 3210 1810 3250
rect 1730 3190 1810 3210
rect 1970 3250 2050 3270
rect 1970 3210 1990 3250
rect 2030 3210 2050 3250
rect 1970 3190 2050 3210
rect 2210 3250 2290 3270
rect 2210 3210 2230 3250
rect 2270 3210 2290 3250
rect 2210 3190 2290 3210
rect 2850 3250 2930 3270
rect 2850 3210 2870 3250
rect 2910 3210 2930 3250
rect 2850 3190 2930 3210
rect 3090 3250 3170 3270
rect 3090 3210 3110 3250
rect 3150 3210 3170 3250
rect 3090 3190 3170 3210
rect 3330 3250 3410 3270
rect 3330 3210 3350 3250
rect 3390 3210 3410 3250
rect 3330 3190 3410 3210
rect 3570 3250 3650 3270
rect 3570 3210 3590 3250
rect 3630 3210 3650 3250
rect 3570 3190 3650 3210
rect -1170 3160 -170 3190
rect 70 3160 1070 3190
rect 1510 3160 2510 3190
rect 2750 3160 3750 3190
rect -1170 2630 -170 2660
rect 70 2630 1070 2660
rect 1510 2630 2510 2660
rect 2750 2630 3750 2660
rect -670 2340 -590 2360
rect -670 2300 -650 2340
rect -610 2300 -590 2340
rect -670 2280 -590 2300
rect -510 2340 -430 2360
rect -510 2300 -490 2340
rect -450 2300 -430 2340
rect -510 2280 -430 2300
rect -350 2340 -270 2360
rect -350 2300 -330 2340
rect -290 2300 -270 2340
rect -350 2280 -270 2300
rect -190 2340 -110 2360
rect -190 2300 -170 2340
rect -130 2300 -110 2340
rect -190 2280 -110 2300
rect -30 2340 50 2360
rect -30 2300 -10 2340
rect 30 2300 50 2340
rect -30 2280 50 2300
rect 130 2340 210 2360
rect 130 2300 150 2340
rect 190 2300 210 2340
rect 130 2280 210 2300
rect 290 2340 370 2360
rect 290 2300 310 2340
rect 350 2300 370 2340
rect 290 2280 370 2300
rect 450 2340 530 2360
rect 450 2300 470 2340
rect 510 2300 530 2340
rect 450 2280 530 2300
rect 610 2340 690 2360
rect 610 2300 630 2340
rect 670 2300 690 2340
rect 610 2280 690 2300
rect 770 2340 850 2360
rect 770 2300 790 2340
rect 830 2300 850 2340
rect 770 2280 850 2300
rect 930 2340 1010 2360
rect 930 2300 950 2340
rect 990 2300 1010 2340
rect 930 2280 1010 2300
rect 1090 2340 1170 2360
rect 1090 2300 1110 2340
rect 1150 2300 1170 2340
rect 1090 2280 1170 2300
rect 1410 2340 1490 2360
rect 1410 2300 1430 2340
rect 1470 2300 1490 2340
rect 1410 2280 1490 2300
rect 1570 2340 1650 2360
rect 1570 2300 1590 2340
rect 1630 2300 1650 2340
rect 1570 2280 1650 2300
rect 1730 2340 1810 2360
rect 1730 2300 1750 2340
rect 1790 2300 1810 2340
rect 1730 2280 1810 2300
rect 1890 2340 1970 2360
rect 1890 2300 1910 2340
rect 1950 2300 1970 2340
rect 1890 2280 1970 2300
rect 2050 2340 2130 2360
rect 2050 2300 2070 2340
rect 2110 2300 2130 2340
rect 2050 2280 2130 2300
rect 2210 2340 2290 2360
rect 2210 2300 2230 2340
rect 2270 2300 2290 2340
rect 2210 2280 2290 2300
rect 2370 2340 2450 2360
rect 2370 2300 2390 2340
rect 2430 2300 2450 2340
rect 2370 2280 2450 2300
rect 2530 2340 2610 2360
rect 2530 2300 2550 2340
rect 2590 2300 2610 2340
rect 2530 2280 2610 2300
rect 2690 2340 2770 2360
rect 2690 2300 2710 2340
rect 2750 2300 2770 2340
rect 2690 2280 2770 2300
rect 2850 2340 2930 2360
rect 2850 2300 2870 2340
rect 2910 2300 2930 2340
rect 2850 2280 2930 2300
rect 3010 2340 3090 2360
rect 3010 2300 3030 2340
rect 3070 2300 3090 2340
rect 3010 2280 3090 2300
rect 3170 2340 3250 2360
rect 3170 2300 3190 2340
rect 3230 2300 3250 2340
rect 3170 2280 3250 2300
rect -750 2250 1250 2280
rect 1330 2250 3330 2280
rect -750 2020 1250 2050
rect 1330 2020 3330 2050
<< polycont >>
rect 11288 14068 11322 14102
rect 11808 14068 11842 14102
rect 12328 14068 12362 14102
rect 12896 14068 12930 14102
rect 410 13270 450 13310
rect 1360 13250 1400 13290
rect 2430 13260 2470 13300
rect 3990 13260 4030 13300
rect 6594 13270 6634 13310
rect 520 13030 560 13070
rect 1100 13030 1140 13070
rect 7150 13120 7190 13160
rect 1440 13030 1480 13070
rect 390 12830 430 12870
rect 1640 12950 1680 12990
rect 2020 13030 2060 13070
rect 2040 12910 2080 12950
rect 2540 13030 2580 13070
rect 2890 13030 2930 13070
rect 3470 13030 3510 13070
rect 3680 13030 3720 13070
rect 3920 13030 3960 13070
rect 4260 13020 4300 13060
rect 4530 12980 4570 13020
rect 3740 12910 3780 12950
rect 4730 12950 4770 12990
rect 5160 13030 5200 13070
rect 5130 12910 5170 12950
rect 5520 13030 5560 13070
rect 5850 13030 5890 13070
rect 6430 13030 6470 13070
rect 6260 12950 6300 12990
rect 6900 13010 6940 13050
rect 7730 13120 7770 13160
rect 8450 13120 8490 13160
rect 8200 13010 8240 13050
rect 7560 12950 7600 12990
rect 9030 13120 9070 13160
rect 9750 13120 9790 13160
rect 9500 13010 9540 13050
rect 8860 12950 8900 12990
rect 10330 13120 10370 13160
rect 11302 13588 11336 13622
rect 11822 13588 11856 13622
rect 12342 13588 12376 13622
rect 11274 13208 11308 13242
rect 11794 13208 11828 13242
rect 12314 13208 12348 13242
rect 10160 12950 10200 12990
rect 10774 13008 10808 13042
rect 5720 12830 5760 12870
rect 1050 12710 1090 12750
rect 1360 12730 1400 12770
rect 2170 12710 2210 12750
rect 2300 12710 2340 12750
rect 3430 12710 3470 12750
rect 5190 12700 5230 12740
rect 7720 12710 7760 12750
rect 9020 12710 9060 12750
rect 10320 12710 10360 12750
rect 11274 12818 11308 12852
rect 11794 12818 11828 12852
rect 12314 12818 12348 12852
rect 11302 12238 11336 12272
rect 11822 12238 11856 12272
rect 12342 12238 12376 12272
rect 11420 11350 11460 11390
rect 11940 11350 11980 11390
rect 12460 11350 12500 11390
rect 12980 11350 13020 11390
rect 3410 10290 3450 10330
rect 1160 9910 1200 9950
rect 1490 9950 1530 9990
rect 2010 9870 2050 9910
rect 2390 9950 2430 9990
rect 1610 9450 1650 9490
rect 3060 9940 3100 9980
rect 3490 9900 3530 9940
rect 3820 9900 3860 9940
rect 4150 9900 4190 9940
rect 4280 9930 4320 9970
rect 4850 9900 4890 9940
rect 5240 9950 5280 9990
rect 5370 9870 5410 9910
rect 5720 9870 5760 9910
rect 7570 9840 7610 9880
rect 2510 9450 2550 9490
rect 10410 9840 10450 9880
rect 3280 9330 3320 9370
rect 8230 9300 8270 9340
rect 8990 9300 9030 9340
rect 9400 9270 9440 9310
rect 10100 9270 10140 9310
rect 1730 9110 1770 9150
rect 4850 9110 4890 9150
rect 1610 8990 1650 9030
rect 1160 8530 1200 8570
rect 1490 8490 1530 8530
rect 2510 8990 2550 9030
rect 2010 8570 2050 8610
rect 2390 8490 2430 8530
rect 7810 8730 7850 8770
rect 8350 8740 8390 8780
rect 9430 8740 9470 8780
rect 9840 8770 9880 8810
rect 10100 8770 10140 8810
rect 3080 8540 3120 8580
rect 3160 8540 3200 8580
rect 3490 8540 3530 8580
rect 3820 8540 3860 8580
rect 4110 8540 4150 8580
rect 4260 8530 4300 8570
rect 4980 8560 5020 8600
rect 5370 8480 5410 8520
rect 4930 8150 4970 8190
rect 5560 8150 5600 8190
rect 7370 8200 7410 8240
rect 10410 8200 10450 8240
rect -340 6920 -300 6960
rect 980 6920 1020 6960
rect 1560 6920 1600 6960
rect 2880 6920 2920 6960
rect -172 6588 -138 6622
rect -62 6588 -28 6622
rect 48 6588 82 6622
rect 158 6588 192 6622
rect 268 6588 302 6622
rect 378 6588 412 6622
rect 488 6588 522 6622
rect 598 6588 632 6622
rect 708 6588 742 6622
rect 818 6588 852 6622
rect 1728 6588 1762 6622
rect 1838 6588 1872 6622
rect 1948 6588 1982 6622
rect 2058 6588 2092 6622
rect 2168 6588 2202 6622
rect 2278 6588 2312 6622
rect 2388 6588 2422 6622
rect 2498 6588 2532 6622
rect 2608 6588 2642 6622
rect 2718 6588 2752 6622
rect -350 6320 -310 6360
rect 2890 6320 2930 6360
rect 7270 6306 7304 6340
rect 8544 6306 8578 6340
rect 3520 6120 3560 6160
rect 3960 6120 4000 6160
rect 8230 6110 8270 6150
rect 8630 6110 8670 6150
rect 3740 5780 3780 5820
rect 7430 5720 7470 5760
rect 9430 5720 9470 5760
rect -80 5580 -40 5620
rect 100 5580 140 5620
rect 280 5580 320 5620
rect 460 5580 500 5620
rect 640 5580 680 5620
rect 820 5580 860 5620
rect 1000 5580 1040 5620
rect 1180 5580 1220 5620
rect 1360 5580 1400 5620
rect 1540 5580 1580 5620
rect 1720 5580 1760 5620
rect 1900 5580 1940 5620
rect 2080 5580 2120 5620
rect 2260 5580 2300 5620
rect 2440 5580 2480 5620
rect 2620 5580 2660 5620
rect 7540 5420 7590 5470
rect 8190 5420 8240 5470
rect 8680 5420 8720 5460
rect 9340 5420 9380 5460
rect 9820 5420 9860 5460
rect 10480 5420 10520 5460
rect 7740 5180 7780 5220
rect 8790 5180 8830 5220
rect 9230 5180 9270 5220
rect 10770 5180 10810 5220
rect 9930 5060 9970 5100
rect 7650 4840 7690 4880
rect 8090 4840 8130 4880
rect 8880 4850 8920 4890
rect 9930 4840 9970 4880
rect -1450 4760 -1410 4800
rect 950 4760 990 4800
rect 1590 4760 1630 4800
rect 3990 4760 4030 4800
rect 10770 4840 10810 4880
rect -1270 4410 -1230 4450
rect -1090 4420 -1050 4460
rect -610 4420 -570 4460
rect -370 4420 -330 4460
rect 110 4420 150 4460
rect 350 4420 390 4460
rect 770 4420 810 4460
rect 7540 4500 7580 4540
rect 8200 4500 8240 4540
rect 8680 4500 8720 4540
rect 9340 4500 9380 4540
rect 9820 4500 9860 4540
rect 10480 4500 10520 4540
rect 1770 4420 1810 4460
rect 2190 4420 2230 4460
rect 2430 4420 2470 4460
rect 2910 4420 2950 4460
rect 3150 4420 3190 4460
rect 3630 4420 3670 4460
rect 3810 4410 3850 4450
rect 7550 4190 7590 4230
rect 9550 4190 9590 4230
rect -446 3818 -412 3852
rect -288 3818 -254 3852
rect 36 3818 70 3852
rect 190 3818 224 3852
rect 514 3818 548 3852
rect -547 3588 -513 3622
rect -187 3588 -153 3622
rect -67 3588 -33 3622
rect 293 3588 327 3622
rect 413 3588 447 3622
rect 2032 3818 2066 3852
rect 2356 3818 2390 3852
rect 2510 3818 2544 3852
rect 2834 3818 2868 3852
rect 2992 3818 3026 3852
rect 2133 3588 2167 3622
rect 2253 3588 2287 3622
rect 2613 3588 2647 3622
rect 2733 3588 2767 3622
rect 3093 3588 3127 3622
rect 8350 3550 8390 3590
rect 8750 3550 8790 3590
rect -1050 3210 -1010 3250
rect -810 3210 -770 3250
rect -570 3210 -530 3250
rect -330 3210 -290 3250
rect 310 3210 350 3250
rect 550 3210 590 3250
rect 790 3210 830 3250
rect 1750 3210 1790 3250
rect 1990 3210 2030 3250
rect 2230 3210 2270 3250
rect 2870 3210 2910 3250
rect 3110 3210 3150 3250
rect 3350 3210 3390 3250
rect 3590 3210 3630 3250
rect -650 2300 -610 2340
rect -490 2300 -450 2340
rect -330 2300 -290 2340
rect -170 2300 -130 2340
rect -10 2300 30 2340
rect 150 2300 190 2340
rect 310 2300 350 2340
rect 470 2300 510 2340
rect 630 2300 670 2340
rect 790 2300 830 2340
rect 950 2300 990 2340
rect 1110 2300 1150 2340
rect 1430 2300 1470 2340
rect 1590 2300 1630 2340
rect 1750 2300 1790 2340
rect 1910 2300 1950 2340
rect 2070 2300 2110 2340
rect 2230 2300 2270 2340
rect 2390 2300 2430 2340
rect 2550 2300 2590 2340
rect 2710 2300 2750 2340
rect 2870 2300 2910 2340
rect 3030 2300 3070 2340
rect 3190 2300 3230 2340
<< xpolycontact >>
rect 11234 6274 11304 6706
rect 11234 5702 11304 6134
rect 11234 3810 11304 4242
rect 11234 3182 11304 3614
rect 642 1720 1082 1790
rect 1510 1720 1950 1790
rect -3536 -1318 -3466 -886
rect -3536 -2128 -3466 -1696
rect -2417 -919 -2347 -487
rect -2749 -2131 -2679 -1699
rect -1636 -388 -1566 44
rect -1304 -2128 -1234 -1696
rect 4016 -388 4086 44
rect 3684 -2128 3754 -1696
rect 4797 -1525 4867 -1093
rect 4797 -2125 4867 -1693
rect 5584 -1318 5654 -886
rect 5584 -2128 5654 -1696
rect 3002 -3176 3434 -3106
rect 4906 -3176 5338 -3106
<< npolyres >>
rect 7684 6290 8164 6356
<< ppolyres >>
rect -3536 -1696 -3466 -1318
rect 5584 -1696 5654 -1318
<< xpolyres >>
rect 11234 6134 11304 6274
rect 11234 3614 11304 3810
rect 1082 1720 1510 1790
rect -2749 -1093 -2513 -1023
rect -2749 -1699 -2679 -1093
rect -2583 -1525 -2513 -1093
rect -2417 -1525 -2347 -919
rect -2583 -1595 -2347 -1525
rect -1636 -1522 -1566 -388
rect -1470 -562 -1234 -492
rect -1470 -1522 -1400 -562
rect -1636 -1592 -1400 -1522
rect -1304 -1696 -1234 -562
rect 3684 -562 3920 -492
rect 3684 -1696 3754 -562
rect 3850 -1522 3920 -562
rect 4016 -1522 4086 -388
rect 3850 -1592 4086 -1522
rect 4797 -1693 4867 -1525
rect 3434 -3176 4906 -3106
<< locali >>
rect 11320 14450 11400 14470
rect 11840 14450 11920 14470
rect 12360 14450 12440 14470
rect 12850 14450 12930 14470
rect 11100 14410 11340 14450
rect 11380 14410 11860 14450
rect 11900 14410 12240 14450
rect 12420 14410 12870 14450
rect 12910 14410 13140 14450
rect 11100 13880 11140 14410
rect 11320 14390 11400 14410
rect 11840 14390 11920 14410
rect 12360 14390 12440 14410
rect 12850 14390 12930 14410
rect 11220 14320 11280 14340
rect 11220 14280 11230 14320
rect 11270 14280 11280 14320
rect 11220 14220 11280 14280
rect 11220 14180 11230 14220
rect 11270 14180 11280 14220
rect 11220 14160 11280 14180
rect 11330 14320 11390 14340
rect 11330 14280 11340 14320
rect 11380 14280 11390 14320
rect 11330 14220 11390 14280
rect 11330 14180 11340 14220
rect 11380 14180 11390 14220
rect 11330 14160 11390 14180
rect 11740 14320 11800 14340
rect 11740 14280 11750 14320
rect 11790 14280 11800 14320
rect 11740 14220 11800 14280
rect 11740 14180 11750 14220
rect 11790 14180 11800 14220
rect 11740 14160 11800 14180
rect 11850 14320 11910 14340
rect 11850 14280 11860 14320
rect 11900 14280 11910 14320
rect 11850 14220 11910 14280
rect 11850 14180 11860 14220
rect 11900 14180 11910 14220
rect 11850 14160 11910 14180
rect 12260 14320 12320 14340
rect 12260 14280 12270 14320
rect 12310 14280 12320 14320
rect 12260 14220 12320 14280
rect 12260 14180 12270 14220
rect 12310 14180 12320 14220
rect 12260 14160 12320 14180
rect 12370 14320 12430 14340
rect 12370 14280 12380 14320
rect 12420 14280 12430 14320
rect 12370 14220 12430 14280
rect 12370 14180 12380 14220
rect 12420 14180 12430 14220
rect 12370 14160 12430 14180
rect 12860 14320 12920 14340
rect 12860 14280 12870 14320
rect 12910 14280 12920 14320
rect 12860 14220 12920 14280
rect 12860 14180 12870 14220
rect 12910 14180 12920 14220
rect 12860 14160 12920 14180
rect 12970 14320 13030 14340
rect 12970 14280 12980 14320
rect 13020 14280 13030 14320
rect 12970 14220 13030 14280
rect 12970 14180 12980 14220
rect 13020 14180 13030 14220
rect 12970 14160 13030 14180
rect 11276 14102 11334 14120
rect 11276 14068 11288 14102
rect 11322 14068 11334 14102
rect 11276 14050 11334 14068
rect 11796 14102 11854 14120
rect 11796 14068 11808 14102
rect 11842 14068 11854 14102
rect 11796 14050 11854 14068
rect 12316 14102 12374 14120
rect 12316 14068 12328 14102
rect 12362 14068 12374 14102
rect 12316 14050 12374 14068
rect 12884 14102 12942 14120
rect 12884 14068 12896 14102
rect 12930 14068 12942 14102
rect 12884 14050 12942 14068
rect 11220 13940 11280 13960
rect 11220 13900 11230 13940
rect 11270 13900 11280 13940
rect 11220 13840 11280 13900
rect 11220 13800 11230 13840
rect 11270 13800 11280 13840
rect 11220 13740 11280 13800
rect 11220 13700 11230 13740
rect 11270 13700 11280 13740
rect 11220 13680 11280 13700
rect 11330 13940 11390 13960
rect 11330 13900 11340 13940
rect 11380 13900 11390 13940
rect 11330 13840 11390 13900
rect 11330 13800 11340 13840
rect 11380 13800 11390 13840
rect 11330 13740 11390 13800
rect 11330 13700 11340 13740
rect 11380 13700 11390 13740
rect 11330 13680 11390 13700
rect 11740 13940 11800 13960
rect 11740 13900 11750 13940
rect 11790 13900 11800 13940
rect 11740 13840 11800 13900
rect 11740 13800 11750 13840
rect 11790 13800 11800 13840
rect 11740 13740 11800 13800
rect 11740 13700 11750 13740
rect 11790 13700 11800 13740
rect 11740 13680 11800 13700
rect 11850 13940 11910 13960
rect 11850 13900 11860 13940
rect 11900 13900 11910 13940
rect 11850 13840 11910 13900
rect 11850 13800 11860 13840
rect 11900 13800 11910 13840
rect 11850 13740 11910 13800
rect 11850 13700 11860 13740
rect 11900 13700 11910 13740
rect 11850 13680 11910 13700
rect 12260 13940 12320 13960
rect 12260 13900 12270 13940
rect 12310 13900 12320 13940
rect 12260 13840 12320 13900
rect 12260 13800 12270 13840
rect 12310 13800 12320 13840
rect 12260 13740 12320 13800
rect 12260 13700 12270 13740
rect 12310 13700 12320 13740
rect 12260 13680 12320 13700
rect 12370 13940 12430 13960
rect 12370 13900 12380 13940
rect 12420 13900 12430 13940
rect 12370 13840 12430 13900
rect 12370 13800 12380 13840
rect 12420 13800 12430 13840
rect 12370 13740 12430 13800
rect 12370 13700 12380 13740
rect 12420 13700 12430 13740
rect 12370 13680 12430 13700
rect 13100 13880 13140 14410
rect 550 13420 630 13440
rect 550 13380 570 13420
rect 610 13380 630 13420
rect 550 13360 630 13380
rect 770 13420 850 13440
rect 770 13380 790 13420
rect 830 13380 850 13420
rect 770 13360 850 13380
rect 1240 13420 1320 13440
rect 1240 13380 1260 13420
rect 1300 13380 1320 13420
rect 1240 13360 1320 13380
rect 1580 13420 1660 13440
rect 1580 13380 1600 13420
rect 1640 13380 1660 13420
rect 1580 13360 1660 13380
rect 1800 13420 1880 13440
rect 1800 13380 1820 13420
rect 1860 13380 1880 13420
rect 1800 13360 1880 13380
rect 2240 13420 2320 13440
rect 2240 13380 2260 13420
rect 2300 13380 2320 13420
rect 2240 13360 2320 13380
rect 2920 13420 3000 13440
rect 2920 13380 2940 13420
rect 2980 13380 3000 13420
rect 2920 13360 3000 13380
rect 3140 13420 3220 13440
rect 3140 13380 3160 13420
rect 3200 13380 3220 13420
rect 3140 13360 3220 13380
rect 3610 13420 3690 13440
rect 3610 13380 3630 13420
rect 3670 13380 3690 13420
rect 3610 13360 3690 13380
rect 4070 13420 4150 13440
rect 4070 13380 4090 13420
rect 4130 13380 4150 13420
rect 4070 13360 4150 13380
rect 4420 13420 4500 13440
rect 4420 13380 4440 13420
rect 4480 13380 4500 13420
rect 4420 13360 4500 13380
rect 4670 13420 4750 13440
rect 4670 13380 4690 13420
rect 4730 13380 4750 13420
rect 4670 13360 4750 13380
rect 4890 13420 4970 13440
rect 4890 13380 4910 13420
rect 4950 13380 4970 13420
rect 4890 13360 4970 13380
rect 5220 13420 5300 13440
rect 5220 13380 5240 13420
rect 5280 13380 5300 13420
rect 5220 13360 5300 13380
rect 5880 13420 5960 13440
rect 5880 13380 5900 13420
rect 5940 13380 5960 13420
rect 5880 13360 5960 13380
rect 6100 13420 6180 13440
rect 6100 13380 6120 13420
rect 6160 13380 6180 13420
rect 6100 13360 6180 13380
rect 6670 13420 6750 13440
rect 6670 13380 6690 13420
rect 6730 13380 6750 13420
rect 6670 13360 6750 13380
rect 6930 13420 7010 13440
rect 6930 13380 6950 13420
rect 6990 13380 7010 13420
rect 6930 13360 7010 13380
rect 7180 13420 7260 13440
rect 7180 13380 7200 13420
rect 7240 13380 7260 13420
rect 7180 13360 7260 13380
rect 7400 13420 7480 13440
rect 7400 13380 7420 13420
rect 7460 13380 7480 13420
rect 7400 13360 7480 13380
rect 7950 13420 8030 13440
rect 7950 13380 7970 13420
rect 8010 13380 8030 13420
rect 7950 13360 8030 13380
rect 8230 13420 8310 13440
rect 8230 13380 8250 13420
rect 8290 13380 8310 13420
rect 8230 13360 8310 13380
rect 8480 13420 8560 13440
rect 8480 13380 8500 13420
rect 8540 13380 8560 13420
rect 8480 13360 8560 13380
rect 8700 13420 8780 13440
rect 8700 13380 8720 13420
rect 8760 13380 8780 13420
rect 8700 13360 8780 13380
rect 9250 13420 9330 13440
rect 9250 13380 9270 13420
rect 9310 13380 9330 13420
rect 9250 13360 9330 13380
rect 9530 13420 9610 13440
rect 9530 13380 9550 13420
rect 9590 13380 9610 13420
rect 9530 13360 9610 13380
rect 9780 13420 9860 13440
rect 9780 13380 9800 13420
rect 9840 13380 9860 13420
rect 9780 13360 9860 13380
rect 10000 13420 10080 13440
rect 10000 13380 10020 13420
rect 10060 13380 10080 13420
rect 10000 13360 10080 13380
rect 10550 13420 10630 13440
rect 10550 13380 10570 13420
rect 10610 13380 10630 13420
rect 10550 13360 10630 13380
rect 390 13310 470 13330
rect 390 13270 410 13310
rect 450 13270 470 13310
rect 390 13250 470 13270
rect 410 13210 450 13250
rect 570 13210 610 13360
rect 790 13210 830 13360
rect 1260 13210 1300 13360
rect 1340 13290 1420 13310
rect 1340 13250 1360 13290
rect 1400 13250 1420 13290
rect 1470 13300 1550 13320
rect 1470 13260 1490 13300
rect 1530 13260 1550 13300
rect 1470 13250 1550 13260
rect 1340 13230 1420 13250
rect 1490 13210 1530 13250
rect 1600 13210 1640 13360
rect 1820 13210 1860 13360
rect 2260 13210 2300 13360
rect 2410 13300 2490 13320
rect 2410 13260 2430 13300
rect 2470 13260 2490 13300
rect 2410 13250 2490 13260
rect 2940 13210 2980 13360
rect 3160 13210 3200 13360
rect 3630 13210 3670 13360
rect 3970 13300 4050 13320
rect 3970 13260 3990 13300
rect 4030 13260 4050 13300
rect 3970 13250 4050 13260
rect 4090 13210 4130 13360
rect 4440 13210 4480 13360
rect 4690 13210 4730 13360
rect 4910 13210 4950 13360
rect 5240 13210 5280 13360
rect 5900 13210 5940 13360
rect 6120 13210 6160 13360
rect 6584 13310 6650 13330
rect 6584 13270 6594 13310
rect 6634 13270 6650 13310
rect 6584 13250 6650 13270
rect 6690 13210 6730 13360
rect 6950 13300 6990 13360
rect 7200 13300 7240 13360
rect 7420 13300 7460 13360
rect 7970 13300 8010 13360
rect 8250 13300 8290 13360
rect 8500 13300 8540 13360
rect 8720 13300 8760 13360
rect 9270 13300 9310 13360
rect 9550 13300 9590 13360
rect 9800 13300 9840 13360
rect 10020 13300 10060 13360
rect 10570 13300 10610 13360
rect 6940 13280 7000 13300
rect 7080 13280 7140 13300
rect 6940 13240 6950 13280
rect 6990 13240 7000 13280
rect 6940 13220 7000 13240
rect 7040 13240 7090 13280
rect 7130 13240 7140 13280
rect 7040 13220 7140 13240
rect 7190 13280 7250 13300
rect 7190 13240 7200 13280
rect 7240 13240 7250 13280
rect 7190 13220 7250 13240
rect 7300 13280 7360 13300
rect 7300 13240 7310 13280
rect 7350 13240 7360 13280
rect 7300 13220 7360 13240
rect 7410 13280 7470 13300
rect 7410 13240 7420 13280
rect 7460 13240 7470 13280
rect 7410 13220 7470 13240
rect 7520 13280 7580 13300
rect 7520 13240 7530 13280
rect 7570 13240 7580 13280
rect 7740 13280 7800 13300
rect 7740 13260 7750 13280
rect 7520 13220 7580 13240
rect 7620 13240 7750 13260
rect 7790 13240 7800 13280
rect 7620 13220 7800 13240
rect 7850 13280 7910 13300
rect 7850 13240 7860 13280
rect 7900 13240 7910 13280
rect 7850 13220 7910 13240
rect 7960 13280 8020 13300
rect 7960 13240 7970 13280
rect 8010 13240 8020 13280
rect 7960 13220 8020 13240
rect 8070 13280 8130 13300
rect 8070 13240 8080 13280
rect 8120 13240 8130 13280
rect 8070 13220 8130 13240
rect 8240 13280 8300 13300
rect 8380 13280 8440 13300
rect 8240 13240 8250 13280
rect 8290 13240 8300 13280
rect 8240 13220 8300 13240
rect 8340 13240 8390 13280
rect 8430 13240 8440 13280
rect 8340 13220 8440 13240
rect 8490 13280 8550 13300
rect 8490 13240 8500 13280
rect 8540 13240 8550 13280
rect 8490 13220 8550 13240
rect 8600 13280 8660 13300
rect 8600 13240 8610 13280
rect 8650 13240 8660 13280
rect 8600 13220 8660 13240
rect 8710 13280 8770 13300
rect 8710 13240 8720 13280
rect 8760 13240 8770 13280
rect 8710 13220 8770 13240
rect 8820 13280 8880 13300
rect 8820 13240 8830 13280
rect 8870 13240 8880 13280
rect 9040 13280 9100 13300
rect 9040 13260 9050 13280
rect 8820 13220 8880 13240
rect 8920 13240 9050 13260
rect 9090 13240 9100 13280
rect 8920 13220 9100 13240
rect 9150 13280 9210 13300
rect 9150 13240 9160 13280
rect 9200 13240 9210 13280
rect 9150 13220 9210 13240
rect 9260 13280 9320 13300
rect 9260 13240 9270 13280
rect 9310 13240 9320 13280
rect 9260 13220 9320 13240
rect 9370 13280 9430 13300
rect 9370 13240 9380 13280
rect 9420 13240 9430 13280
rect 9370 13220 9430 13240
rect 9540 13280 9600 13300
rect 9680 13280 9740 13300
rect 9540 13240 9550 13280
rect 9590 13240 9600 13280
rect 9540 13220 9600 13240
rect 9640 13240 9690 13280
rect 9730 13240 9740 13280
rect 9640 13220 9740 13240
rect 9790 13280 9850 13300
rect 9790 13240 9800 13280
rect 9840 13240 9850 13280
rect 9790 13220 9850 13240
rect 9900 13280 9960 13300
rect 9900 13240 9910 13280
rect 9950 13240 9960 13280
rect 9900 13220 9960 13240
rect 10010 13280 10070 13300
rect 10010 13240 10020 13280
rect 10060 13240 10070 13280
rect 10010 13220 10070 13240
rect 10120 13280 10180 13300
rect 10120 13240 10130 13280
rect 10170 13240 10180 13280
rect 10340 13280 10400 13300
rect 10340 13260 10350 13280
rect 10120 13220 10180 13240
rect 10220 13240 10350 13260
rect 10390 13240 10400 13280
rect 10220 13220 10400 13240
rect 10450 13280 10510 13300
rect 10450 13240 10460 13280
rect 10500 13240 10510 13280
rect 10450 13220 10510 13240
rect 10560 13280 10620 13300
rect 10560 13240 10570 13280
rect 10610 13240 10620 13280
rect 10560 13220 10620 13240
rect 10670 13280 10730 13300
rect 10670 13240 10680 13280
rect 10720 13240 10730 13280
rect 10670 13220 10730 13240
rect 410 13190 510 13210
rect 410 13150 460 13190
rect 500 13150 510 13190
rect 410 13130 510 13150
rect 560 13190 620 13210
rect 560 13150 570 13190
rect 610 13150 620 13190
rect 560 13130 620 13150
rect 670 13190 730 13210
rect 670 13150 680 13190
rect 720 13150 730 13190
rect 670 13130 730 13150
rect 780 13190 840 13210
rect 780 13150 790 13190
rect 830 13150 840 13190
rect 780 13130 840 13150
rect 890 13190 950 13210
rect 1030 13190 1090 13210
rect 890 13150 900 13190
rect 940 13150 950 13190
rect 890 13130 950 13150
rect 990 13150 1040 13190
rect 1080 13150 1090 13190
rect 990 13130 1090 13150
rect 1140 13190 1200 13210
rect 1140 13150 1150 13190
rect 1190 13150 1200 13190
rect 1140 13130 1200 13150
rect 1250 13190 1310 13210
rect 1250 13150 1260 13190
rect 1300 13150 1310 13190
rect 1250 13130 1310 13150
rect 1480 13190 1540 13210
rect 1480 13150 1490 13190
rect 1530 13150 1540 13190
rect 1480 13130 1540 13150
rect 1590 13190 1650 13210
rect 1590 13150 1600 13190
rect 1640 13150 1650 13190
rect 1590 13130 1650 13150
rect 1700 13190 1760 13210
rect 1700 13150 1710 13190
rect 1750 13150 1760 13190
rect 1700 13130 1760 13150
rect 1810 13190 1870 13210
rect 1810 13150 1820 13190
rect 1860 13150 1870 13190
rect 1810 13130 1870 13150
rect 1920 13190 1980 13210
rect 1920 13150 1930 13190
rect 1970 13150 1980 13190
rect 1920 13130 1980 13150
rect 2140 13190 2200 13210
rect 2140 13150 2150 13190
rect 2190 13150 2200 13190
rect 2140 13130 2200 13150
rect 2250 13190 2310 13210
rect 2250 13150 2260 13190
rect 2300 13150 2310 13190
rect 2250 13130 2310 13150
rect 2360 13190 2420 13210
rect 2360 13150 2370 13190
rect 2410 13150 2420 13190
rect 2360 13130 2420 13150
rect 2470 13190 2530 13210
rect 2470 13150 2480 13190
rect 2520 13150 2530 13190
rect 2470 13130 2530 13150
rect 2580 13190 2640 13210
rect 2820 13190 2880 13210
rect 2580 13150 2590 13190
rect 2630 13150 2680 13190
rect 2580 13130 2680 13150
rect 410 13060 450 13130
rect 680 13090 720 13130
rect 900 13090 940 13130
rect 330 13040 450 13060
rect 330 13000 350 13040
rect 390 13000 450 13040
rect 500 13070 940 13090
rect 500 13030 520 13070
rect 560 13050 940 13070
rect 560 13030 580 13050
rect 500 13010 580 13030
rect 330 12980 450 13000
rect 410 12890 450 12980
rect 370 12870 450 12890
rect 610 12870 670 12890
rect 370 12830 390 12870
rect 430 12830 620 12870
rect 660 12830 670 12870
rect 370 12810 450 12830
rect 610 12810 670 12830
rect 720 12870 860 12890
rect 720 12830 730 12870
rect 770 12830 810 12870
rect 850 12830 860 12870
rect 900 12870 940 13050
rect 990 12970 1030 13130
rect 1480 13090 1520 13130
rect 1700 13090 1740 13130
rect 1920 13090 1960 13130
rect 2150 13090 2190 13130
rect 2370 13090 2410 13130
rect 1080 13070 1160 13090
rect 1420 13070 1520 13090
rect 1080 13030 1100 13070
rect 1140 13030 1440 13070
rect 1480 13030 1520 13070
rect 1080 13010 1160 13030
rect 1420 13010 1520 13030
rect 1660 13050 1960 13090
rect 1660 13010 1700 13050
rect 990 12930 1300 12970
rect 1260 12890 1300 12930
rect 1030 12870 1090 12890
rect 900 12830 1040 12870
rect 1080 12830 1090 12870
rect 720 12810 860 12830
rect 1030 12810 1090 12830
rect 1140 12870 1200 12890
rect 1140 12830 1150 12870
rect 1190 12830 1200 12870
rect 1140 12810 1200 12830
rect 1250 12870 1310 12890
rect 1250 12830 1260 12870
rect 1300 12830 1310 12870
rect 1480 12870 1520 13010
rect 1620 12990 1700 13010
rect 1620 12950 1640 12990
rect 1680 12950 1700 12990
rect 1620 12930 1700 12950
rect 1920 12890 1960 13050
rect 2000 13070 2080 13090
rect 2000 13030 2020 13070
rect 2060 13030 2080 13070
rect 2150 13050 2410 13090
rect 2520 13070 2600 13090
rect 2000 13020 2080 13030
rect 2520 13030 2540 13070
rect 2580 13030 2600 13070
rect 2520 13020 2600 13030
rect 2640 12970 2680 13130
rect 2020 12950 2680 12970
rect 2020 12910 2040 12950
rect 2080 12930 2680 12950
rect 2780 13150 2830 13190
rect 2870 13150 2880 13190
rect 2780 13130 2880 13150
rect 2930 13190 2990 13210
rect 2930 13150 2940 13190
rect 2980 13150 2990 13190
rect 2930 13130 2990 13150
rect 3040 13190 3100 13210
rect 3040 13150 3050 13190
rect 3090 13150 3100 13190
rect 3040 13130 3100 13150
rect 3150 13190 3210 13210
rect 3150 13150 3160 13190
rect 3200 13150 3210 13190
rect 3150 13130 3210 13150
rect 3260 13190 3320 13210
rect 3400 13190 3460 13210
rect 3260 13150 3270 13190
rect 3310 13150 3320 13190
rect 3260 13130 3320 13150
rect 3360 13150 3410 13190
rect 3450 13150 3460 13190
rect 3360 13130 3460 13150
rect 3510 13190 3570 13210
rect 3510 13150 3520 13190
rect 3560 13150 3570 13190
rect 3510 13130 3570 13150
rect 3620 13190 3760 13210
rect 3960 13190 4020 13210
rect 3620 13150 3630 13190
rect 3670 13150 3710 13190
rect 3750 13150 3760 13190
rect 3620 13130 3760 13150
rect 3800 13150 3970 13190
rect 4010 13150 4020 13190
rect 2080 12910 2100 12930
rect 2020 12890 2100 12910
rect 2150 12890 2190 12930
rect 2480 12890 2520 12930
rect 2780 12890 2820 13130
rect 3050 13090 3090 13130
rect 3270 13090 3310 13130
rect 2870 13070 3310 13090
rect 2870 13030 2890 13070
rect 2930 13050 3310 13070
rect 2930 13030 2950 13050
rect 2870 13020 2950 13030
rect 1700 12870 1760 12890
rect 1480 12830 1710 12870
rect 1750 12830 1760 12870
rect 1250 12810 1310 12830
rect 1700 12810 1760 12830
rect 1810 12870 1870 12890
rect 1810 12830 1820 12870
rect 1860 12830 1870 12870
rect 1810 12810 1870 12830
rect 1920 12870 1980 12890
rect 1920 12830 1930 12870
rect 1970 12830 1980 12870
rect 1920 12810 1980 12830
rect 2140 12870 2200 12890
rect 2140 12830 2150 12870
rect 2190 12830 2200 12870
rect 2140 12810 2200 12830
rect 2250 12870 2310 12890
rect 2250 12830 2260 12870
rect 2300 12830 2310 12870
rect 2250 12810 2310 12830
rect 2360 12870 2430 12890
rect 2360 12830 2370 12870
rect 2410 12830 2430 12870
rect 2360 12810 2430 12830
rect 2470 12870 2530 12890
rect 2470 12830 2480 12870
rect 2520 12830 2530 12870
rect 2470 12810 2530 12830
rect 2740 12870 2820 12890
rect 2980 12870 3040 12890
rect 2740 12830 2760 12870
rect 2800 12830 2990 12870
rect 3030 12830 3040 12870
rect 2740 12810 2820 12830
rect 2980 12810 3040 12830
rect 3090 12870 3230 12890
rect 3090 12830 3100 12870
rect 3140 12830 3180 12870
rect 3220 12830 3230 12870
rect 3270 12870 3310 13050
rect 3360 12970 3400 13130
rect 3450 13070 3530 13090
rect 3660 13070 3740 13090
rect 3450 13030 3470 13070
rect 3510 13030 3680 13070
rect 3720 13030 3740 13070
rect 3450 13010 3530 13030
rect 3660 13020 3740 13030
rect 3800 12970 3840 13150
rect 3960 13130 4020 13150
rect 4070 13190 4130 13210
rect 4070 13150 4080 13190
rect 4120 13150 4130 13190
rect 4070 13130 4130 13150
rect 4320 13190 4380 13210
rect 4320 13150 4330 13190
rect 4370 13150 4380 13190
rect 4320 13130 4380 13150
rect 4430 13190 4490 13210
rect 4430 13150 4440 13190
rect 4480 13150 4490 13190
rect 4430 13130 4490 13150
rect 4570 13190 4630 13210
rect 4570 13150 4580 13190
rect 4620 13150 4630 13190
rect 4570 13130 4630 13150
rect 4680 13190 4740 13210
rect 4680 13150 4690 13190
rect 4730 13150 4740 13190
rect 4680 13130 4740 13150
rect 4790 13190 4850 13210
rect 4790 13150 4800 13190
rect 4840 13150 4850 13190
rect 4790 13130 4850 13150
rect 4900 13190 4960 13210
rect 4900 13150 4910 13190
rect 4950 13150 4960 13190
rect 4900 13130 4960 13150
rect 5010 13190 5070 13210
rect 5010 13150 5020 13190
rect 5060 13150 5070 13190
rect 5010 13130 5070 13150
rect 5150 13190 5290 13210
rect 5150 13150 5160 13190
rect 5200 13150 5240 13190
rect 5280 13150 5290 13190
rect 5150 13130 5290 13150
rect 5340 13190 5400 13210
rect 5340 13150 5350 13190
rect 5390 13150 5400 13190
rect 5340 13130 5400 13150
rect 5450 13190 5510 13210
rect 5450 13150 5460 13190
rect 5500 13150 5510 13190
rect 5450 13130 5510 13150
rect 5560 13190 5620 13210
rect 5780 13190 5840 13210
rect 5560 13150 5570 13190
rect 5610 13150 5660 13190
rect 5560 13130 5660 13150
rect 3900 13070 3980 13090
rect 4330 13080 4370 13130
rect 3900 13030 3920 13070
rect 3960 13050 3980 13070
rect 4240 13060 4370 13080
rect 4240 13050 4260 13060
rect 3960 13030 4260 13050
rect 3900 13020 4260 13030
rect 4300 13020 4370 13060
rect 4570 13040 4610 13130
rect 4790 13090 4830 13130
rect 5010 13090 5050 13130
rect 3900 13010 4370 13020
rect 4240 13000 4370 13010
rect 3360 12930 3670 12970
rect 3630 12890 3670 12930
rect 3720 12950 4120 12970
rect 3720 12910 3740 12950
rect 3780 12930 4120 12950
rect 3780 12910 3800 12930
rect 3720 12890 3800 12910
rect 3860 12890 3900 12930
rect 4080 12890 4120 12930
rect 4330 12890 4370 13000
rect 4510 13020 4610 13040
rect 4510 12980 4530 13020
rect 4570 12980 4610 13020
rect 4750 13050 5050 13090
rect 4750 13010 4790 13050
rect 4510 12960 4610 12980
rect 3400 12870 3460 12890
rect 3270 12830 3410 12870
rect 3450 12830 3460 12870
rect 3090 12810 3230 12830
rect 3400 12810 3460 12830
rect 3510 12870 3570 12890
rect 3510 12830 3520 12870
rect 3560 12830 3570 12870
rect 3510 12810 3570 12830
rect 3620 12870 3680 12890
rect 3620 12830 3630 12870
rect 3670 12830 3680 12870
rect 3620 12810 3680 12830
rect 3850 12870 3910 12890
rect 3850 12830 3860 12870
rect 3900 12830 3910 12870
rect 3850 12810 3910 12830
rect 3960 12870 4020 12890
rect 3960 12830 3970 12870
rect 4010 12830 4020 12870
rect 3960 12810 4020 12830
rect 4070 12870 4130 12890
rect 4070 12830 4080 12870
rect 4120 12830 4130 12870
rect 4070 12810 4130 12830
rect 4210 12870 4270 12890
rect 4210 12830 4220 12870
rect 4260 12830 4270 12870
rect 4210 12810 4270 12830
rect 4320 12870 4380 12890
rect 4320 12830 4330 12870
rect 4370 12830 4380 12870
rect 4320 12810 4380 12830
rect 4430 12870 4490 12890
rect 4430 12830 4440 12870
rect 4480 12830 4490 12870
rect 4570 12870 4610 12960
rect 4710 12990 4790 13010
rect 4710 12950 4730 12990
rect 4770 12950 4790 12990
rect 4710 12930 4790 12950
rect 5010 12890 5050 13050
rect 5140 13070 5220 13090
rect 5500 13070 5580 13090
rect 5140 13030 5160 13070
rect 5200 13030 5520 13070
rect 5560 13030 5580 13070
rect 5140 13020 5220 13030
rect 5500 13020 5580 13030
rect 5110 12950 5500 12970
rect 5110 12910 5130 12950
rect 5170 12930 5500 12950
rect 5170 12910 5190 12930
rect 5110 12890 5190 12910
rect 5240 12890 5280 12930
rect 5460 12890 5500 12930
rect 4790 12870 4850 12890
rect 4570 12830 4800 12870
rect 4840 12830 4850 12870
rect 4430 12810 4490 12830
rect 4790 12810 4850 12830
rect 4900 12870 4960 12890
rect 4900 12830 4910 12870
rect 4950 12830 4960 12870
rect 4900 12810 4960 12830
rect 5010 12870 5070 12890
rect 5010 12830 5020 12870
rect 5060 12830 5070 12870
rect 5010 12810 5070 12830
rect 5230 12870 5290 12890
rect 5230 12830 5240 12870
rect 5280 12830 5290 12870
rect 5230 12810 5290 12830
rect 5340 12870 5400 12890
rect 5340 12830 5350 12870
rect 5390 12830 5400 12870
rect 5340 12810 5400 12830
rect 5450 12870 5510 12890
rect 5620 12870 5660 13130
rect 5740 13150 5790 13190
rect 5830 13150 5840 13190
rect 5740 13130 5840 13150
rect 5890 13190 5950 13210
rect 5890 13150 5900 13190
rect 5940 13150 5950 13190
rect 5890 13130 5950 13150
rect 6000 13190 6060 13210
rect 6000 13150 6010 13190
rect 6050 13150 6060 13190
rect 6000 13130 6060 13150
rect 6110 13190 6170 13210
rect 6110 13150 6120 13190
rect 6160 13150 6170 13190
rect 6110 13130 6170 13150
rect 6220 13190 6280 13210
rect 6220 13150 6230 13190
rect 6270 13150 6280 13190
rect 6440 13190 6500 13210
rect 6440 13170 6450 13190
rect 6220 13130 6280 13150
rect 6320 13150 6450 13170
rect 6490 13150 6500 13190
rect 6320 13130 6500 13150
rect 6550 13190 6610 13210
rect 6550 13150 6560 13190
rect 6600 13150 6610 13190
rect 6550 13130 6610 13150
rect 6660 13190 6730 13210
rect 6660 13150 6670 13190
rect 6710 13150 6730 13190
rect 6660 13130 6730 13150
rect 6770 13190 6830 13210
rect 6770 13150 6780 13190
rect 6820 13150 6830 13190
rect 6770 13130 6830 13150
rect 5740 12890 5780 13130
rect 6010 13090 6050 13130
rect 6230 13090 6270 13130
rect 5830 13070 6270 13090
rect 5830 13030 5850 13070
rect 5890 13050 6270 13070
rect 5890 13030 5910 13050
rect 5830 13020 5910 13030
rect 6160 12890 6200 13050
rect 6320 13010 6360 13130
rect 6780 13090 6820 13130
rect 6410 13070 6820 13090
rect 6410 13030 6430 13070
rect 6470 13050 6820 13070
rect 6470 13030 6490 13050
rect 6410 13010 6490 13030
rect 6240 12990 6360 13010
rect 6240 12950 6260 12990
rect 6300 12970 6360 12990
rect 6300 12950 6460 12970
rect 6240 12930 6460 12950
rect 6420 12890 6460 12930
rect 6560 12890 6600 13050
rect 6780 12890 6820 13050
rect 6880 13050 6960 13070
rect 6880 13010 6900 13050
rect 6940 13030 6960 13050
rect 7040 13030 7080 13220
rect 7310 13180 7350 13220
rect 7530 13180 7570 13220
rect 7130 13160 7570 13180
rect 7130 13120 7150 13160
rect 7190 13140 7570 13160
rect 7190 13120 7210 13140
rect 7130 13100 7210 13120
rect 6940 13010 7080 13030
rect 6880 12990 7080 13010
rect 5450 12830 5460 12870
rect 5500 12830 5660 12870
rect 5700 12870 5780 12890
rect 5850 12870 5910 12890
rect 5700 12830 5720 12870
rect 5760 12830 5860 12870
rect 5900 12830 5910 12870
rect 5450 12810 5510 12830
rect 5700 12810 5780 12830
rect 5850 12810 5910 12830
rect 5960 12870 6100 12890
rect 5960 12830 5970 12870
rect 6010 12830 6050 12870
rect 6090 12830 6100 12870
rect 5960 12810 6100 12830
rect 6160 12870 6250 12890
rect 6160 12830 6200 12870
rect 6240 12830 6250 12870
rect 6160 12810 6250 12830
rect 6300 12870 6360 12890
rect 6300 12830 6310 12870
rect 6350 12830 6360 12870
rect 6300 12810 6360 12830
rect 6410 12870 6470 12890
rect 6410 12830 6420 12870
rect 6460 12830 6470 12870
rect 6410 12810 6470 12830
rect 6550 12870 6610 12890
rect 6550 12830 6560 12870
rect 6600 12830 6610 12870
rect 6550 12810 6610 12830
rect 6660 12870 6720 12890
rect 6660 12830 6670 12870
rect 6710 12830 6720 12870
rect 6660 12810 6720 12830
rect 6770 12870 6830 12890
rect 6770 12830 6780 12870
rect 6820 12830 6830 12870
rect 7040 12870 7080 12990
rect 7460 12890 7500 13140
rect 7620 13010 7660 13220
rect 8080 13180 8120 13220
rect 7710 13160 8120 13180
rect 7710 13120 7730 13160
rect 7770 13140 8120 13160
rect 7770 13120 7790 13140
rect 7710 13100 7790 13120
rect 7540 12990 7660 13010
rect 7540 12950 7560 12990
rect 7600 12970 7660 12990
rect 7600 12950 7760 12970
rect 7540 12930 7760 12950
rect 7720 12890 7760 12930
rect 7860 12890 7900 13140
rect 8080 12890 8120 13140
rect 8180 13050 8260 13070
rect 8180 13010 8200 13050
rect 8240 13030 8260 13050
rect 8340 13030 8380 13220
rect 8610 13180 8650 13220
rect 8830 13180 8870 13220
rect 8430 13160 8870 13180
rect 8430 13120 8450 13160
rect 8490 13140 8870 13160
rect 8490 13120 8510 13140
rect 8430 13100 8510 13120
rect 8240 13010 8380 13030
rect 8180 12990 8380 13010
rect 7150 12870 7210 12890
rect 7040 12830 7160 12870
rect 7200 12830 7210 12870
rect 6770 12810 6830 12830
rect 7150 12810 7210 12830
rect 7260 12870 7400 12890
rect 7260 12830 7270 12870
rect 7310 12830 7350 12870
rect 7390 12830 7400 12870
rect 7260 12810 7400 12830
rect 7460 12870 7550 12890
rect 7460 12830 7500 12870
rect 7540 12830 7550 12870
rect 7460 12810 7550 12830
rect 7600 12870 7660 12890
rect 7600 12830 7610 12870
rect 7650 12830 7660 12870
rect 7600 12810 7660 12830
rect 7710 12870 7770 12890
rect 7710 12830 7720 12870
rect 7760 12830 7770 12870
rect 7710 12810 7770 12830
rect 7850 12870 7910 12890
rect 7850 12830 7860 12870
rect 7900 12830 7910 12870
rect 7850 12810 7910 12830
rect 7960 12870 8020 12890
rect 7960 12830 7970 12870
rect 8010 12830 8020 12870
rect 7960 12810 8020 12830
rect 8070 12870 8130 12890
rect 8070 12830 8080 12870
rect 8120 12830 8130 12870
rect 8340 12870 8380 12990
rect 8760 12890 8800 13140
rect 8920 13010 8960 13220
rect 9380 13180 9420 13220
rect 9010 13160 9420 13180
rect 9010 13120 9030 13160
rect 9070 13140 9420 13160
rect 9070 13120 9090 13140
rect 9010 13100 9090 13120
rect 8840 12990 8960 13010
rect 8840 12950 8860 12990
rect 8900 12970 8960 12990
rect 8900 12950 9060 12970
rect 8840 12930 9060 12950
rect 9020 12890 9060 12930
rect 9160 12890 9200 13140
rect 9380 12890 9420 13140
rect 9480 13050 9560 13070
rect 9480 13010 9500 13050
rect 9540 13030 9560 13050
rect 9640 13030 9680 13220
rect 9910 13180 9950 13220
rect 10130 13180 10170 13220
rect 9730 13160 10170 13180
rect 9730 13120 9750 13160
rect 9790 13140 10170 13160
rect 9790 13120 9810 13140
rect 9730 13100 9810 13120
rect 9540 13010 9680 13030
rect 9480 12990 9680 13010
rect 8450 12870 8510 12890
rect 8340 12830 8460 12870
rect 8500 12830 8510 12870
rect 8070 12810 8130 12830
rect 8450 12810 8510 12830
rect 8560 12870 8700 12890
rect 8560 12830 8570 12870
rect 8610 12830 8650 12870
rect 8690 12830 8700 12870
rect 8560 12810 8700 12830
rect 8760 12870 8850 12890
rect 8760 12830 8800 12870
rect 8840 12830 8850 12870
rect 8760 12810 8850 12830
rect 8900 12870 8960 12890
rect 8900 12830 8910 12870
rect 8950 12830 8960 12870
rect 8900 12810 8960 12830
rect 9010 12870 9070 12890
rect 9010 12830 9020 12870
rect 9060 12830 9070 12870
rect 9010 12810 9070 12830
rect 9150 12870 9210 12890
rect 9150 12830 9160 12870
rect 9200 12830 9210 12870
rect 9150 12810 9210 12830
rect 9260 12870 9320 12890
rect 9260 12830 9270 12870
rect 9310 12830 9320 12870
rect 9260 12810 9320 12830
rect 9370 12870 9430 12890
rect 9370 12830 9380 12870
rect 9420 12830 9430 12870
rect 9640 12870 9680 12990
rect 10060 12890 10100 13140
rect 10220 13010 10260 13220
rect 10680 13180 10720 13220
rect 10310 13160 10720 13180
rect 10310 13120 10330 13160
rect 10370 13140 10720 13160
rect 10370 13120 10390 13140
rect 10310 13100 10390 13120
rect 10140 12990 10260 13010
rect 10140 12950 10160 12990
rect 10200 12970 10260 12990
rect 10200 12950 10360 12970
rect 10140 12930 10360 12950
rect 10320 12890 10360 12930
rect 10460 12890 10500 13140
rect 10680 12890 10720 13140
rect 11100 13150 11140 13670
rect 11290 13622 11348 13640
rect 11290 13588 11302 13622
rect 11336 13588 11348 13622
rect 11290 13570 11348 13588
rect 11810 13622 11868 13640
rect 11810 13588 11822 13622
rect 11856 13588 11868 13622
rect 11810 13570 11868 13588
rect 12330 13622 12388 13640
rect 12330 13588 12342 13622
rect 12376 13588 12388 13622
rect 12330 13570 12388 13588
rect 11218 13460 11278 13480
rect 11218 13420 11228 13460
rect 11268 13420 11278 13460
rect 11218 13360 11278 13420
rect 11218 13320 11228 13360
rect 11268 13320 11278 13360
rect 11218 13300 11278 13320
rect 11330 13460 11390 13480
rect 11330 13420 11340 13460
rect 11380 13420 11390 13460
rect 11330 13360 11390 13420
rect 11330 13320 11340 13360
rect 11380 13320 11390 13360
rect 11330 13300 11390 13320
rect 11738 13460 11798 13480
rect 11738 13420 11748 13460
rect 11788 13420 11798 13460
rect 11738 13360 11798 13420
rect 11738 13320 11748 13360
rect 11788 13320 11798 13360
rect 11738 13300 11798 13320
rect 11850 13460 11910 13480
rect 11850 13420 11860 13460
rect 11900 13420 11910 13460
rect 11850 13360 11910 13420
rect 11850 13320 11860 13360
rect 11900 13320 11910 13360
rect 11850 13300 11910 13320
rect 12258 13460 12318 13480
rect 12258 13420 12268 13460
rect 12308 13420 12318 13460
rect 12258 13360 12318 13420
rect 12258 13320 12268 13360
rect 12308 13320 12318 13360
rect 12258 13300 12318 13320
rect 12370 13460 12430 13480
rect 12370 13420 12380 13460
rect 12420 13420 12430 13460
rect 12370 13360 12430 13420
rect 12370 13320 12380 13360
rect 12420 13320 12430 13360
rect 12370 13300 12430 13320
rect 11262 13242 11320 13260
rect 11262 13208 11274 13242
rect 11308 13208 11320 13242
rect 11262 13190 11320 13208
rect 11782 13242 11840 13260
rect 11782 13208 11794 13242
rect 11828 13208 11840 13242
rect 11782 13190 11840 13208
rect 12302 13242 12360 13260
rect 12302 13208 12314 13242
rect 12348 13208 12360 13242
rect 12302 13190 12360 13208
rect 13100 13150 13140 13670
rect 11100 13110 12240 13150
rect 12380 13110 13140 13150
rect 10762 13042 10820 13070
rect 10762 13008 10774 13042
rect 10808 13008 10820 13042
rect 10762 12990 10820 13008
rect 11100 12910 12120 12950
rect 12280 12910 13330 12950
rect 9750 12870 9810 12890
rect 9640 12830 9760 12870
rect 9800 12830 9810 12870
rect 9370 12810 9430 12830
rect 9750 12810 9810 12830
rect 9860 12870 10000 12890
rect 9860 12830 9870 12870
rect 9910 12830 9950 12870
rect 9990 12830 10000 12870
rect 9860 12810 10000 12830
rect 10060 12870 10150 12890
rect 10060 12830 10100 12870
rect 10140 12830 10150 12870
rect 10060 12810 10150 12830
rect 10200 12870 10260 12890
rect 10200 12830 10210 12870
rect 10250 12830 10260 12870
rect 10200 12810 10260 12830
rect 10310 12870 10370 12890
rect 10310 12830 10320 12870
rect 10360 12830 10370 12870
rect 10310 12810 10370 12830
rect 10450 12870 10510 12890
rect 10450 12830 10460 12870
rect 10500 12830 10510 12870
rect 10450 12810 10510 12830
rect 10560 12870 10620 12890
rect 10560 12830 10570 12870
rect 10610 12830 10620 12870
rect 10560 12810 10620 12830
rect 10670 12870 10730 12890
rect 10670 12830 10680 12870
rect 10720 12830 10730 12870
rect 10670 12810 10730 12830
rect 730 12660 770 12810
rect 1030 12750 1110 12770
rect 1030 12710 1050 12750
rect 1090 12710 1110 12750
rect 1030 12690 1110 12710
rect 1150 12660 1190 12810
rect 1260 12770 1300 12810
rect 1230 12750 1300 12770
rect 1230 12710 1240 12750
rect 1280 12710 1300 12750
rect 1340 12770 1420 12790
rect 1340 12730 1360 12770
rect 1400 12730 1420 12770
rect 1340 12710 1420 12730
rect 1230 12690 1300 12710
rect 1820 12660 1860 12810
rect 2150 12750 2230 12770
rect 2150 12710 2170 12750
rect 2210 12710 2230 12750
rect 2150 12690 2230 12710
rect 2290 12750 2350 12770
rect 2290 12710 2300 12750
rect 2340 12710 2350 12750
rect 2290 12690 2350 12710
rect 2390 12660 2430 12810
rect 3100 12660 3140 12810
rect 3410 12750 3490 12770
rect 3410 12710 3430 12750
rect 3470 12710 3490 12750
rect 3410 12690 3490 12710
rect 3530 12660 3570 12810
rect 3630 12770 3670 12810
rect 3630 12750 3710 12770
rect 3630 12710 3650 12750
rect 3690 12710 3710 12750
rect 3630 12690 3710 12710
rect 3970 12660 4010 12810
rect 4220 12660 4260 12810
rect 4440 12660 4480 12810
rect 4800 12760 4840 12810
rect 4760 12740 4840 12760
rect 4760 12700 4780 12740
rect 4820 12700 4840 12740
rect 4760 12690 4840 12700
rect 4910 12660 4950 12810
rect 5170 12740 5250 12760
rect 5170 12700 5190 12740
rect 5230 12700 5250 12740
rect 5170 12690 5250 12700
rect 5350 12660 5390 12810
rect 5970 12660 6010 12810
rect 6310 12660 6350 12810
rect 6670 12660 6710 12810
rect 7160 12770 7200 12810
rect 7120 12750 7200 12770
rect 7120 12710 7140 12750
rect 7180 12710 7200 12750
rect 7120 12690 7200 12710
rect 7270 12660 7310 12810
rect 7610 12660 7650 12810
rect 7700 12750 7780 12770
rect 7700 12710 7720 12750
rect 7760 12710 7780 12750
rect 7700 12690 7780 12710
rect 7970 12660 8010 12810
rect 8460 12770 8500 12810
rect 8420 12750 8500 12770
rect 8420 12710 8440 12750
rect 8480 12710 8500 12750
rect 8420 12690 8500 12710
rect 8570 12660 8610 12810
rect 8910 12660 8950 12810
rect 9000 12750 9080 12770
rect 9000 12710 9020 12750
rect 9060 12710 9080 12750
rect 9000 12690 9080 12710
rect 9270 12660 9310 12810
rect 9760 12770 9800 12810
rect 9720 12750 9800 12770
rect 9720 12710 9740 12750
rect 9780 12710 9800 12750
rect 9720 12690 9800 12710
rect 9870 12660 9910 12810
rect 10210 12660 10250 12810
rect 10300 12750 10380 12770
rect 10300 12710 10320 12750
rect 10360 12710 10380 12750
rect 10300 12690 10380 12710
rect 10570 12660 10610 12810
rect 710 12640 790 12660
rect 710 12600 730 12640
rect 770 12600 790 12640
rect 710 12580 790 12600
rect 1130 12640 1210 12660
rect 1130 12600 1150 12640
rect 1190 12600 1210 12640
rect 1130 12580 1210 12600
rect 1800 12640 1880 12660
rect 1800 12600 1820 12640
rect 1860 12600 1880 12640
rect 1800 12580 1880 12600
rect 2370 12640 2450 12660
rect 2370 12600 2390 12640
rect 2430 12600 2450 12640
rect 2370 12580 2450 12600
rect 3080 12640 3160 12660
rect 3080 12600 3100 12640
rect 3140 12600 3160 12640
rect 3080 12580 3160 12600
rect 3510 12640 3590 12660
rect 3510 12600 3530 12640
rect 3570 12600 3590 12640
rect 3510 12580 3590 12600
rect 3950 12640 4030 12660
rect 3950 12600 3970 12640
rect 4010 12600 4030 12640
rect 3950 12580 4030 12600
rect 4200 12640 4280 12660
rect 4200 12600 4220 12640
rect 4260 12600 4280 12640
rect 4200 12580 4280 12600
rect 4420 12640 4500 12660
rect 4420 12600 4440 12640
rect 4480 12600 4500 12640
rect 4420 12580 4500 12600
rect 4890 12640 4970 12660
rect 4890 12600 4910 12640
rect 4950 12600 4970 12640
rect 4890 12580 4970 12600
rect 5330 12640 5410 12660
rect 5330 12600 5350 12640
rect 5390 12600 5410 12640
rect 5330 12580 5410 12600
rect 5950 12640 6030 12660
rect 5950 12600 5970 12640
rect 6010 12600 6030 12640
rect 5950 12580 6030 12600
rect 6290 12640 6370 12660
rect 6290 12600 6310 12640
rect 6350 12600 6370 12640
rect 6290 12580 6370 12600
rect 6650 12640 6730 12660
rect 6650 12600 6670 12640
rect 6710 12600 6730 12640
rect 6650 12580 6730 12600
rect 7250 12640 7330 12660
rect 7250 12600 7270 12640
rect 7310 12600 7330 12640
rect 7250 12580 7330 12600
rect 7590 12640 7670 12660
rect 7590 12600 7610 12640
rect 7650 12600 7670 12640
rect 7590 12580 7670 12600
rect 7950 12640 8030 12660
rect 7950 12600 7970 12640
rect 8010 12600 8030 12640
rect 7950 12580 8030 12600
rect 8550 12640 8630 12660
rect 8550 12600 8570 12640
rect 8610 12600 8630 12640
rect 8550 12580 8630 12600
rect 8890 12640 8970 12660
rect 8890 12600 8910 12640
rect 8950 12600 8970 12640
rect 8890 12580 8970 12600
rect 9250 12640 9330 12660
rect 9250 12600 9270 12640
rect 9310 12600 9330 12640
rect 9250 12580 9330 12600
rect 9850 12640 9930 12660
rect 9850 12600 9870 12640
rect 9910 12600 9930 12640
rect 9850 12580 9930 12600
rect 10190 12640 10270 12660
rect 10190 12600 10210 12640
rect 10250 12600 10270 12640
rect 10190 12580 10270 12600
rect 10550 12640 10630 12660
rect 10550 12600 10570 12640
rect 10610 12600 10630 12640
rect 10550 12580 10630 12600
rect 11100 11600 11140 12910
rect 11262 12852 11320 12870
rect 11262 12818 11274 12852
rect 11308 12818 11320 12852
rect 11262 12800 11320 12818
rect 11782 12852 11840 12870
rect 11782 12818 11794 12852
rect 11828 12818 11840 12852
rect 11782 12800 11840 12818
rect 12302 12852 12360 12870
rect 12302 12818 12314 12852
rect 12348 12818 12360 12852
rect 12302 12800 12360 12818
rect 11218 12740 11278 12760
rect 11218 12700 11228 12740
rect 11268 12700 11278 12740
rect 11218 12640 11278 12700
rect 11218 12600 11228 12640
rect 11268 12600 11278 12640
rect 11218 12540 11278 12600
rect 11218 12500 11228 12540
rect 11268 12500 11278 12540
rect 11218 12440 11278 12500
rect 11218 12400 11228 12440
rect 11268 12400 11278 12440
rect 11218 12380 11278 12400
rect 11330 12740 11390 12760
rect 11330 12700 11340 12740
rect 11380 12700 11390 12740
rect 11330 12640 11390 12700
rect 11330 12600 11340 12640
rect 11380 12600 11390 12640
rect 11330 12540 11390 12600
rect 11330 12500 11340 12540
rect 11380 12500 11390 12540
rect 11330 12440 11390 12500
rect 11330 12400 11340 12440
rect 11380 12400 11390 12440
rect 11330 12380 11390 12400
rect 11738 12740 11798 12760
rect 11738 12700 11748 12740
rect 11788 12700 11798 12740
rect 11738 12640 11798 12700
rect 11738 12600 11748 12640
rect 11788 12600 11798 12640
rect 11738 12540 11798 12600
rect 11738 12500 11748 12540
rect 11788 12500 11798 12540
rect 11738 12440 11798 12500
rect 11738 12400 11748 12440
rect 11788 12400 11798 12440
rect 11738 12380 11798 12400
rect 11850 12740 11910 12760
rect 11850 12700 11860 12740
rect 11900 12700 11910 12740
rect 11850 12640 11910 12700
rect 11850 12600 11860 12640
rect 11900 12600 11910 12640
rect 11850 12540 11910 12600
rect 11850 12500 11860 12540
rect 11900 12500 11910 12540
rect 11850 12440 11910 12500
rect 11850 12400 11860 12440
rect 11900 12400 11910 12440
rect 11850 12380 11910 12400
rect 12258 12740 12318 12760
rect 12258 12700 12268 12740
rect 12308 12700 12318 12740
rect 12258 12640 12318 12700
rect 12258 12600 12268 12640
rect 12308 12600 12318 12640
rect 12258 12540 12318 12600
rect 12258 12500 12268 12540
rect 12308 12500 12318 12540
rect 12258 12440 12318 12500
rect 12258 12400 12268 12440
rect 12308 12400 12318 12440
rect 12258 12380 12318 12400
rect 12370 12740 12430 12760
rect 12370 12700 12380 12740
rect 12420 12700 12430 12740
rect 12370 12640 12430 12700
rect 12370 12600 12380 12640
rect 12420 12600 12430 12640
rect 12370 12540 12430 12600
rect 12370 12500 12380 12540
rect 12420 12500 12430 12540
rect 12370 12440 12430 12500
rect 12370 12400 12380 12440
rect 12420 12400 12430 12440
rect 12370 12380 12430 12400
rect 11290 12272 11348 12290
rect 11290 12238 11302 12272
rect 11336 12238 11348 12272
rect 11290 12220 11348 12238
rect 11810 12272 11868 12290
rect 11810 12238 11822 12272
rect 11856 12238 11868 12272
rect 11810 12220 11868 12238
rect 12330 12272 12388 12290
rect 12330 12238 12342 12272
rect 12376 12238 12388 12272
rect 12330 12220 12388 12238
rect 11220 12160 11280 12180
rect 11220 12120 11230 12160
rect 11270 12120 11280 12160
rect 11220 12060 11280 12120
rect 11220 12020 11230 12060
rect 11270 12020 11280 12060
rect 11220 11960 11280 12020
rect 11220 11920 11230 11960
rect 11270 11920 11280 11960
rect 11220 11860 11280 11920
rect 11220 11820 11230 11860
rect 11270 11820 11280 11860
rect 11220 11760 11280 11820
rect 11220 11720 11230 11760
rect 11270 11720 11280 11760
rect 11220 11660 11280 11720
rect 11220 11620 11230 11660
rect 11270 11620 11280 11660
rect 11220 11600 11280 11620
rect 11330 12160 11390 12180
rect 11330 12120 11340 12160
rect 11380 12120 11390 12160
rect 11330 12060 11390 12120
rect 11330 12020 11340 12060
rect 11380 12020 11390 12060
rect 11330 11960 11390 12020
rect 11330 11920 11340 11960
rect 11380 11920 11390 11960
rect 11330 11860 11390 11920
rect 11330 11820 11340 11860
rect 11380 11820 11390 11860
rect 11330 11760 11390 11820
rect 11330 11720 11340 11760
rect 11380 11720 11390 11760
rect 11330 11660 11390 11720
rect 11330 11620 11340 11660
rect 11380 11620 11390 11660
rect 11330 11600 11390 11620
rect 11740 12160 11800 12180
rect 11740 12120 11750 12160
rect 11790 12120 11800 12160
rect 11740 12060 11800 12120
rect 11740 12020 11750 12060
rect 11790 12020 11800 12060
rect 11740 11960 11800 12020
rect 11740 11920 11750 11960
rect 11790 11920 11800 11960
rect 11740 11860 11800 11920
rect 11740 11820 11750 11860
rect 11790 11820 11800 11860
rect 11740 11760 11800 11820
rect 11740 11720 11750 11760
rect 11790 11720 11800 11760
rect 11740 11660 11800 11720
rect 11740 11620 11750 11660
rect 11790 11620 11800 11660
rect 11740 11600 11800 11620
rect 11850 12160 11910 12180
rect 11850 12120 11860 12160
rect 11900 12120 11910 12160
rect 11850 12060 11910 12120
rect 11850 12020 11860 12060
rect 11900 12020 11910 12060
rect 11850 11960 11910 12020
rect 11850 11920 11860 11960
rect 11900 11920 11910 11960
rect 11850 11860 11910 11920
rect 11850 11820 11860 11860
rect 11900 11820 11910 11860
rect 11850 11760 11910 11820
rect 11850 11720 11860 11760
rect 11900 11720 11910 11760
rect 11850 11660 11910 11720
rect 11850 11620 11860 11660
rect 11900 11620 11910 11660
rect 11850 11600 11910 11620
rect 12260 12160 12320 12180
rect 12260 12120 12270 12160
rect 12310 12120 12320 12160
rect 12260 12060 12320 12120
rect 12260 12020 12270 12060
rect 12310 12020 12320 12060
rect 12260 11960 12320 12020
rect 12260 11920 12270 11960
rect 12310 11920 12320 11960
rect 12260 11860 12320 11920
rect 12260 11820 12270 11860
rect 12310 11820 12320 11860
rect 12260 11760 12320 11820
rect 12260 11720 12270 11760
rect 12310 11720 12320 11760
rect 12260 11660 12320 11720
rect 12260 11620 12270 11660
rect 12310 11620 12320 11660
rect 12260 11600 12320 11620
rect 12370 12160 12430 12180
rect 12370 12120 12380 12160
rect 12420 12120 12430 12160
rect 12370 12060 12430 12120
rect 12370 12020 12380 12060
rect 12420 12020 12430 12060
rect 12370 11960 12430 12020
rect 12370 11920 12380 11960
rect 12420 11920 12430 11960
rect 12370 11860 12430 11920
rect 12370 11820 12380 11860
rect 12420 11820 12430 11860
rect 12370 11760 12430 11820
rect 12370 11720 12380 11760
rect 12420 11720 12430 11760
rect 12370 11660 12430 11720
rect 12370 11620 12380 11660
rect 12420 11620 12430 11660
rect 12370 11600 12430 11620
rect 13290 11600 13330 12910
rect 11400 11390 11480 11410
rect 11400 11350 11420 11390
rect 11460 11350 11480 11390
rect 11400 11330 11480 11350
rect 11920 11390 12000 11410
rect 11920 11350 11940 11390
rect 11980 11350 12000 11390
rect 11920 11330 12000 11350
rect 12440 11390 12520 11410
rect 12440 11350 12460 11390
rect 12500 11350 12520 11390
rect 12440 11330 12520 11350
rect 12970 11390 13030 11410
rect 12970 11350 12980 11390
rect 13020 11350 13030 11390
rect 12970 11330 13030 11350
rect 11100 10840 11140 11270
rect 11220 11270 11280 11290
rect 11220 11230 11230 11270
rect 11270 11230 11280 11270
rect 11220 11170 11280 11230
rect 11220 11130 11230 11170
rect 11270 11130 11280 11170
rect 11220 11070 11280 11130
rect 11220 11030 11230 11070
rect 11270 11030 11280 11070
rect 11220 10970 11280 11030
rect 11220 10930 11230 10970
rect 11270 10930 11280 10970
rect 11220 10910 11280 10930
rect 11600 11270 11660 11290
rect 11600 11230 11610 11270
rect 11650 11230 11660 11270
rect 11600 11170 11660 11230
rect 11600 11130 11610 11170
rect 11650 11130 11660 11170
rect 11600 11070 11660 11130
rect 11600 11030 11610 11070
rect 11650 11030 11660 11070
rect 11600 10970 11660 11030
rect 11600 10930 11610 10970
rect 11650 10930 11660 10970
rect 11600 10910 11660 10930
rect 11740 11270 11800 11290
rect 11740 11230 11750 11270
rect 11790 11230 11800 11270
rect 11740 11170 11800 11230
rect 11740 11130 11750 11170
rect 11790 11130 11800 11170
rect 11740 11070 11800 11130
rect 11740 11030 11750 11070
rect 11790 11030 11800 11070
rect 11740 10970 11800 11030
rect 11740 10930 11750 10970
rect 11790 10930 11800 10970
rect 11740 10910 11800 10930
rect 12120 11270 12180 11290
rect 12120 11230 12130 11270
rect 12170 11230 12180 11270
rect 12120 11170 12180 11230
rect 12120 11130 12130 11170
rect 12170 11130 12180 11170
rect 12120 11070 12180 11130
rect 12120 11030 12130 11070
rect 12170 11030 12180 11070
rect 12120 10970 12180 11030
rect 12120 10930 12130 10970
rect 12170 10930 12180 10970
rect 12120 10910 12180 10930
rect 12260 11270 12320 11290
rect 12260 11230 12270 11270
rect 12310 11230 12320 11270
rect 12260 11170 12320 11230
rect 12260 11130 12270 11170
rect 12310 11130 12320 11170
rect 12260 11070 12320 11130
rect 12260 11030 12270 11070
rect 12310 11030 12320 11070
rect 12260 10970 12320 11030
rect 12260 10930 12270 10970
rect 12310 10930 12320 10970
rect 12260 10910 12320 10930
rect 12640 11270 12700 11290
rect 12640 11230 12650 11270
rect 12690 11230 12700 11270
rect 12640 11170 12700 11230
rect 12640 11130 12650 11170
rect 12690 11130 12700 11170
rect 12640 11070 12700 11130
rect 12640 11030 12650 11070
rect 12690 11030 12700 11070
rect 12640 10970 12700 11030
rect 12640 10930 12650 10970
rect 12690 10930 12700 10970
rect 12640 10910 12700 10930
rect 12780 11270 12840 11290
rect 12780 11230 12790 11270
rect 12830 11230 12840 11270
rect 12780 11170 12840 11230
rect 12780 11130 12790 11170
rect 12830 11130 12840 11170
rect 12780 11070 12840 11130
rect 12780 11030 12790 11070
rect 12830 11030 12840 11070
rect 12780 10970 12840 11030
rect 12780 10930 12790 10970
rect 12830 10930 12840 10970
rect 12780 10910 12840 10930
rect 13160 11270 13220 11290
rect 13160 11230 13170 11270
rect 13210 11230 13220 11270
rect 13160 11170 13220 11230
rect 13160 11130 13170 11170
rect 13210 11130 13220 11170
rect 13160 11070 13220 11130
rect 13160 11030 13170 11070
rect 13210 11030 13220 11070
rect 13160 10970 13220 11030
rect 13160 10930 13170 10970
rect 13210 10930 13220 10970
rect 13160 10910 13220 10930
rect 11590 10840 11670 10860
rect 12110 10840 12190 10860
rect 12630 10840 12710 10860
rect 13150 10840 13230 10860
rect 13290 10840 13330 11270
rect 11100 10800 11610 10840
rect 11650 10800 12120 10840
rect 12280 10800 12650 10840
rect 12690 10800 13160 10840
rect 13230 10800 13330 10840
rect 11590 10780 11670 10800
rect 12110 10780 12190 10800
rect 12630 10780 12710 10800
rect 13150 10780 13230 10800
rect 10990 10520 11100 10540
rect 1260 10440 1340 10460
rect 1260 10400 1280 10440
rect 1320 10400 1340 10440
rect 1260 10380 1340 10400
rect 1480 10440 1560 10460
rect 1480 10400 1500 10440
rect 1540 10400 1560 10440
rect 1480 10380 1560 10400
rect 1780 10440 1860 10460
rect 1780 10400 1800 10440
rect 1840 10400 1860 10440
rect 1780 10380 1860 10400
rect 2000 10440 2080 10460
rect 2000 10400 2020 10440
rect 2060 10400 2080 10440
rect 2000 10380 2080 10400
rect 2160 10440 2240 10460
rect 2160 10400 2180 10440
rect 2220 10400 2240 10440
rect 2160 10380 2240 10400
rect 2380 10440 2460 10460
rect 2380 10400 2400 10440
rect 2440 10400 2460 10440
rect 2380 10380 2460 10400
rect 2680 10440 2760 10460
rect 2680 10400 2700 10440
rect 2740 10400 2760 10440
rect 2680 10380 2760 10400
rect 2900 10440 2980 10460
rect 2900 10400 2920 10440
rect 2960 10400 2980 10440
rect 2900 10380 2980 10400
rect 3200 10440 3280 10460
rect 3200 10400 3220 10440
rect 3260 10400 3280 10440
rect 3200 10380 3280 10400
rect 3640 10440 3720 10460
rect 3640 10400 3660 10440
rect 3700 10400 3720 10440
rect 3640 10380 3720 10400
rect 3970 10440 4050 10460
rect 3970 10400 3990 10440
rect 4030 10400 4050 10440
rect 3970 10380 4050 10400
rect 4400 10440 4480 10460
rect 4400 10400 4420 10440
rect 4460 10400 4480 10440
rect 4400 10380 4480 10400
rect 4790 10440 4870 10460
rect 4790 10400 4810 10440
rect 4850 10400 4870 10440
rect 4790 10380 4870 10400
rect 5180 10440 5260 10460
rect 5180 10400 5200 10440
rect 5240 10400 5260 10440
rect 10990 10450 11010 10520
rect 11080 10450 11100 10520
rect 10990 10430 11100 10450
rect 5180 10380 5260 10400
rect 1280 10230 1320 10380
rect 1500 10230 1540 10380
rect 1670 10330 1750 10350
rect 1670 10290 1690 10330
rect 1730 10290 1750 10330
rect 1670 10270 1750 10290
rect 1190 10210 1330 10230
rect 1190 10170 1200 10210
rect 1240 10170 1280 10210
rect 1320 10170 1330 10210
rect 1190 10110 1330 10170
rect 1190 10070 1200 10110
rect 1240 10070 1280 10110
rect 1320 10070 1330 10110
rect 1190 10050 1330 10070
rect 1380 10210 1440 10230
rect 1380 10170 1390 10210
rect 1430 10170 1440 10210
rect 1380 10110 1440 10170
rect 1380 10070 1390 10110
rect 1430 10070 1440 10110
rect 1380 10050 1440 10070
rect 1490 10210 1550 10230
rect 1490 10170 1500 10210
rect 1540 10170 1550 10210
rect 1490 10110 1550 10170
rect 1490 10070 1500 10110
rect 1540 10070 1550 10110
rect 1490 10050 1550 10070
rect 1140 9950 1220 9970
rect 1140 9910 1160 9950
rect 1200 9910 1220 9950
rect 1140 9890 1220 9910
rect 1380 9890 1420 10050
rect 1470 9990 1550 10010
rect 1470 9950 1490 9990
rect 1530 9970 1550 9990
rect 1710 9970 1750 10270
rect 1800 10230 1840 10380
rect 2020 10230 2060 10380
rect 2180 10230 2220 10380
rect 2400 10230 2440 10380
rect 2700 10230 2740 10380
rect 2920 10230 2960 10380
rect 3220 10230 3260 10380
rect 3390 10330 3470 10350
rect 3390 10290 3410 10330
rect 3450 10290 3470 10330
rect 3390 10270 3470 10290
rect 3660 10230 3700 10380
rect 3990 10230 4030 10380
rect 4420 10230 4460 10380
rect 4810 10230 4850 10380
rect 5200 10230 5240 10380
rect 5470 10330 5550 10350
rect 5470 10290 5490 10330
rect 5530 10290 5550 10330
rect 5470 10270 5550 10290
rect 5490 10230 5530 10270
rect 1790 10210 1850 10230
rect 1790 10170 1800 10210
rect 1840 10170 1850 10210
rect 1790 10110 1850 10170
rect 1790 10070 1800 10110
rect 1840 10070 1850 10110
rect 1790 10050 1850 10070
rect 1900 10210 1960 10230
rect 1900 10170 1910 10210
rect 1950 10170 1960 10210
rect 1900 10110 1960 10170
rect 1900 10070 1910 10110
rect 1950 10070 1960 10110
rect 1900 10050 1960 10070
rect 2010 10210 2230 10230
rect 2010 10170 2020 10210
rect 2060 10170 2100 10210
rect 2140 10170 2180 10210
rect 2220 10170 2230 10210
rect 2010 10110 2230 10170
rect 2010 10070 2020 10110
rect 2060 10070 2100 10110
rect 2140 10070 2180 10110
rect 2220 10070 2230 10110
rect 2010 10050 2230 10070
rect 2280 10210 2340 10230
rect 2280 10170 2290 10210
rect 2330 10170 2340 10210
rect 2280 10110 2340 10170
rect 2280 10070 2290 10110
rect 2330 10070 2340 10110
rect 2280 10050 2340 10070
rect 2390 10210 2450 10230
rect 2390 10170 2400 10210
rect 2440 10170 2450 10210
rect 2390 10110 2450 10170
rect 2390 10070 2400 10110
rect 2440 10070 2450 10110
rect 2390 10050 2450 10070
rect 2690 10210 2750 10230
rect 2690 10170 2700 10210
rect 2740 10170 2750 10210
rect 2690 10110 2750 10170
rect 2690 10070 2700 10110
rect 2740 10070 2750 10110
rect 2690 10050 2750 10070
rect 2800 10210 2860 10230
rect 2800 10170 2810 10210
rect 2850 10170 2860 10210
rect 2800 10110 2860 10170
rect 2800 10070 2810 10110
rect 2850 10070 2860 10110
rect 2800 10050 2860 10070
rect 2910 10210 3050 10230
rect 2910 10170 2920 10210
rect 2960 10170 3000 10210
rect 3040 10170 3050 10210
rect 2910 10110 3050 10170
rect 2910 10070 2920 10110
rect 2960 10070 3000 10110
rect 3040 10070 3050 10110
rect 2910 10050 3050 10070
rect 3130 10210 3270 10230
rect 3130 10170 3140 10210
rect 3180 10170 3220 10210
rect 3260 10170 3270 10210
rect 3130 10110 3270 10170
rect 3130 10070 3140 10110
rect 3180 10070 3220 10110
rect 3260 10070 3270 10110
rect 3130 10050 3270 10070
rect 3320 10210 3380 10230
rect 3320 10170 3330 10210
rect 3370 10170 3380 10210
rect 3320 10110 3380 10170
rect 3320 10070 3330 10110
rect 3370 10070 3380 10110
rect 3320 10050 3380 10070
rect 3430 10210 3490 10230
rect 3430 10170 3440 10210
rect 3480 10170 3490 10210
rect 3430 10110 3490 10170
rect 3430 10070 3440 10110
rect 3480 10070 3490 10110
rect 3430 10050 3490 10070
rect 3570 10210 3710 10230
rect 3570 10170 3580 10210
rect 3620 10170 3660 10210
rect 3700 10170 3710 10210
rect 3570 10110 3710 10170
rect 3570 10070 3580 10110
rect 3620 10070 3660 10110
rect 3700 10070 3710 10110
rect 3570 10050 3710 10070
rect 3760 10210 3820 10230
rect 3760 10170 3770 10210
rect 3810 10170 3820 10210
rect 3760 10110 3820 10170
rect 3760 10070 3770 10110
rect 3810 10070 3820 10110
rect 3760 10050 3820 10070
rect 3900 10210 4040 10230
rect 3900 10170 3910 10210
rect 3950 10170 3990 10210
rect 4030 10170 4040 10210
rect 3900 10110 4040 10170
rect 3900 10070 3910 10110
rect 3950 10070 3990 10110
rect 4030 10070 4040 10110
rect 3900 10050 4040 10070
rect 4090 10210 4150 10230
rect 4090 10170 4100 10210
rect 4140 10170 4150 10210
rect 4090 10110 4150 10170
rect 4090 10070 4100 10110
rect 4140 10070 4150 10110
rect 4090 10050 4150 10070
rect 4320 10210 4480 10230
rect 4320 10170 4330 10210
rect 4370 10170 4420 10210
rect 4460 10170 4480 10210
rect 4320 10110 4480 10170
rect 4320 10070 4330 10110
rect 4370 10070 4420 10110
rect 4460 10070 4480 10110
rect 4320 10050 4480 10070
rect 4530 10210 4610 10230
rect 4530 10170 4550 10210
rect 4590 10170 4610 10210
rect 4530 10110 4610 10170
rect 4530 10070 4550 10110
rect 4590 10070 4610 10110
rect 4530 10050 4610 10070
rect 4710 10210 4870 10230
rect 4710 10170 4720 10210
rect 4760 10170 4810 10210
rect 4850 10170 4870 10210
rect 4710 10110 4870 10170
rect 4710 10070 4720 10110
rect 4760 10070 4810 10110
rect 4850 10070 4870 10110
rect 4710 10050 4870 10070
rect 4920 10210 5000 10230
rect 4920 10170 4940 10210
rect 4980 10170 5000 10210
rect 4920 10110 5000 10170
rect 4920 10070 4940 10110
rect 4980 10070 5000 10110
rect 4920 10050 5000 10070
rect 5100 10210 5260 10230
rect 5100 10170 5110 10210
rect 5150 10170 5200 10210
rect 5240 10170 5260 10210
rect 5100 10110 5260 10170
rect 5100 10070 5110 10110
rect 5150 10070 5200 10110
rect 5240 10070 5260 10110
rect 5100 10050 5260 10070
rect 5310 10210 5390 10230
rect 5310 10170 5330 10210
rect 5370 10170 5390 10210
rect 5310 10110 5390 10170
rect 5310 10070 5330 10110
rect 5370 10070 5390 10110
rect 5310 10050 5390 10070
rect 5470 10210 5550 10230
rect 5470 10170 5490 10210
rect 5530 10170 5550 10210
rect 5470 10110 5550 10170
rect 5470 10070 5490 10110
rect 5530 10070 5550 10110
rect 5470 10050 5550 10070
rect 5600 10210 5680 10230
rect 5600 10170 5620 10210
rect 5660 10170 5680 10210
rect 5600 10110 5680 10170
rect 5600 10070 5620 10110
rect 5660 10070 5680 10110
rect 5600 10050 5680 10070
rect 1530 9950 1750 9970
rect 1470 9930 1750 9950
rect 1380 9850 1540 9890
rect 1500 9810 1540 9850
rect 1190 9790 1330 9810
rect 1190 9750 1200 9790
rect 1240 9750 1280 9790
rect 1320 9750 1330 9790
rect 1190 9690 1330 9750
rect 1190 9650 1200 9690
rect 1240 9650 1280 9690
rect 1320 9650 1330 9690
rect 1190 9590 1330 9650
rect 1190 9550 1200 9590
rect 1240 9550 1280 9590
rect 1320 9550 1330 9590
rect 1190 9490 1330 9550
rect 1190 9450 1200 9490
rect 1240 9450 1280 9490
rect 1320 9450 1330 9490
rect 1190 9430 1330 9450
rect 1380 9790 1440 9810
rect 1380 9750 1390 9790
rect 1430 9750 1440 9790
rect 1380 9690 1440 9750
rect 1380 9650 1390 9690
rect 1430 9650 1440 9690
rect 1380 9590 1440 9650
rect 1380 9550 1390 9590
rect 1430 9550 1440 9590
rect 1380 9490 1440 9550
rect 1380 9450 1390 9490
rect 1430 9450 1440 9490
rect 1380 9430 1440 9450
rect 1490 9790 1550 9810
rect 1490 9750 1500 9790
rect 1540 9750 1550 9790
rect 1490 9690 1550 9750
rect 1490 9650 1500 9690
rect 1540 9650 1550 9690
rect 1490 9590 1550 9650
rect 1490 9550 1500 9590
rect 1540 9550 1550 9590
rect 1490 9490 1550 9550
rect 1490 9450 1500 9490
rect 1540 9480 1550 9490
rect 1590 9490 1670 9510
rect 1590 9480 1610 9490
rect 1540 9450 1610 9480
rect 1650 9450 1670 9490
rect 1490 9430 1670 9450
rect 1710 9470 1750 9930
rect 1910 9890 1950 10050
rect 1800 9850 1950 9890
rect 1990 9910 2070 9930
rect 1990 9870 2010 9910
rect 2050 9890 2070 9910
rect 2280 9890 2320 10050
rect 2370 9990 2450 10010
rect 2370 9950 2390 9990
rect 2430 9970 2450 9990
rect 2430 9950 2650 9970
rect 2370 9930 2650 9950
rect 2050 9870 2440 9890
rect 1990 9850 2440 9870
rect 1800 9810 1840 9850
rect 2400 9810 2440 9850
rect 1790 9790 1850 9810
rect 1790 9750 1800 9790
rect 1840 9750 1850 9790
rect 1790 9690 1850 9750
rect 1790 9650 1800 9690
rect 1840 9650 1850 9690
rect 1790 9590 1850 9650
rect 1790 9550 1800 9590
rect 1840 9550 1850 9590
rect 1790 9490 1850 9550
rect 1790 9470 1800 9490
rect 1710 9450 1800 9470
rect 1840 9450 1850 9490
rect 1710 9430 1850 9450
rect 1900 9790 1960 9810
rect 1900 9750 1910 9790
rect 1950 9750 1960 9790
rect 1900 9690 1960 9750
rect 1900 9650 1910 9690
rect 1950 9650 1960 9690
rect 1900 9590 1960 9650
rect 1900 9550 1910 9590
rect 1950 9550 1960 9590
rect 1900 9490 1960 9550
rect 1900 9450 1910 9490
rect 1950 9450 1960 9490
rect 1900 9430 1960 9450
rect 2010 9790 2230 9810
rect 2010 9750 2020 9790
rect 2060 9750 2100 9790
rect 2140 9750 2180 9790
rect 2220 9750 2230 9790
rect 2010 9690 2230 9750
rect 2010 9650 2020 9690
rect 2060 9650 2100 9690
rect 2140 9650 2180 9690
rect 2220 9650 2230 9690
rect 2010 9590 2230 9650
rect 2010 9550 2020 9590
rect 2060 9550 2100 9590
rect 2140 9550 2180 9590
rect 2220 9550 2230 9590
rect 2010 9490 2230 9550
rect 2010 9450 2020 9490
rect 2060 9450 2100 9490
rect 2140 9450 2180 9490
rect 2220 9450 2230 9490
rect 2010 9430 2230 9450
rect 2280 9790 2340 9810
rect 2280 9750 2290 9790
rect 2330 9750 2340 9790
rect 2280 9690 2340 9750
rect 2280 9650 2290 9690
rect 2330 9650 2340 9690
rect 2280 9590 2340 9650
rect 2280 9550 2290 9590
rect 2330 9550 2340 9590
rect 2280 9490 2340 9550
rect 2280 9450 2290 9490
rect 2330 9450 2340 9490
rect 2280 9430 2340 9450
rect 2390 9790 2450 9810
rect 2390 9750 2400 9790
rect 2440 9750 2450 9790
rect 2390 9690 2450 9750
rect 2390 9650 2400 9690
rect 2440 9650 2450 9690
rect 2390 9590 2450 9650
rect 2390 9550 2400 9590
rect 2440 9550 2450 9590
rect 2390 9490 2450 9550
rect 2390 9450 2400 9490
rect 2440 9480 2450 9490
rect 2490 9490 2570 9510
rect 2490 9480 2510 9490
rect 2440 9450 2510 9480
rect 2550 9450 2570 9490
rect 2390 9430 2570 9450
rect 2610 9470 2650 9930
rect 2810 9890 2850 10050
rect 3040 9980 3120 10000
rect 3040 9940 3060 9980
rect 3100 9940 3120 9980
rect 3040 9920 3120 9940
rect 3440 9960 3480 10050
rect 3780 9960 3820 10050
rect 4110 9960 4150 10050
rect 4260 9970 4340 9990
rect 3440 9940 3550 9960
rect 3440 9920 3490 9940
rect 2700 9850 2850 9890
rect 3330 9900 3490 9920
rect 3530 9900 3550 9940
rect 3330 9880 3550 9900
rect 3780 9940 3880 9960
rect 3780 9900 3820 9940
rect 3860 9900 3880 9940
rect 3780 9880 3880 9900
rect 4110 9940 4210 9960
rect 4110 9900 4150 9940
rect 4190 9900 4210 9940
rect 4260 9930 4280 9970
rect 4320 9930 4340 9970
rect 4260 9910 4340 9930
rect 4570 9940 4610 10050
rect 4960 9970 5000 10050
rect 5220 9990 5300 10010
rect 5220 9970 5240 9990
rect 4830 9940 4910 9960
rect 4110 9880 4210 9900
rect 4570 9900 4850 9940
rect 4890 9900 4910 9940
rect 2700 9810 2740 9850
rect 3330 9810 3370 9880
rect 3780 9810 3820 9880
rect 4110 9810 4150 9880
rect 4570 9810 4610 9900
rect 4830 9880 4910 9900
rect 4960 9950 5240 9970
rect 5280 9950 5300 9990
rect 4960 9930 5300 9950
rect 5350 9930 5390 10050
rect 4960 9810 5000 9930
rect 5350 9910 5430 9930
rect 5350 9870 5370 9910
rect 5410 9870 5430 9910
rect 5350 9850 5430 9870
rect 5350 9810 5390 9850
rect 5490 9810 5530 10050
rect 5620 10010 5660 10050
rect 5620 9990 6090 10010
rect 5620 9970 6030 9990
rect 5620 9810 5660 9970
rect 6010 9950 6030 9970
rect 6070 9950 6090 9990
rect 6010 9930 6090 9950
rect 5700 9910 5780 9930
rect 5700 9870 5720 9910
rect 5760 9870 5780 9910
rect 5700 9850 5780 9870
rect 6010 9810 6050 9930
rect 7550 9880 7630 9900
rect 7550 9840 7570 9880
rect 7610 9840 7630 9880
rect 7550 9820 7630 9840
rect 10390 9880 10470 9900
rect 10390 9840 10410 9880
rect 10450 9840 10470 9880
rect 10390 9820 10470 9840
rect 2690 9790 2750 9810
rect 2690 9750 2700 9790
rect 2740 9750 2750 9790
rect 2690 9690 2750 9750
rect 2690 9650 2700 9690
rect 2740 9650 2750 9690
rect 2690 9590 2750 9650
rect 2690 9550 2700 9590
rect 2740 9550 2750 9590
rect 2690 9490 2750 9550
rect 2690 9470 2700 9490
rect 2610 9450 2700 9470
rect 2740 9450 2750 9490
rect 2610 9430 2750 9450
rect 2800 9790 2860 9810
rect 2800 9750 2810 9790
rect 2850 9750 2860 9790
rect 2800 9690 2860 9750
rect 2800 9650 2810 9690
rect 2850 9650 2860 9690
rect 2800 9590 2860 9650
rect 2800 9550 2810 9590
rect 2850 9550 2860 9590
rect 2800 9490 2860 9550
rect 2800 9450 2810 9490
rect 2850 9450 2860 9490
rect 2800 9430 2860 9450
rect 2910 9790 3050 9810
rect 2910 9750 2920 9790
rect 2960 9750 3000 9790
rect 3040 9750 3050 9790
rect 2910 9690 3050 9750
rect 2910 9650 2920 9690
rect 2960 9650 3000 9690
rect 3040 9650 3050 9690
rect 2910 9590 3050 9650
rect 2910 9550 2920 9590
rect 2960 9550 3000 9590
rect 3040 9550 3050 9590
rect 2910 9490 3050 9550
rect 2910 9450 2920 9490
rect 2960 9450 3000 9490
rect 3040 9450 3050 9490
rect 2910 9430 3050 9450
rect 3130 9790 3270 9810
rect 3130 9750 3140 9790
rect 3180 9750 3220 9790
rect 3260 9750 3270 9790
rect 3130 9690 3270 9750
rect 3130 9650 3140 9690
rect 3180 9650 3220 9690
rect 3260 9650 3270 9690
rect 3130 9590 3270 9650
rect 3130 9550 3140 9590
rect 3180 9550 3220 9590
rect 3260 9550 3270 9590
rect 3130 9490 3270 9550
rect 3130 9450 3140 9490
rect 3180 9450 3220 9490
rect 3260 9450 3270 9490
rect 3130 9430 3270 9450
rect 3320 9790 3380 9810
rect 3320 9750 3330 9790
rect 3370 9750 3380 9790
rect 3320 9690 3380 9750
rect 3320 9650 3330 9690
rect 3370 9650 3380 9690
rect 3320 9590 3380 9650
rect 3320 9550 3330 9590
rect 3370 9550 3380 9590
rect 3320 9490 3380 9550
rect 3320 9450 3330 9490
rect 3370 9450 3380 9490
rect 3320 9430 3380 9450
rect 3430 9790 3490 9810
rect 3430 9750 3440 9790
rect 3480 9750 3490 9790
rect 3430 9690 3490 9750
rect 3430 9650 3440 9690
rect 3480 9650 3490 9690
rect 3430 9590 3490 9650
rect 3430 9550 3440 9590
rect 3480 9550 3490 9590
rect 3430 9490 3490 9550
rect 3430 9450 3440 9490
rect 3480 9450 3490 9490
rect 3430 9430 3490 9450
rect 3570 9790 3710 9810
rect 3570 9750 3580 9790
rect 3620 9750 3660 9790
rect 3700 9750 3710 9790
rect 3570 9690 3710 9750
rect 3570 9650 3580 9690
rect 3620 9650 3660 9690
rect 3700 9650 3710 9690
rect 3570 9590 3710 9650
rect 3570 9550 3580 9590
rect 3620 9550 3660 9590
rect 3700 9550 3710 9590
rect 3570 9490 3710 9550
rect 3570 9450 3580 9490
rect 3620 9450 3660 9490
rect 3700 9450 3710 9490
rect 3570 9430 3710 9450
rect 3760 9790 3820 9810
rect 3760 9750 3770 9790
rect 3810 9750 3820 9790
rect 3760 9690 3820 9750
rect 3760 9650 3770 9690
rect 3810 9650 3820 9690
rect 3760 9590 3820 9650
rect 3760 9550 3770 9590
rect 3810 9550 3820 9590
rect 3760 9490 3820 9550
rect 3760 9450 3770 9490
rect 3810 9450 3820 9490
rect 3760 9430 3820 9450
rect 3900 9790 4040 9810
rect 3900 9750 3910 9790
rect 3950 9750 3990 9790
rect 4030 9750 4040 9790
rect 3900 9690 4040 9750
rect 3900 9650 3910 9690
rect 3950 9650 3990 9690
rect 4030 9650 4040 9690
rect 3900 9590 4040 9650
rect 3900 9550 3910 9590
rect 3950 9550 3990 9590
rect 4030 9550 4040 9590
rect 3900 9490 4040 9550
rect 3900 9450 3910 9490
rect 3950 9450 3990 9490
rect 4030 9450 4040 9490
rect 3900 9430 4040 9450
rect 4090 9790 4150 9810
rect 4090 9750 4100 9790
rect 4140 9750 4150 9790
rect 4090 9690 4150 9750
rect 4090 9650 4100 9690
rect 4140 9650 4150 9690
rect 4090 9590 4150 9650
rect 4090 9550 4100 9590
rect 4140 9550 4150 9590
rect 4090 9490 4150 9550
rect 4090 9450 4100 9490
rect 4140 9450 4150 9490
rect 4090 9430 4150 9450
rect 4300 9790 4480 9810
rect 4300 9750 4320 9790
rect 4360 9750 4420 9790
rect 4460 9750 4480 9790
rect 4300 9690 4480 9750
rect 4300 9650 4320 9690
rect 4360 9650 4420 9690
rect 4460 9650 4480 9690
rect 4300 9590 4480 9650
rect 4300 9550 4320 9590
rect 4360 9550 4420 9590
rect 4460 9550 4480 9590
rect 4300 9490 4480 9550
rect 4300 9450 4320 9490
rect 4360 9450 4420 9490
rect 4460 9450 4480 9490
rect 4300 9430 4480 9450
rect 4530 9790 4610 9810
rect 4530 9750 4550 9790
rect 4590 9750 4610 9790
rect 4530 9690 4610 9750
rect 4530 9650 4550 9690
rect 4590 9650 4610 9690
rect 4530 9590 4610 9650
rect 4530 9550 4550 9590
rect 4590 9550 4610 9590
rect 4530 9490 4610 9550
rect 4530 9450 4550 9490
rect 4590 9450 4610 9490
rect 4530 9430 4610 9450
rect 4690 9790 4870 9810
rect 4690 9750 4710 9790
rect 4750 9750 4810 9790
rect 4850 9750 4870 9790
rect 4690 9690 4870 9750
rect 4690 9650 4710 9690
rect 4750 9650 4810 9690
rect 4850 9650 4870 9690
rect 4690 9590 4870 9650
rect 4690 9550 4710 9590
rect 4750 9550 4810 9590
rect 4850 9550 4870 9590
rect 4690 9490 4870 9550
rect 4690 9450 4710 9490
rect 4750 9450 4810 9490
rect 4850 9450 4870 9490
rect 4690 9430 4870 9450
rect 4920 9790 5000 9810
rect 4920 9750 4940 9790
rect 4980 9750 5000 9790
rect 4920 9690 5000 9750
rect 4920 9650 4940 9690
rect 4980 9650 5000 9690
rect 4920 9590 5000 9650
rect 4920 9550 4940 9590
rect 4980 9550 5000 9590
rect 4920 9490 5000 9550
rect 4920 9450 4940 9490
rect 4980 9450 5000 9490
rect 4920 9430 5000 9450
rect 5080 9790 5260 9810
rect 5080 9750 5100 9790
rect 5140 9750 5200 9790
rect 5240 9750 5260 9790
rect 5080 9690 5260 9750
rect 5080 9650 5100 9690
rect 5140 9650 5200 9690
rect 5240 9650 5260 9690
rect 5080 9590 5260 9650
rect 5080 9550 5100 9590
rect 5140 9550 5200 9590
rect 5240 9550 5260 9590
rect 5080 9490 5260 9550
rect 5080 9450 5100 9490
rect 5140 9450 5200 9490
rect 5240 9450 5260 9490
rect 5080 9430 5260 9450
rect 5310 9790 5390 9810
rect 5310 9750 5330 9790
rect 5370 9750 5390 9790
rect 5310 9690 5390 9750
rect 5310 9650 5330 9690
rect 5370 9650 5390 9690
rect 5310 9590 5390 9650
rect 5310 9550 5330 9590
rect 5370 9550 5390 9590
rect 5310 9490 5390 9550
rect 5310 9450 5330 9490
rect 5370 9450 5390 9490
rect 5310 9430 5390 9450
rect 5470 9790 5550 9810
rect 5470 9750 5490 9790
rect 5530 9750 5550 9790
rect 5470 9690 5550 9750
rect 5470 9650 5490 9690
rect 5530 9650 5550 9690
rect 5470 9590 5550 9650
rect 5470 9550 5490 9590
rect 5530 9550 5550 9590
rect 5470 9490 5550 9550
rect 5470 9450 5490 9490
rect 5530 9450 5550 9490
rect 5470 9430 5550 9450
rect 5600 9790 5680 9810
rect 5600 9750 5620 9790
rect 5660 9750 5680 9790
rect 5600 9690 5680 9750
rect 5600 9650 5620 9690
rect 5660 9650 5680 9690
rect 5600 9590 5680 9650
rect 5600 9550 5620 9590
rect 5660 9550 5680 9590
rect 5600 9490 5680 9550
rect 5600 9450 5620 9490
rect 5660 9450 5680 9490
rect 5600 9430 5680 9450
rect 5760 9790 5940 9810
rect 5760 9750 5780 9790
rect 5820 9750 5880 9790
rect 5920 9750 5940 9790
rect 5760 9690 5940 9750
rect 5760 9650 5780 9690
rect 5820 9650 5880 9690
rect 5920 9650 5940 9690
rect 5760 9590 5940 9650
rect 5760 9550 5780 9590
rect 5820 9550 5880 9590
rect 5920 9550 5940 9590
rect 5760 9490 5940 9550
rect 5760 9450 5780 9490
rect 5820 9450 5880 9490
rect 5920 9450 5940 9490
rect 5760 9430 5940 9450
rect 5990 9790 6070 9810
rect 5990 9750 6010 9790
rect 6050 9750 6070 9790
rect 5990 9690 6070 9750
rect 5990 9650 6010 9690
rect 6050 9650 6070 9690
rect 5990 9590 6070 9650
rect 5990 9550 6010 9590
rect 6050 9550 6070 9590
rect 5990 9490 6070 9550
rect 5990 9450 6010 9490
rect 6050 9450 6070 9490
rect 5990 9430 6070 9450
rect 7450 9760 7630 9780
rect 7450 9720 7470 9760
rect 7510 9720 7570 9760
rect 7610 9720 7630 9760
rect 7450 9660 7630 9720
rect 7450 9620 7470 9660
rect 7510 9620 7570 9660
rect 7610 9620 7630 9660
rect 7450 9560 7630 9620
rect 7450 9520 7470 9560
rect 7510 9520 7570 9560
rect 7610 9520 7630 9560
rect 7450 9460 7630 9520
rect 1280 9280 1320 9430
rect 2020 9280 2060 9430
rect 2180 9280 2220 9430
rect 2920 9280 2960 9430
rect 3180 9280 3220 9430
rect 3260 9370 3340 9390
rect 3260 9330 3280 9370
rect 3320 9330 3340 9370
rect 3260 9320 3340 9330
rect 3440 9280 3480 9430
rect 3660 9280 3700 9430
rect 3990 9280 4030 9430
rect 4420 9280 4460 9430
rect 4810 9280 4850 9430
rect 5200 9280 5240 9430
rect 5880 9280 5920 9430
rect 7450 9420 7470 9460
rect 7510 9420 7570 9460
rect 7610 9420 7630 9460
rect 7450 9400 7630 9420
rect 7770 9760 7850 9780
rect 7770 9720 7790 9760
rect 7830 9720 7850 9760
rect 7770 9660 7850 9720
rect 7770 9620 7790 9660
rect 7830 9620 7850 9660
rect 7770 9560 7850 9620
rect 7770 9520 7790 9560
rect 7830 9520 7850 9560
rect 7770 9460 7850 9520
rect 7770 9420 7790 9460
rect 7830 9420 7850 9460
rect 7770 9400 7850 9420
rect 7990 9760 8070 9780
rect 7990 9720 8010 9760
rect 8050 9720 8070 9760
rect 7990 9660 8070 9720
rect 7990 9620 8010 9660
rect 8050 9620 8070 9660
rect 7990 9560 8070 9620
rect 7990 9520 8010 9560
rect 8050 9520 8070 9560
rect 7990 9460 8070 9520
rect 7990 9420 8010 9460
rect 8050 9420 8070 9460
rect 7990 9400 8070 9420
rect 8210 9760 8290 9780
rect 8210 9720 8230 9760
rect 8270 9720 8290 9760
rect 8210 9660 8290 9720
rect 8210 9620 8230 9660
rect 8270 9620 8290 9660
rect 8210 9560 8290 9620
rect 8210 9520 8230 9560
rect 8270 9520 8290 9560
rect 8210 9460 8290 9520
rect 8210 9420 8230 9460
rect 8270 9420 8290 9460
rect 8210 9400 8290 9420
rect 8430 9760 8510 9780
rect 8430 9720 8450 9760
rect 8490 9720 8510 9760
rect 8430 9660 8510 9720
rect 8430 9620 8450 9660
rect 8490 9620 8510 9660
rect 8430 9560 8510 9620
rect 8430 9520 8450 9560
rect 8490 9520 8510 9560
rect 8430 9460 8510 9520
rect 8430 9420 8450 9460
rect 8490 9420 8510 9460
rect 8430 9400 8510 9420
rect 8650 9760 8730 9780
rect 8650 9720 8670 9760
rect 8710 9720 8730 9760
rect 8650 9660 8730 9720
rect 8650 9620 8670 9660
rect 8710 9620 8730 9660
rect 8650 9560 8730 9620
rect 8650 9520 8670 9560
rect 8710 9520 8730 9560
rect 8650 9460 8730 9520
rect 8650 9420 8670 9460
rect 8710 9420 8730 9460
rect 8650 9400 8730 9420
rect 8870 9760 9150 9780
rect 8870 9720 8890 9760
rect 8930 9720 8990 9760
rect 9030 9720 9090 9760
rect 9130 9720 9150 9760
rect 8870 9660 9150 9720
rect 8870 9620 8890 9660
rect 8930 9620 8990 9660
rect 9030 9620 9090 9660
rect 9130 9620 9150 9660
rect 8870 9560 9150 9620
rect 8870 9520 8890 9560
rect 8930 9520 8990 9560
rect 9030 9520 9090 9560
rect 9130 9520 9150 9560
rect 8870 9460 9150 9520
rect 8870 9420 8890 9460
rect 8930 9420 8990 9460
rect 9030 9420 9090 9460
rect 9130 9420 9150 9460
rect 8870 9400 9150 9420
rect 9290 9760 9370 9780
rect 9290 9720 9310 9760
rect 9350 9720 9370 9760
rect 9290 9660 9370 9720
rect 9290 9620 9310 9660
rect 9350 9620 9370 9660
rect 9290 9560 9370 9620
rect 9290 9520 9310 9560
rect 9350 9520 9370 9560
rect 9290 9460 9370 9520
rect 9290 9420 9310 9460
rect 9350 9420 9370 9460
rect 9290 9400 9370 9420
rect 9510 9760 9590 9780
rect 9510 9720 9530 9760
rect 9570 9720 9590 9760
rect 9510 9660 9590 9720
rect 9510 9620 9530 9660
rect 9570 9620 9590 9660
rect 9510 9560 9590 9620
rect 9510 9520 9530 9560
rect 9570 9520 9590 9560
rect 9510 9460 9590 9520
rect 9510 9420 9530 9460
rect 9570 9420 9590 9460
rect 9510 9400 9590 9420
rect 9730 9760 9810 9780
rect 9730 9720 9750 9760
rect 9790 9720 9810 9760
rect 9730 9660 9810 9720
rect 9730 9620 9750 9660
rect 9790 9620 9810 9660
rect 9730 9560 9810 9620
rect 9730 9520 9750 9560
rect 9790 9520 9810 9560
rect 9730 9460 9810 9520
rect 9730 9420 9750 9460
rect 9790 9420 9810 9460
rect 9730 9400 9810 9420
rect 9950 9760 10030 9780
rect 9950 9720 9970 9760
rect 10010 9720 10030 9760
rect 9950 9660 10030 9720
rect 9950 9620 9970 9660
rect 10010 9620 10030 9660
rect 9950 9560 10030 9620
rect 9950 9520 9970 9560
rect 10010 9520 10030 9560
rect 9950 9460 10030 9520
rect 9950 9420 9970 9460
rect 10010 9420 10030 9460
rect 9950 9400 10030 9420
rect 10170 9760 10250 9780
rect 10170 9720 10190 9760
rect 10230 9720 10250 9760
rect 10170 9660 10250 9720
rect 10170 9620 10190 9660
rect 10230 9620 10250 9660
rect 10170 9560 10250 9620
rect 10170 9520 10190 9560
rect 10230 9520 10250 9560
rect 10170 9460 10250 9520
rect 10170 9420 10190 9460
rect 10230 9420 10250 9460
rect 10170 9400 10250 9420
rect 10390 9760 10570 9780
rect 10390 9720 10410 9760
rect 10450 9720 10510 9760
rect 10550 9720 10570 9760
rect 10390 9660 10570 9720
rect 10390 9620 10410 9660
rect 10450 9620 10510 9660
rect 10550 9620 10570 9660
rect 10390 9560 10570 9620
rect 10390 9520 10410 9560
rect 10450 9520 10510 9560
rect 10550 9520 10570 9560
rect 10390 9460 10570 9520
rect 10390 9420 10410 9460
rect 10450 9420 10510 9460
rect 10550 9420 10570 9460
rect 10390 9400 10570 9420
rect 8210 9340 8290 9360
rect 8210 9300 8230 9340
rect 8270 9300 8290 9340
rect 8210 9280 8290 9300
rect 8970 9340 9050 9400
rect 8970 9300 8990 9340
rect 9030 9300 9050 9340
rect 10750 9340 10860 9360
rect 8970 9280 9050 9300
rect 9380 9310 9460 9330
rect 1260 9260 1340 9280
rect 1260 9220 1280 9260
rect 1320 9220 1340 9260
rect 1260 9200 1340 9220
rect 2000 9260 2080 9280
rect 2000 9220 2020 9260
rect 2060 9220 2080 9260
rect 2000 9200 2080 9220
rect 2160 9260 2240 9280
rect 2160 9220 2180 9260
rect 2220 9220 2240 9260
rect 2160 9200 2240 9220
rect 2900 9260 2980 9280
rect 2900 9220 2920 9260
rect 2960 9220 2980 9260
rect 2900 9200 2980 9220
rect 3150 9260 3230 9280
rect 3150 9220 3170 9260
rect 3210 9220 3230 9260
rect 3150 9200 3230 9220
rect 3340 9260 3500 9280
rect 3340 9220 3360 9260
rect 3400 9220 3440 9260
rect 3480 9220 3500 9260
rect 3340 9200 3500 9220
rect 3630 9260 3710 9280
rect 3630 9220 3650 9260
rect 3690 9220 3710 9260
rect 3630 9200 3710 9220
rect 3960 9260 4040 9280
rect 3960 9220 3980 9260
rect 4020 9220 4040 9260
rect 3960 9200 4040 9220
rect 4400 9260 4480 9280
rect 4400 9220 4420 9260
rect 4460 9220 4480 9260
rect 4400 9200 4480 9220
rect 4790 9260 4870 9280
rect 4790 9220 4810 9260
rect 4850 9220 4870 9260
rect 4790 9200 4870 9220
rect 5180 9260 5260 9280
rect 5180 9220 5200 9260
rect 5240 9220 5260 9260
rect 5180 9200 5260 9220
rect 5860 9260 5940 9280
rect 5860 9220 5880 9260
rect 5920 9220 5940 9260
rect 9380 9270 9400 9310
rect 9440 9270 9460 9310
rect 9380 9250 9460 9270
rect 10080 9310 10160 9330
rect 10080 9270 10100 9310
rect 10140 9270 10160 9310
rect 10080 9250 10160 9270
rect 10750 9270 10770 9340
rect 10840 9270 10860 9340
rect 10750 9250 10860 9270
rect 5860 9200 5940 9220
rect 1280 9050 1320 9200
rect 1710 9150 1790 9170
rect 1710 9110 1730 9150
rect 1770 9110 1790 9150
rect 1710 9090 1790 9110
rect 1710 9050 1750 9090
rect 2020 9050 2060 9200
rect 2180 9050 2220 9200
rect 2920 9050 2960 9200
rect 3340 9050 3380 9200
rect 3650 9050 3690 9200
rect 3980 9050 4020 9200
rect 4420 9050 4460 9200
rect 4830 9150 4910 9160
rect 4830 9110 4850 9150
rect 4890 9110 4910 9150
rect 4830 9090 4910 9110
rect 5200 9050 5240 9200
rect 5470 9150 5550 9170
rect 5470 9110 5490 9150
rect 5530 9110 5550 9150
rect 5470 9090 5550 9110
rect 5490 9050 5530 9090
rect 1190 9030 1330 9050
rect 1190 8990 1200 9030
rect 1240 8990 1280 9030
rect 1320 8990 1330 9030
rect 1190 8930 1330 8990
rect 1190 8890 1200 8930
rect 1240 8890 1280 8930
rect 1320 8890 1330 8930
rect 1190 8830 1330 8890
rect 1190 8790 1200 8830
rect 1240 8790 1280 8830
rect 1320 8790 1330 8830
rect 1190 8730 1330 8790
rect 1190 8690 1200 8730
rect 1240 8690 1280 8730
rect 1320 8690 1330 8730
rect 1190 8670 1330 8690
rect 1380 9030 1440 9050
rect 1380 8990 1390 9030
rect 1430 8990 1440 9030
rect 1380 8930 1440 8990
rect 1380 8890 1390 8930
rect 1430 8890 1440 8930
rect 1380 8830 1440 8890
rect 1380 8790 1390 8830
rect 1430 8790 1440 8830
rect 1380 8730 1440 8790
rect 1380 8690 1390 8730
rect 1430 8690 1440 8730
rect 1380 8670 1440 8690
rect 1490 9030 1670 9050
rect 1490 8990 1500 9030
rect 1540 9000 1610 9030
rect 1540 8990 1550 9000
rect 1490 8930 1550 8990
rect 1590 8990 1610 9000
rect 1650 8990 1670 9030
rect 1590 8970 1670 8990
rect 1710 9030 1850 9050
rect 1710 9010 1800 9030
rect 1490 8890 1500 8930
rect 1540 8890 1550 8930
rect 1490 8830 1550 8890
rect 1490 8790 1500 8830
rect 1540 8790 1550 8830
rect 1490 8730 1550 8790
rect 1490 8690 1500 8730
rect 1540 8690 1550 8730
rect 1490 8670 1550 8690
rect 1500 8630 1540 8670
rect 1380 8590 1540 8630
rect 1140 8570 1220 8590
rect 1140 8530 1160 8570
rect 1200 8530 1220 8570
rect 1140 8510 1220 8530
rect 1380 8430 1420 8590
rect 1710 8550 1750 9010
rect 1790 8990 1800 9010
rect 1840 8990 1850 9030
rect 1790 8930 1850 8990
rect 1790 8890 1800 8930
rect 1840 8890 1850 8930
rect 1790 8830 1850 8890
rect 1790 8790 1800 8830
rect 1840 8790 1850 8830
rect 1790 8730 1850 8790
rect 1790 8690 1800 8730
rect 1840 8690 1850 8730
rect 1790 8670 1850 8690
rect 1900 9030 1960 9050
rect 1900 8990 1910 9030
rect 1950 8990 1960 9030
rect 1900 8930 1960 8990
rect 1900 8890 1910 8930
rect 1950 8890 1960 8930
rect 1900 8830 1960 8890
rect 1900 8790 1910 8830
rect 1950 8790 1960 8830
rect 1900 8730 1960 8790
rect 1900 8690 1910 8730
rect 1950 8690 1960 8730
rect 1900 8670 1960 8690
rect 2010 9030 2230 9050
rect 2010 8990 2020 9030
rect 2060 8990 2100 9030
rect 2140 8990 2180 9030
rect 2220 8990 2230 9030
rect 2010 8930 2230 8990
rect 2010 8890 2020 8930
rect 2060 8890 2100 8930
rect 2140 8890 2180 8930
rect 2220 8890 2230 8930
rect 2010 8830 2230 8890
rect 2010 8790 2020 8830
rect 2060 8790 2100 8830
rect 2140 8790 2180 8830
rect 2220 8790 2230 8830
rect 2010 8730 2230 8790
rect 2010 8690 2020 8730
rect 2060 8690 2100 8730
rect 2140 8690 2180 8730
rect 2220 8690 2230 8730
rect 2010 8670 2230 8690
rect 2280 9030 2340 9050
rect 2280 8990 2290 9030
rect 2330 8990 2340 9030
rect 2280 8930 2340 8990
rect 2280 8890 2290 8930
rect 2330 8890 2340 8930
rect 2280 8830 2340 8890
rect 2280 8790 2290 8830
rect 2330 8790 2340 8830
rect 2280 8730 2340 8790
rect 2280 8690 2290 8730
rect 2330 8690 2340 8730
rect 2280 8670 2340 8690
rect 2390 9030 2570 9050
rect 2390 8990 2400 9030
rect 2440 9000 2510 9030
rect 2440 8990 2450 9000
rect 2390 8930 2450 8990
rect 2490 8990 2510 9000
rect 2550 8990 2570 9030
rect 2490 8970 2570 8990
rect 2610 9030 2750 9050
rect 2610 9010 2700 9030
rect 2390 8890 2400 8930
rect 2440 8890 2450 8930
rect 2390 8830 2450 8890
rect 2390 8790 2400 8830
rect 2440 8790 2450 8830
rect 2390 8730 2450 8790
rect 2390 8690 2400 8730
rect 2440 8690 2450 8730
rect 2390 8670 2450 8690
rect 1800 8630 1840 8670
rect 2400 8630 2440 8670
rect 1800 8590 1950 8630
rect 1470 8530 1750 8550
rect 1470 8490 1490 8530
rect 1530 8510 1750 8530
rect 1530 8490 1550 8510
rect 1470 8470 1550 8490
rect 1910 8430 1950 8590
rect 1990 8610 2440 8630
rect 1990 8570 2010 8610
rect 2050 8590 2440 8610
rect 2050 8570 2070 8590
rect 1990 8550 2070 8570
rect 2280 8430 2320 8590
rect 2610 8550 2650 9010
rect 2690 8990 2700 9010
rect 2740 8990 2750 9030
rect 2690 8930 2750 8990
rect 2690 8890 2700 8930
rect 2740 8890 2750 8930
rect 2690 8830 2750 8890
rect 2690 8790 2700 8830
rect 2740 8790 2750 8830
rect 2690 8730 2750 8790
rect 2690 8690 2700 8730
rect 2740 8690 2750 8730
rect 2690 8670 2750 8690
rect 2800 9030 2860 9050
rect 2800 8990 2810 9030
rect 2850 8990 2860 9030
rect 2800 8930 2860 8990
rect 2800 8890 2810 8930
rect 2850 8890 2860 8930
rect 2800 8830 2860 8890
rect 2800 8790 2810 8830
rect 2850 8790 2860 8830
rect 2800 8730 2860 8790
rect 2800 8690 2810 8730
rect 2850 8690 2860 8730
rect 2800 8670 2860 8690
rect 2910 9030 3050 9050
rect 2910 8990 2920 9030
rect 2960 8990 3000 9030
rect 3040 8990 3050 9030
rect 2910 8930 3050 8990
rect 2910 8890 2920 8930
rect 2960 8890 3000 8930
rect 3040 8890 3050 8930
rect 2910 8830 3050 8890
rect 2910 8790 2920 8830
rect 2960 8790 3000 8830
rect 3040 8790 3050 8830
rect 2910 8730 3050 8790
rect 2910 8690 2920 8730
rect 2960 8690 3000 8730
rect 3040 8690 3050 8730
rect 2910 8670 3050 8690
rect 3200 9030 3260 9050
rect 3200 8990 3210 9030
rect 3250 8990 3260 9030
rect 3200 8930 3260 8990
rect 3200 8890 3210 8930
rect 3250 8890 3260 8930
rect 3200 8830 3260 8890
rect 3200 8790 3210 8830
rect 3250 8790 3260 8830
rect 3200 8730 3260 8790
rect 3200 8690 3210 8730
rect 3250 8690 3260 8730
rect 3200 8670 3260 8690
rect 3310 9030 3450 9050
rect 3310 8990 3320 9030
rect 3360 8990 3400 9030
rect 3440 8990 3450 9030
rect 3310 8930 3450 8990
rect 3310 8890 3320 8930
rect 3360 8890 3400 8930
rect 3440 8890 3450 8930
rect 3310 8830 3450 8890
rect 3310 8790 3320 8830
rect 3360 8790 3400 8830
rect 3440 8790 3450 8830
rect 3310 8730 3450 8790
rect 3310 8690 3320 8730
rect 3360 8690 3400 8730
rect 3440 8690 3450 8730
rect 3310 8670 3450 8690
rect 3530 9030 3590 9050
rect 3530 8990 3540 9030
rect 3580 8990 3590 9030
rect 3530 8930 3590 8990
rect 3530 8890 3540 8930
rect 3580 8890 3590 8930
rect 3530 8830 3590 8890
rect 3530 8790 3540 8830
rect 3580 8790 3590 8830
rect 3530 8730 3590 8790
rect 3530 8690 3540 8730
rect 3580 8690 3590 8730
rect 3530 8670 3590 8690
rect 3640 9030 3780 9050
rect 3640 8990 3650 9030
rect 3690 8990 3730 9030
rect 3770 8990 3780 9030
rect 3640 8930 3780 8990
rect 3640 8890 3650 8930
rect 3690 8890 3730 8930
rect 3770 8890 3780 8930
rect 3640 8830 3780 8890
rect 3640 8790 3650 8830
rect 3690 8790 3730 8830
rect 3770 8790 3780 8830
rect 3640 8730 3780 8790
rect 3640 8690 3650 8730
rect 3690 8690 3730 8730
rect 3770 8690 3780 8730
rect 3640 8670 3780 8690
rect 3860 9030 3920 9050
rect 3860 8990 3870 9030
rect 3910 8990 3920 9030
rect 3860 8930 3920 8990
rect 3860 8890 3870 8930
rect 3910 8890 3920 8930
rect 3860 8830 3920 8890
rect 3860 8790 3870 8830
rect 3910 8790 3920 8830
rect 3860 8730 3920 8790
rect 3860 8690 3870 8730
rect 3910 8690 3920 8730
rect 3860 8670 3920 8690
rect 3970 9030 4110 9050
rect 3970 8990 3980 9030
rect 4020 8990 4060 9030
rect 4100 8990 4110 9030
rect 3970 8930 4110 8990
rect 3970 8890 3980 8930
rect 4020 8890 4060 8930
rect 4100 8890 4110 8930
rect 3970 8830 4110 8890
rect 3970 8790 3980 8830
rect 4020 8790 4060 8830
rect 4100 8790 4110 8830
rect 3970 8730 4110 8790
rect 3970 8690 3980 8730
rect 4020 8690 4060 8730
rect 4100 8690 4110 8730
rect 3970 8670 4110 8690
rect 4300 9030 4480 9050
rect 4300 8990 4320 9030
rect 4360 8990 4420 9030
rect 4460 8990 4480 9030
rect 4300 8930 4480 8990
rect 4300 8890 4320 8930
rect 4360 8890 4420 8930
rect 4460 8890 4480 8930
rect 4300 8830 4480 8890
rect 4300 8790 4320 8830
rect 4360 8790 4420 8830
rect 4460 8790 4480 8830
rect 4300 8730 4480 8790
rect 4300 8690 4320 8730
rect 4360 8690 4420 8730
rect 4460 8690 4480 8730
rect 4300 8670 4480 8690
rect 4530 9030 4610 9050
rect 4530 8990 4550 9030
rect 4590 8990 4610 9030
rect 4530 8930 4610 8990
rect 4530 8890 4550 8930
rect 4590 8890 4610 8930
rect 4530 8830 4610 8890
rect 4530 8790 4550 8830
rect 4590 8790 4610 8830
rect 4530 8730 4610 8790
rect 4530 8690 4550 8730
rect 4590 8690 4610 8730
rect 4530 8670 4610 8690
rect 4790 9030 4870 9050
rect 4790 8990 4810 9030
rect 4850 8990 4870 9030
rect 4790 8930 4870 8990
rect 4790 8890 4810 8930
rect 4850 8890 4870 8930
rect 4790 8830 4870 8890
rect 4790 8790 4810 8830
rect 4850 8790 4870 8830
rect 4790 8730 4870 8790
rect 4790 8690 4810 8730
rect 4850 8690 4870 8730
rect 4790 8670 4870 8690
rect 4920 9030 5000 9050
rect 4920 8990 4940 9030
rect 4980 8990 5000 9030
rect 4920 8930 5000 8990
rect 4920 8890 4940 8930
rect 4980 8890 5000 8930
rect 4920 8830 5000 8890
rect 4920 8790 4940 8830
rect 4980 8790 5000 8830
rect 4920 8730 5000 8790
rect 4920 8690 4940 8730
rect 4980 8690 5000 8730
rect 4920 8670 5000 8690
rect 5080 9030 5260 9050
rect 5080 8990 5100 9030
rect 5140 8990 5200 9030
rect 5240 8990 5260 9030
rect 5080 8930 5260 8990
rect 5080 8890 5100 8930
rect 5140 8890 5200 8930
rect 5240 8890 5260 8930
rect 5080 8830 5260 8890
rect 5080 8790 5100 8830
rect 5140 8790 5200 8830
rect 5240 8790 5260 8830
rect 5080 8730 5260 8790
rect 5080 8690 5100 8730
rect 5140 8690 5200 8730
rect 5240 8690 5260 8730
rect 5080 8670 5260 8690
rect 5310 9030 5390 9050
rect 5310 8990 5330 9030
rect 5370 8990 5390 9030
rect 5310 8930 5390 8990
rect 5310 8890 5330 8930
rect 5370 8890 5390 8930
rect 5310 8830 5390 8890
rect 5310 8790 5330 8830
rect 5370 8790 5390 8830
rect 5310 8730 5390 8790
rect 5310 8690 5330 8730
rect 5370 8690 5390 8730
rect 5310 8670 5390 8690
rect 5470 9030 5550 9050
rect 5470 8990 5490 9030
rect 5530 8990 5550 9030
rect 5470 8930 5550 8990
rect 5470 8890 5490 8930
rect 5530 8890 5550 8930
rect 5470 8830 5550 8890
rect 5470 8790 5490 8830
rect 5530 8790 5550 8830
rect 5470 8730 5550 8790
rect 5470 8690 5490 8730
rect 5530 8690 5550 8730
rect 5470 8670 5550 8690
rect 5600 9030 5680 9050
rect 5600 8990 5620 9030
rect 5660 8990 5680 9030
rect 5600 8930 5680 8990
rect 5600 8890 5620 8930
rect 5660 8890 5680 8930
rect 5600 8830 5680 8890
rect 5600 8790 5620 8830
rect 5660 8790 5680 8830
rect 9820 8810 9900 8830
rect 5600 8730 5680 8790
rect 5600 8690 5620 8730
rect 5660 8690 5680 8730
rect 5600 8670 5680 8690
rect 7790 8770 7870 8790
rect 7790 8730 7810 8770
rect 7850 8730 7870 8770
rect 2700 8630 2740 8670
rect 2700 8590 2850 8630
rect 3200 8600 3240 8670
rect 3530 8600 3570 8670
rect 3860 8600 3900 8670
rect 4550 8630 4590 8670
rect 4810 8630 4850 8670
rect 2370 8530 2650 8550
rect 2370 8490 2390 8530
rect 2430 8510 2650 8530
rect 2430 8490 2450 8510
rect 2370 8470 2450 8490
rect 2810 8430 2850 8590
rect 3060 8580 3240 8600
rect 3060 8540 3080 8580
rect 3120 8540 3160 8580
rect 3200 8540 3240 8580
rect 3060 8520 3240 8540
rect 3470 8580 3570 8600
rect 3470 8540 3490 8580
rect 3530 8540 3570 8580
rect 3470 8520 3570 8540
rect 3800 8580 3900 8600
rect 3800 8540 3820 8580
rect 3860 8540 3900 8580
rect 3800 8520 3900 8540
rect 4090 8580 4170 8600
rect 4550 8590 4850 8630
rect 4090 8540 4110 8580
rect 4150 8540 4170 8580
rect 4090 8520 4170 8540
rect 4240 8570 4320 8590
rect 4240 8530 4260 8570
rect 4300 8530 4320 8570
rect 3200 8430 3240 8520
rect 3530 8430 3570 8520
rect 3860 8430 3900 8520
rect 4240 8510 4320 8530
rect 4550 8430 4590 8590
rect 4810 8430 4850 8590
rect 4940 8620 4980 8670
rect 4940 8600 5040 8620
rect 4940 8560 4980 8600
rect 5020 8560 5040 8600
rect 4940 8540 5040 8560
rect 4940 8430 4980 8540
rect 5350 8530 5390 8670
rect 5350 8520 5430 8530
rect 5350 8480 5370 8520
rect 5410 8480 5430 8520
rect 5350 8460 5430 8480
rect 5350 8430 5390 8460
rect 5490 8430 5530 8670
rect 5620 8550 5660 8670
rect 7250 8660 7430 8680
rect 7250 8620 7270 8660
rect 7310 8620 7370 8660
rect 7410 8620 7430 8660
rect 7250 8560 7430 8620
rect 5620 8530 6090 8550
rect 5620 8510 6030 8530
rect 5620 8430 5660 8510
rect 6010 8490 6030 8510
rect 6070 8490 6090 8530
rect 6010 8470 6090 8490
rect 7250 8520 7270 8560
rect 7310 8520 7370 8560
rect 7410 8520 7430 8560
rect 6010 8430 6050 8470
rect 7250 8460 7430 8520
rect 1190 8410 1330 8430
rect 1190 8370 1200 8410
rect 1240 8370 1280 8410
rect 1320 8370 1330 8410
rect 1190 8310 1330 8370
rect 1190 8270 1200 8310
rect 1240 8270 1280 8310
rect 1320 8270 1330 8310
rect 1190 8250 1330 8270
rect 1380 8410 1440 8430
rect 1380 8370 1390 8410
rect 1430 8370 1440 8410
rect 1380 8310 1440 8370
rect 1380 8270 1390 8310
rect 1430 8270 1440 8310
rect 1380 8250 1440 8270
rect 1490 8410 1550 8430
rect 1490 8370 1500 8410
rect 1540 8370 1550 8410
rect 1490 8310 1550 8370
rect 1490 8270 1500 8310
rect 1540 8270 1550 8310
rect 1490 8250 1550 8270
rect 1790 8410 1850 8430
rect 1790 8370 1800 8410
rect 1840 8370 1850 8410
rect 1790 8310 1850 8370
rect 1790 8270 1800 8310
rect 1840 8270 1850 8310
rect 1790 8250 1850 8270
rect 1900 8410 1960 8430
rect 1900 8370 1910 8410
rect 1950 8370 1960 8410
rect 1900 8310 1960 8370
rect 1900 8270 1910 8310
rect 1950 8270 1960 8310
rect 1900 8250 1960 8270
rect 2010 8410 2230 8430
rect 2010 8370 2020 8410
rect 2060 8370 2100 8410
rect 2140 8370 2180 8410
rect 2220 8370 2230 8410
rect 2010 8310 2230 8370
rect 2010 8270 2020 8310
rect 2060 8270 2100 8310
rect 2140 8270 2180 8310
rect 2220 8270 2230 8310
rect 2010 8250 2230 8270
rect 2280 8410 2340 8430
rect 2280 8370 2290 8410
rect 2330 8370 2340 8410
rect 2280 8310 2340 8370
rect 2280 8270 2290 8310
rect 2330 8270 2340 8310
rect 2280 8250 2340 8270
rect 2390 8410 2450 8430
rect 2390 8370 2400 8410
rect 2440 8370 2450 8410
rect 2390 8310 2450 8370
rect 2390 8270 2400 8310
rect 2440 8270 2450 8310
rect 2390 8250 2450 8270
rect 2690 8410 2750 8430
rect 2690 8370 2700 8410
rect 2740 8370 2750 8410
rect 2690 8310 2750 8370
rect 2690 8270 2700 8310
rect 2740 8270 2750 8310
rect 2690 8250 2750 8270
rect 2800 8410 2860 8430
rect 2800 8370 2810 8410
rect 2850 8370 2860 8410
rect 2800 8310 2860 8370
rect 2800 8270 2810 8310
rect 2850 8270 2860 8310
rect 2800 8250 2860 8270
rect 2910 8410 3050 8430
rect 2910 8370 2920 8410
rect 2960 8370 3000 8410
rect 3040 8370 3050 8410
rect 2910 8310 3050 8370
rect 2910 8270 2920 8310
rect 2960 8270 3000 8310
rect 3040 8270 3050 8310
rect 2910 8250 3050 8270
rect 3200 8410 3260 8430
rect 3200 8370 3210 8410
rect 3250 8370 3260 8410
rect 3200 8310 3260 8370
rect 3200 8270 3210 8310
rect 3250 8270 3260 8310
rect 3200 8250 3260 8270
rect 3310 8410 3450 8430
rect 3310 8370 3320 8410
rect 3360 8370 3400 8410
rect 3440 8370 3450 8410
rect 3310 8310 3450 8370
rect 3310 8270 3320 8310
rect 3360 8270 3400 8310
rect 3440 8270 3450 8310
rect 3310 8250 3450 8270
rect 3530 8410 3590 8430
rect 3530 8370 3540 8410
rect 3580 8370 3590 8410
rect 3530 8310 3590 8370
rect 3530 8270 3540 8310
rect 3580 8270 3590 8310
rect 3530 8250 3590 8270
rect 3640 8410 3780 8430
rect 3640 8370 3650 8410
rect 3690 8370 3730 8410
rect 3770 8370 3780 8410
rect 3640 8310 3780 8370
rect 3640 8270 3650 8310
rect 3690 8270 3730 8310
rect 3770 8270 3780 8310
rect 3640 8250 3780 8270
rect 3860 8410 3920 8430
rect 3860 8370 3870 8410
rect 3910 8370 3920 8410
rect 3860 8310 3920 8370
rect 3860 8270 3870 8310
rect 3910 8270 3920 8310
rect 3860 8250 3920 8270
rect 3970 8410 4110 8430
rect 3970 8370 3980 8410
rect 4020 8370 4060 8410
rect 4100 8370 4110 8410
rect 3970 8310 4110 8370
rect 3970 8270 3980 8310
rect 4020 8270 4060 8310
rect 4100 8270 4110 8310
rect 3970 8250 4110 8270
rect 4300 8410 4480 8430
rect 4300 8370 4320 8410
rect 4360 8370 4420 8410
rect 4460 8370 4480 8410
rect 4300 8310 4480 8370
rect 4300 8270 4320 8310
rect 4360 8270 4420 8310
rect 4460 8270 4480 8310
rect 4300 8250 4480 8270
rect 4530 8410 4610 8430
rect 4530 8370 4550 8410
rect 4590 8370 4610 8410
rect 4530 8310 4610 8370
rect 4530 8270 4550 8310
rect 4590 8270 4610 8310
rect 4530 8250 4610 8270
rect 4790 8410 4870 8430
rect 4790 8370 4810 8410
rect 4850 8370 4870 8410
rect 4790 8310 4870 8370
rect 4790 8270 4810 8310
rect 4850 8270 4870 8310
rect 4790 8250 4870 8270
rect 4920 8410 5000 8430
rect 4920 8370 4940 8410
rect 4980 8370 5000 8410
rect 4920 8310 5000 8370
rect 4920 8270 4940 8310
rect 4980 8270 5000 8310
rect 4920 8250 5000 8270
rect 5080 8410 5260 8430
rect 5080 8370 5100 8410
rect 5140 8370 5200 8410
rect 5240 8370 5260 8410
rect 5080 8310 5260 8370
rect 5080 8270 5100 8310
rect 5140 8270 5200 8310
rect 5240 8270 5260 8310
rect 5080 8250 5260 8270
rect 5310 8410 5390 8430
rect 5310 8370 5330 8410
rect 5370 8370 5390 8410
rect 5310 8310 5390 8370
rect 5310 8270 5330 8310
rect 5370 8270 5390 8310
rect 5310 8250 5390 8270
rect 5470 8410 5550 8430
rect 5470 8370 5490 8410
rect 5530 8370 5550 8410
rect 5470 8310 5550 8370
rect 5470 8270 5490 8310
rect 5530 8270 5550 8310
rect 5470 8250 5550 8270
rect 5600 8410 5680 8430
rect 5600 8370 5620 8410
rect 5660 8370 5680 8410
rect 5600 8310 5680 8370
rect 5600 8270 5620 8310
rect 5660 8270 5680 8310
rect 5600 8250 5680 8270
rect 5760 8410 5940 8430
rect 5760 8370 5780 8410
rect 5820 8370 5880 8410
rect 5920 8370 5940 8410
rect 5760 8310 5940 8370
rect 5760 8270 5780 8310
rect 5820 8270 5880 8310
rect 5920 8270 5940 8310
rect 5760 8250 5940 8270
rect 5990 8410 6070 8430
rect 5990 8370 6010 8410
rect 6050 8370 6070 8410
rect 5990 8310 6070 8370
rect 5990 8270 6010 8310
rect 6050 8270 6070 8310
rect 7250 8420 7270 8460
rect 7310 8420 7370 8460
rect 7410 8420 7430 8460
rect 7250 8360 7430 8420
rect 7250 8320 7270 8360
rect 7310 8320 7370 8360
rect 7410 8320 7430 8360
rect 7250 8300 7430 8320
rect 7570 8660 7650 8680
rect 7570 8620 7590 8660
rect 7630 8620 7650 8660
rect 7570 8560 7650 8620
rect 7570 8520 7590 8560
rect 7630 8520 7650 8560
rect 7570 8460 7650 8520
rect 7570 8420 7590 8460
rect 7630 8420 7650 8460
rect 7570 8360 7650 8420
rect 7570 8320 7590 8360
rect 7630 8320 7650 8360
rect 7570 8300 7650 8320
rect 7790 8660 7870 8730
rect 8330 8780 8410 8800
rect 8330 8740 8350 8780
rect 8390 8740 8410 8780
rect 8330 8680 8410 8740
rect 9410 8780 9490 8800
rect 9410 8740 9430 8780
rect 9470 8740 9490 8780
rect 9820 8770 9840 8810
rect 9880 8770 9900 8810
rect 9820 8750 9900 8770
rect 10080 8810 10160 8830
rect 10080 8770 10100 8810
rect 10140 8770 10160 8810
rect 10080 8750 10160 8770
rect 10750 8810 10860 8830
rect 9410 8680 9490 8740
rect 10750 8740 10770 8810
rect 10840 8740 10860 8810
rect 10750 8720 10860 8740
rect 7790 8620 7810 8660
rect 7850 8620 7870 8660
rect 7790 8560 7870 8620
rect 7790 8520 7810 8560
rect 7850 8520 7870 8560
rect 7790 8460 7870 8520
rect 7790 8420 7810 8460
rect 7850 8420 7870 8460
rect 7790 8360 7870 8420
rect 7790 8320 7810 8360
rect 7850 8320 7870 8360
rect 7790 8300 7870 8320
rect 8010 8660 8090 8680
rect 8010 8620 8030 8660
rect 8070 8620 8090 8660
rect 8010 8560 8090 8620
rect 8010 8520 8030 8560
rect 8070 8520 8090 8560
rect 8010 8460 8090 8520
rect 8010 8420 8030 8460
rect 8070 8420 8090 8460
rect 8010 8360 8090 8420
rect 8010 8320 8030 8360
rect 8070 8320 8090 8360
rect 8010 8300 8090 8320
rect 8230 8660 8510 8680
rect 8230 8620 8250 8660
rect 8290 8620 8350 8660
rect 8390 8620 8450 8660
rect 8490 8620 8510 8660
rect 8230 8560 8510 8620
rect 8230 8520 8250 8560
rect 8290 8520 8350 8560
rect 8390 8520 8450 8560
rect 8490 8520 8510 8560
rect 8230 8460 8510 8520
rect 8230 8420 8250 8460
rect 8290 8420 8350 8460
rect 8390 8420 8450 8460
rect 8490 8420 8510 8460
rect 8230 8360 8510 8420
rect 8230 8320 8250 8360
rect 8290 8320 8350 8360
rect 8390 8320 8450 8360
rect 8490 8320 8510 8360
rect 8230 8300 8510 8320
rect 8650 8660 8730 8680
rect 8650 8620 8670 8660
rect 8710 8620 8730 8660
rect 8650 8560 8730 8620
rect 8650 8520 8670 8560
rect 8710 8520 8730 8560
rect 8650 8460 8730 8520
rect 8650 8420 8670 8460
rect 8710 8420 8730 8460
rect 8650 8360 8730 8420
rect 8650 8320 8670 8360
rect 8710 8320 8730 8360
rect 8650 8300 8730 8320
rect 8870 8660 8950 8680
rect 8870 8620 8890 8660
rect 8930 8620 8950 8660
rect 8870 8560 8950 8620
rect 8870 8520 8890 8560
rect 8930 8520 8950 8560
rect 8870 8460 8950 8520
rect 8870 8420 8890 8460
rect 8930 8420 8950 8460
rect 8870 8360 8950 8420
rect 8870 8320 8890 8360
rect 8930 8320 8950 8360
rect 8870 8300 8950 8320
rect 9090 8660 9170 8680
rect 9090 8620 9110 8660
rect 9150 8620 9170 8660
rect 9090 8560 9170 8620
rect 9090 8520 9110 8560
rect 9150 8520 9170 8560
rect 9090 8460 9170 8520
rect 9090 8420 9110 8460
rect 9150 8420 9170 8460
rect 9090 8360 9170 8420
rect 9090 8320 9110 8360
rect 9150 8320 9170 8360
rect 9090 8300 9170 8320
rect 9310 8660 9590 8680
rect 9310 8620 9330 8660
rect 9370 8620 9430 8660
rect 9470 8620 9530 8660
rect 9570 8620 9590 8660
rect 9310 8560 9590 8620
rect 9310 8520 9330 8560
rect 9370 8520 9430 8560
rect 9470 8520 9530 8560
rect 9570 8520 9590 8560
rect 9310 8460 9590 8520
rect 9310 8420 9330 8460
rect 9370 8420 9430 8460
rect 9470 8420 9530 8460
rect 9570 8420 9590 8460
rect 9310 8360 9590 8420
rect 9310 8320 9330 8360
rect 9370 8320 9430 8360
rect 9470 8320 9530 8360
rect 9570 8320 9590 8360
rect 9310 8300 9590 8320
rect 9730 8660 9810 8680
rect 9730 8620 9750 8660
rect 9790 8620 9810 8660
rect 9730 8560 9810 8620
rect 9730 8520 9750 8560
rect 9790 8520 9810 8560
rect 9730 8460 9810 8520
rect 9730 8420 9750 8460
rect 9790 8420 9810 8460
rect 9730 8360 9810 8420
rect 9730 8320 9750 8360
rect 9790 8320 9810 8360
rect 9730 8300 9810 8320
rect 9950 8660 10030 8680
rect 9950 8620 9970 8660
rect 10010 8620 10030 8660
rect 9950 8560 10030 8620
rect 9950 8520 9970 8560
rect 10010 8520 10030 8560
rect 9950 8460 10030 8520
rect 9950 8420 9970 8460
rect 10010 8420 10030 8460
rect 9950 8360 10030 8420
rect 9950 8320 9970 8360
rect 10010 8320 10030 8360
rect 9950 8300 10030 8320
rect 10170 8660 10250 8680
rect 10170 8620 10190 8660
rect 10230 8620 10250 8660
rect 10170 8560 10250 8620
rect 10170 8520 10190 8560
rect 10230 8520 10250 8560
rect 10170 8460 10250 8520
rect 10170 8420 10190 8460
rect 10230 8420 10250 8460
rect 10170 8360 10250 8420
rect 10170 8320 10190 8360
rect 10230 8320 10250 8360
rect 10170 8300 10250 8320
rect 10390 8660 10570 8680
rect 10390 8620 10410 8660
rect 10450 8620 10510 8660
rect 10550 8620 10570 8660
rect 10390 8560 10570 8620
rect 10390 8520 10410 8560
rect 10450 8520 10510 8560
rect 10550 8520 10570 8560
rect 10390 8460 10570 8520
rect 10390 8420 10410 8460
rect 10450 8420 10510 8460
rect 10550 8420 10570 8460
rect 10390 8360 10570 8420
rect 10390 8320 10410 8360
rect 10450 8320 10510 8360
rect 10550 8320 10570 8360
rect 10390 8300 10570 8320
rect 5990 8250 6070 8270
rect 1280 8100 1320 8250
rect 1500 8100 1540 8250
rect 1800 8100 1840 8250
rect 2030 8100 2070 8250
rect 2180 8100 2220 8250
rect 2400 8100 2440 8250
rect 2700 8100 2740 8250
rect 2920 8100 2960 8250
rect 3320 8100 3360 8250
rect 3650 8100 3690 8250
rect 3980 8100 4020 8250
rect 4420 8100 4460 8250
rect 4910 8190 4990 8210
rect 4910 8150 4930 8190
rect 4970 8150 4990 8190
rect 4910 8130 4990 8150
rect 5200 8100 5240 8250
rect 5540 8190 5620 8210
rect 5540 8150 5560 8190
rect 5600 8150 5620 8190
rect 5540 8130 5620 8150
rect 5880 8100 5920 8250
rect 7350 8240 7430 8260
rect 7350 8200 7370 8240
rect 7410 8200 7430 8240
rect 7350 8180 7430 8200
rect 10390 8240 10470 8260
rect 10390 8200 10410 8240
rect 10450 8200 10470 8240
rect 10390 8180 10470 8200
rect 1260 8080 1340 8100
rect 1260 8040 1280 8080
rect 1320 8040 1340 8080
rect 1260 8020 1340 8040
rect 1480 8080 1560 8100
rect 1480 8040 1500 8080
rect 1540 8040 1560 8080
rect 1480 8020 1560 8040
rect 1780 8080 1860 8100
rect 1780 8040 1800 8080
rect 1840 8040 1860 8080
rect 1780 8020 1860 8040
rect 2010 8080 2090 8100
rect 2010 8040 2030 8080
rect 2070 8040 2090 8080
rect 2010 8020 2090 8040
rect 2160 8080 2240 8100
rect 2160 8040 2180 8080
rect 2220 8040 2240 8080
rect 2160 8020 2240 8040
rect 2380 8080 2460 8100
rect 2380 8040 2400 8080
rect 2440 8040 2460 8080
rect 2380 8020 2460 8040
rect 2680 8080 2760 8100
rect 2680 8040 2700 8080
rect 2740 8040 2760 8080
rect 2680 8020 2760 8040
rect 2900 8080 2980 8100
rect 2900 8040 2920 8080
rect 2960 8040 2980 8080
rect 2900 8020 2980 8040
rect 3300 8080 3380 8100
rect 3300 8040 3320 8080
rect 3360 8040 3380 8080
rect 3300 8020 3380 8040
rect 3630 8080 3710 8100
rect 3630 8040 3650 8080
rect 3690 8040 3710 8080
rect 3630 8020 3710 8040
rect 3960 8080 4040 8100
rect 3960 8040 3980 8080
rect 4020 8040 4040 8080
rect 3960 8020 4040 8040
rect 4400 8080 4480 8100
rect 4400 8040 4420 8080
rect 4460 8040 4480 8080
rect 4400 8020 4480 8040
rect 5180 8080 5260 8100
rect 5180 8040 5200 8080
rect 5240 8040 5260 8080
rect 5180 8020 5260 8040
rect 5860 8080 5940 8100
rect 5860 8040 5880 8080
rect 5920 8040 5940 8080
rect 5860 8020 5940 8040
rect 11100 8020 11210 8040
rect 11100 7950 11120 8020
rect 11190 7950 11210 8020
rect 11100 7930 11210 7950
rect 11220 7260 11320 7280
rect 11220 7200 11240 7260
rect 11300 7200 11320 7260
rect 11220 7180 11320 7200
rect -360 6960 -280 6980
rect -360 6920 -340 6960
rect -300 6920 -280 6960
rect -360 6900 -280 6920
rect 960 6960 1040 6980
rect 960 6920 980 6960
rect 1020 6920 1040 6960
rect 960 6900 1040 6920
rect 1540 6960 1620 6980
rect 1540 6920 1560 6960
rect 1600 6920 1620 6960
rect 1540 6900 1620 6920
rect 2860 6960 2940 6980
rect 2860 6920 2880 6960
rect 2920 6920 2940 6960
rect 2860 6900 2940 6920
rect -430 6840 -290 6860
rect -430 6800 -420 6840
rect -380 6800 -340 6840
rect -300 6800 -290 6840
rect -430 6740 -290 6800
rect -430 6700 -420 6740
rect -380 6700 -340 6740
rect -300 6700 -290 6740
rect -430 6680 -290 6700
rect -240 6840 -180 6860
rect -240 6800 -230 6840
rect -190 6800 -180 6840
rect -240 6740 -180 6800
rect -240 6700 -230 6740
rect -190 6700 -180 6740
rect -240 6680 -180 6700
rect -130 6840 -70 6860
rect -130 6800 -120 6840
rect -80 6800 -70 6840
rect -130 6740 -70 6800
rect -130 6700 -120 6740
rect -80 6700 -70 6740
rect -130 6680 -70 6700
rect -20 6840 40 6860
rect -20 6800 -10 6840
rect 30 6800 40 6840
rect -20 6740 40 6800
rect -20 6700 -10 6740
rect 30 6700 40 6740
rect -20 6680 40 6700
rect 90 6840 150 6860
rect 90 6800 100 6840
rect 140 6800 150 6840
rect 90 6740 150 6800
rect 90 6700 100 6740
rect 140 6700 150 6740
rect 90 6680 150 6700
rect 200 6840 260 6860
rect 200 6800 210 6840
rect 250 6800 260 6840
rect 200 6740 260 6800
rect 200 6700 210 6740
rect 250 6700 260 6740
rect 200 6680 260 6700
rect 310 6840 370 6860
rect 310 6800 320 6840
rect 360 6800 370 6840
rect 310 6740 370 6800
rect 310 6700 320 6740
rect 360 6700 370 6740
rect 310 6680 370 6700
rect 420 6840 480 6860
rect 420 6800 430 6840
rect 470 6800 480 6840
rect 420 6740 480 6800
rect 420 6700 430 6740
rect 470 6700 480 6740
rect 420 6680 480 6700
rect 530 6840 590 6860
rect 530 6800 540 6840
rect 580 6800 590 6840
rect 530 6740 590 6800
rect 530 6700 540 6740
rect 580 6700 590 6740
rect 530 6680 590 6700
rect 640 6840 700 6860
rect 640 6800 650 6840
rect 690 6800 700 6840
rect 640 6740 700 6800
rect 640 6700 650 6740
rect 690 6700 700 6740
rect 640 6680 700 6700
rect 750 6840 810 6860
rect 750 6800 760 6840
rect 800 6800 810 6840
rect 750 6740 810 6800
rect 750 6700 760 6740
rect 800 6700 810 6740
rect 750 6680 810 6700
rect 860 6840 920 6860
rect 860 6800 870 6840
rect 910 6800 920 6840
rect 860 6740 920 6800
rect 860 6700 870 6740
rect 910 6700 920 6740
rect 860 6680 920 6700
rect 970 6840 1110 6860
rect 970 6800 980 6840
rect 1020 6800 1060 6840
rect 1100 6800 1110 6840
rect 970 6740 1110 6800
rect 970 6700 980 6740
rect 1020 6700 1060 6740
rect 1100 6700 1110 6740
rect 970 6680 1110 6700
rect 1470 6840 1610 6860
rect 1470 6800 1480 6840
rect 1520 6800 1560 6840
rect 1600 6800 1610 6840
rect 1470 6740 1610 6800
rect 1470 6700 1480 6740
rect 1520 6700 1560 6740
rect 1600 6700 1610 6740
rect 1470 6680 1610 6700
rect 1660 6840 1720 6860
rect 1660 6800 1670 6840
rect 1710 6800 1720 6840
rect 1660 6740 1720 6800
rect 1660 6700 1670 6740
rect 1710 6700 1720 6740
rect 1660 6680 1720 6700
rect 1770 6840 1830 6860
rect 1770 6800 1780 6840
rect 1820 6800 1830 6840
rect 1770 6740 1830 6800
rect 1770 6700 1780 6740
rect 1820 6700 1830 6740
rect 1770 6680 1830 6700
rect 1880 6840 1940 6860
rect 1880 6800 1890 6840
rect 1930 6800 1940 6840
rect 1880 6740 1940 6800
rect 1880 6700 1890 6740
rect 1930 6700 1940 6740
rect 1880 6680 1940 6700
rect 1990 6840 2050 6860
rect 1990 6800 2000 6840
rect 2040 6800 2050 6840
rect 1990 6740 2050 6800
rect 1990 6700 2000 6740
rect 2040 6700 2050 6740
rect 1990 6680 2050 6700
rect 2100 6840 2160 6860
rect 2100 6800 2110 6840
rect 2150 6800 2160 6840
rect 2100 6740 2160 6800
rect 2100 6700 2110 6740
rect 2150 6700 2160 6740
rect 2100 6680 2160 6700
rect 2210 6840 2270 6860
rect 2210 6800 2220 6840
rect 2260 6800 2270 6840
rect 2210 6740 2270 6800
rect 2210 6700 2220 6740
rect 2260 6700 2270 6740
rect 2210 6680 2270 6700
rect 2320 6840 2380 6860
rect 2320 6800 2330 6840
rect 2370 6800 2380 6840
rect 2320 6740 2380 6800
rect 2320 6700 2330 6740
rect 2370 6700 2380 6740
rect 2320 6680 2380 6700
rect 2430 6840 2490 6860
rect 2430 6800 2440 6840
rect 2480 6800 2490 6840
rect 2430 6740 2490 6800
rect 2430 6700 2440 6740
rect 2480 6700 2490 6740
rect 2430 6680 2490 6700
rect 2540 6840 2600 6860
rect 2540 6800 2550 6840
rect 2590 6800 2600 6840
rect 2540 6740 2600 6800
rect 2540 6700 2550 6740
rect 2590 6700 2600 6740
rect 2540 6680 2600 6700
rect 2650 6840 2710 6860
rect 2650 6800 2660 6840
rect 2700 6800 2710 6840
rect 2650 6740 2710 6800
rect 2650 6700 2660 6740
rect 2700 6700 2710 6740
rect 2650 6680 2710 6700
rect 2760 6840 2820 6860
rect 2760 6800 2770 6840
rect 2810 6800 2820 6840
rect 2760 6740 2820 6800
rect 2760 6700 2770 6740
rect 2810 6700 2820 6740
rect 2760 6680 2820 6700
rect 2870 6840 3010 6860
rect 2870 6800 2880 6840
rect 2920 6800 2960 6840
rect 3000 6800 3010 6840
rect 2870 6740 3010 6800
rect 11043 6811 11139 6845
rect 11399 6811 11495 6845
rect 11043 6750 11077 6811
rect 2870 6700 2880 6740
rect 2920 6700 2960 6740
rect 3000 6700 3010 6740
rect 2870 6680 3010 6700
rect 11020 6749 11100 6750
rect 11020 6730 11043 6749
rect 11077 6730 11100 6749
rect 11020 6690 11040 6730
rect 11080 6690 11100 6730
rect 11461 6749 11495 6811
rect 11020 6670 11043 6690
rect -184 6622 -126 6640
rect -184 6588 -172 6622
rect -138 6588 -126 6622
rect -184 6570 -126 6588
rect -74 6622 -16 6640
rect -74 6588 -62 6622
rect -28 6588 -16 6622
rect -74 6570 -16 6588
rect 36 6622 94 6640
rect 36 6588 48 6622
rect 82 6588 94 6622
rect 36 6570 94 6588
rect 146 6622 204 6640
rect 146 6588 158 6622
rect 192 6588 204 6622
rect 146 6570 204 6588
rect 256 6622 314 6640
rect 256 6588 268 6622
rect 302 6588 314 6622
rect 256 6570 314 6588
rect 366 6622 424 6640
rect 366 6588 378 6622
rect 412 6588 424 6622
rect 366 6570 424 6588
rect 476 6622 534 6640
rect 476 6588 488 6622
rect 522 6588 534 6622
rect 476 6570 534 6588
rect 586 6622 644 6640
rect 586 6588 598 6622
rect 632 6588 644 6622
rect 586 6570 644 6588
rect 696 6622 754 6640
rect 696 6588 708 6622
rect 742 6588 754 6622
rect 696 6570 754 6588
rect 806 6622 864 6640
rect 806 6588 818 6622
rect 852 6588 864 6622
rect 806 6570 864 6588
rect 1716 6622 1774 6640
rect 1716 6588 1728 6622
rect 1762 6588 1774 6622
rect 1716 6570 1774 6588
rect 1826 6622 1884 6640
rect 1826 6588 1838 6622
rect 1872 6588 1884 6622
rect 1826 6570 1884 6588
rect 1936 6622 1994 6640
rect 1936 6588 1948 6622
rect 1982 6588 1994 6622
rect 1936 6570 1994 6588
rect 2046 6622 2104 6640
rect 2046 6588 2058 6622
rect 2092 6588 2104 6622
rect 2046 6570 2104 6588
rect 2156 6622 2214 6640
rect 2156 6588 2168 6622
rect 2202 6588 2214 6622
rect 2156 6570 2214 6588
rect 2266 6622 2324 6640
rect 2266 6588 2278 6622
rect 2312 6588 2324 6622
rect 2266 6570 2324 6588
rect 2376 6622 2434 6640
rect 2376 6588 2388 6622
rect 2422 6588 2434 6622
rect 2376 6570 2434 6588
rect 2486 6622 2544 6640
rect 2486 6588 2498 6622
rect 2532 6588 2544 6622
rect 2486 6570 2544 6588
rect 2596 6622 2654 6640
rect 2596 6588 2608 6622
rect 2642 6588 2654 6622
rect 2596 6570 2654 6588
rect 2706 6622 2764 6640
rect 2706 6588 2718 6622
rect 2752 6588 2764 6622
rect 2706 6570 2764 6588
rect -370 6360 -290 6380
rect -370 6320 -350 6360
rect -310 6320 -290 6360
rect -370 6300 -290 6320
rect -10 6360 70 6380
rect -10 6320 10 6360
rect 50 6320 70 6360
rect -10 6300 70 6320
rect 350 6360 430 6380
rect 350 6320 370 6360
rect 410 6320 430 6360
rect 350 6300 430 6320
rect 710 6360 790 6380
rect 710 6320 730 6360
rect 770 6320 790 6360
rect 710 6300 790 6320
rect 1070 6360 1150 6380
rect 1070 6320 1090 6360
rect 1130 6320 1150 6360
rect 1070 6300 1150 6320
rect 1430 6360 1510 6380
rect 1430 6320 1450 6360
rect 1490 6320 1510 6360
rect 1430 6300 1510 6320
rect 1790 6360 1870 6380
rect 1790 6320 1810 6360
rect 1850 6320 1870 6360
rect 1790 6300 1870 6320
rect 2150 6360 2230 6380
rect 2150 6320 2170 6360
rect 2210 6320 2230 6360
rect 2150 6300 2230 6320
rect 2510 6360 2590 6380
rect 2510 6320 2530 6360
rect 2570 6320 2590 6360
rect 2510 6300 2590 6320
rect 2870 6360 2950 6380
rect 2870 6320 2890 6360
rect 2930 6320 2950 6360
rect 2870 6300 2950 6320
rect 7150 6356 7270 6360
rect 8570 6356 8690 6360
rect 7150 6340 7304 6356
rect 7150 6300 7170 6340
rect 7210 6306 7270 6340
rect 7210 6300 7304 6306
rect -350 6260 -310 6300
rect 10 6260 50 6300
rect 370 6260 410 6300
rect 730 6260 770 6300
rect 1090 6260 1130 6300
rect 1450 6260 1490 6300
rect 1810 6260 1850 6300
rect 2170 6260 2210 6300
rect 2530 6260 2570 6300
rect 2890 6260 2930 6300
rect 7150 6290 7304 6300
rect 8544 6340 8690 6356
rect 8578 6306 8690 6340
rect 8544 6290 8690 6306
rect 7150 6280 7270 6290
rect -440 6240 -300 6260
rect -440 6200 -430 6240
rect -390 6200 -350 6240
rect -310 6200 -300 6240
rect -440 6140 -300 6200
rect -440 6100 -430 6140
rect -390 6100 -350 6140
rect -310 6100 -300 6140
rect -440 6040 -300 6100
rect -440 6000 -430 6040
rect -390 6000 -350 6040
rect -310 6000 -300 6040
rect -440 5940 -300 6000
rect -440 5900 -430 5940
rect -390 5900 -350 5940
rect -310 5900 -300 5940
rect -440 5840 -300 5900
rect -440 5800 -430 5840
rect -390 5800 -350 5840
rect -310 5800 -300 5840
rect -440 5740 -300 5800
rect -440 5700 -430 5740
rect -390 5700 -350 5740
rect -310 5700 -300 5740
rect -440 5680 -300 5700
rect -180 6240 -120 6260
rect -180 6200 -170 6240
rect -130 6200 -120 6240
rect -180 6140 -120 6200
rect -180 6100 -170 6140
rect -130 6100 -120 6140
rect -180 6040 -120 6100
rect -180 6000 -170 6040
rect -130 6000 -120 6040
rect -180 5940 -120 6000
rect -180 5900 -170 5940
rect -130 5900 -120 5940
rect -180 5840 -120 5900
rect -180 5800 -170 5840
rect -130 5800 -120 5840
rect -180 5740 -120 5800
rect -180 5700 -170 5740
rect -130 5700 -120 5740
rect -180 5680 -120 5700
rect 0 6240 60 6260
rect 0 6200 10 6240
rect 50 6200 60 6240
rect 0 6140 60 6200
rect 0 6100 10 6140
rect 50 6100 60 6140
rect 0 6040 60 6100
rect 0 6000 10 6040
rect 50 6000 60 6040
rect 0 5940 60 6000
rect 0 5900 10 5940
rect 50 5900 60 5940
rect 0 5840 60 5900
rect 0 5800 10 5840
rect 50 5800 60 5840
rect 0 5740 60 5800
rect 0 5700 10 5740
rect 50 5700 60 5740
rect 0 5680 60 5700
rect 180 6240 240 6260
rect 180 6200 190 6240
rect 230 6200 240 6240
rect 180 6140 240 6200
rect 180 6100 190 6140
rect 230 6100 240 6140
rect 180 6040 240 6100
rect 180 6000 190 6040
rect 230 6000 240 6040
rect 180 5940 240 6000
rect 180 5900 190 5940
rect 230 5900 240 5940
rect 180 5840 240 5900
rect 180 5800 190 5840
rect 230 5800 240 5840
rect 180 5740 240 5800
rect 180 5700 190 5740
rect 230 5700 240 5740
rect 180 5680 240 5700
rect 360 6240 420 6260
rect 360 6200 370 6240
rect 410 6200 420 6240
rect 360 6140 420 6200
rect 360 6100 370 6140
rect 410 6100 420 6140
rect 360 6040 420 6100
rect 360 6000 370 6040
rect 410 6000 420 6040
rect 360 5940 420 6000
rect 360 5900 370 5940
rect 410 5900 420 5940
rect 360 5840 420 5900
rect 360 5800 370 5840
rect 410 5800 420 5840
rect 360 5740 420 5800
rect 360 5700 370 5740
rect 410 5700 420 5740
rect 360 5680 420 5700
rect 540 6240 600 6260
rect 540 6200 550 6240
rect 590 6200 600 6240
rect 540 6140 600 6200
rect 540 6100 550 6140
rect 590 6100 600 6140
rect 540 6040 600 6100
rect 540 6000 550 6040
rect 590 6000 600 6040
rect 540 5940 600 6000
rect 540 5900 550 5940
rect 590 5900 600 5940
rect 540 5840 600 5900
rect 540 5800 550 5840
rect 590 5800 600 5840
rect 540 5740 600 5800
rect 540 5700 550 5740
rect 590 5700 600 5740
rect 540 5680 600 5700
rect 720 6240 780 6260
rect 720 6200 730 6240
rect 770 6200 780 6240
rect 720 6140 780 6200
rect 720 6100 730 6140
rect 770 6100 780 6140
rect 720 6040 780 6100
rect 720 6000 730 6040
rect 770 6000 780 6040
rect 720 5940 780 6000
rect 720 5900 730 5940
rect 770 5900 780 5940
rect 720 5840 780 5900
rect 720 5800 730 5840
rect 770 5800 780 5840
rect 720 5740 780 5800
rect 720 5700 730 5740
rect 770 5700 780 5740
rect 720 5680 780 5700
rect 900 6240 960 6260
rect 900 6200 910 6240
rect 950 6200 960 6240
rect 900 6140 960 6200
rect 900 6100 910 6140
rect 950 6100 960 6140
rect 900 6040 960 6100
rect 900 6000 910 6040
rect 950 6000 960 6040
rect 900 5940 960 6000
rect 900 5900 910 5940
rect 950 5900 960 5940
rect 900 5840 960 5900
rect 900 5800 910 5840
rect 950 5800 960 5840
rect 900 5740 960 5800
rect 900 5700 910 5740
rect 950 5700 960 5740
rect 900 5680 960 5700
rect 1080 6240 1140 6260
rect 1080 6200 1090 6240
rect 1130 6200 1140 6240
rect 1080 6140 1140 6200
rect 1080 6100 1090 6140
rect 1130 6100 1140 6140
rect 1080 6040 1140 6100
rect 1080 6000 1090 6040
rect 1130 6000 1140 6040
rect 1080 5940 1140 6000
rect 1080 5900 1090 5940
rect 1130 5900 1140 5940
rect 1080 5840 1140 5900
rect 1080 5800 1090 5840
rect 1130 5800 1140 5840
rect 1080 5740 1140 5800
rect 1080 5700 1090 5740
rect 1130 5700 1140 5740
rect 1080 5680 1140 5700
rect 1260 6240 1320 6260
rect 1260 6200 1270 6240
rect 1310 6200 1320 6240
rect 1260 6140 1320 6200
rect 1260 6100 1270 6140
rect 1310 6100 1320 6140
rect 1260 6040 1320 6100
rect 1260 6000 1270 6040
rect 1310 6000 1320 6040
rect 1260 5940 1320 6000
rect 1260 5900 1270 5940
rect 1310 5900 1320 5940
rect 1260 5840 1320 5900
rect 1260 5800 1270 5840
rect 1310 5800 1320 5840
rect 1260 5740 1320 5800
rect 1260 5700 1270 5740
rect 1310 5700 1320 5740
rect 1260 5680 1320 5700
rect 1440 6240 1500 6260
rect 1440 6200 1450 6240
rect 1490 6200 1500 6240
rect 1440 6140 1500 6200
rect 1440 6100 1450 6140
rect 1490 6100 1500 6140
rect 1440 6040 1500 6100
rect 1440 6000 1450 6040
rect 1490 6000 1500 6040
rect 1440 5940 1500 6000
rect 1440 5900 1450 5940
rect 1490 5900 1500 5940
rect 1440 5840 1500 5900
rect 1440 5800 1450 5840
rect 1490 5800 1500 5840
rect 1440 5740 1500 5800
rect 1440 5700 1450 5740
rect 1490 5700 1500 5740
rect 1440 5680 1500 5700
rect 1620 6240 1680 6260
rect 1620 6200 1630 6240
rect 1670 6200 1680 6240
rect 1620 6140 1680 6200
rect 1620 6100 1630 6140
rect 1670 6100 1680 6140
rect 1620 6040 1680 6100
rect 1620 6000 1630 6040
rect 1670 6000 1680 6040
rect 1620 5940 1680 6000
rect 1620 5900 1630 5940
rect 1670 5900 1680 5940
rect 1620 5840 1680 5900
rect 1620 5800 1630 5840
rect 1670 5800 1680 5840
rect 1620 5740 1680 5800
rect 1620 5700 1630 5740
rect 1670 5700 1680 5740
rect 1620 5680 1680 5700
rect 1800 6240 1860 6260
rect 1800 6200 1810 6240
rect 1850 6200 1860 6240
rect 1800 6140 1860 6200
rect 1800 6100 1810 6140
rect 1850 6100 1860 6140
rect 1800 6040 1860 6100
rect 1800 6000 1810 6040
rect 1850 6000 1860 6040
rect 1800 5940 1860 6000
rect 1800 5900 1810 5940
rect 1850 5900 1860 5940
rect 1800 5840 1860 5900
rect 1800 5800 1810 5840
rect 1850 5800 1860 5840
rect 1800 5740 1860 5800
rect 1800 5700 1810 5740
rect 1850 5700 1860 5740
rect 1800 5680 1860 5700
rect 1980 6240 2040 6260
rect 1980 6200 1990 6240
rect 2030 6200 2040 6240
rect 1980 6140 2040 6200
rect 1980 6100 1990 6140
rect 2030 6100 2040 6140
rect 1980 6040 2040 6100
rect 1980 6000 1990 6040
rect 2030 6000 2040 6040
rect 1980 5940 2040 6000
rect 1980 5900 1990 5940
rect 2030 5900 2040 5940
rect 1980 5840 2040 5900
rect 1980 5800 1990 5840
rect 2030 5800 2040 5840
rect 1980 5740 2040 5800
rect 1980 5700 1990 5740
rect 2030 5700 2040 5740
rect 1980 5680 2040 5700
rect 2160 6240 2220 6260
rect 2160 6200 2170 6240
rect 2210 6200 2220 6240
rect 2160 6140 2220 6200
rect 2160 6100 2170 6140
rect 2210 6100 2220 6140
rect 2160 6040 2220 6100
rect 2160 6000 2170 6040
rect 2210 6000 2220 6040
rect 2160 5940 2220 6000
rect 2160 5900 2170 5940
rect 2210 5900 2220 5940
rect 2160 5840 2220 5900
rect 2160 5800 2170 5840
rect 2210 5800 2220 5840
rect 2160 5740 2220 5800
rect 2160 5700 2170 5740
rect 2210 5700 2220 5740
rect 2160 5680 2220 5700
rect 2340 6240 2400 6260
rect 2340 6200 2350 6240
rect 2390 6200 2400 6240
rect 2340 6140 2400 6200
rect 2340 6100 2350 6140
rect 2390 6100 2400 6140
rect 2340 6040 2400 6100
rect 2340 6000 2350 6040
rect 2390 6000 2400 6040
rect 2340 5940 2400 6000
rect 2340 5900 2350 5940
rect 2390 5900 2400 5940
rect 2340 5840 2400 5900
rect 2340 5800 2350 5840
rect 2390 5800 2400 5840
rect 2340 5740 2400 5800
rect 2340 5700 2350 5740
rect 2390 5700 2400 5740
rect 2340 5680 2400 5700
rect 2520 6240 2580 6260
rect 2520 6200 2530 6240
rect 2570 6200 2580 6240
rect 2520 6140 2580 6200
rect 2520 6100 2530 6140
rect 2570 6100 2580 6140
rect 2520 6040 2580 6100
rect 2520 6000 2530 6040
rect 2570 6000 2580 6040
rect 2520 5940 2580 6000
rect 2520 5900 2530 5940
rect 2570 5900 2580 5940
rect 2520 5840 2580 5900
rect 2520 5800 2530 5840
rect 2570 5800 2580 5840
rect 2520 5740 2580 5800
rect 2520 5700 2530 5740
rect 2570 5700 2580 5740
rect 2520 5680 2580 5700
rect 2700 6240 2760 6260
rect 2700 6200 2710 6240
rect 2750 6200 2760 6240
rect 2700 6140 2760 6200
rect 2700 6100 2710 6140
rect 2750 6100 2760 6140
rect 2700 6040 2760 6100
rect 2700 6000 2710 6040
rect 2750 6000 2760 6040
rect 2700 5940 2760 6000
rect 2700 5900 2710 5940
rect 2750 5900 2760 5940
rect 2700 5840 2760 5900
rect 2700 5800 2710 5840
rect 2750 5800 2760 5840
rect 2700 5740 2760 5800
rect 2700 5700 2710 5740
rect 2750 5700 2760 5740
rect 2700 5680 2760 5700
rect 2880 6240 3020 6260
rect 2880 6200 2890 6240
rect 2930 6200 2970 6240
rect 3010 6200 3020 6240
rect 2880 6140 3020 6200
rect 2880 6100 2890 6140
rect 2930 6100 2970 6140
rect 3010 6100 3020 6140
rect 3500 6160 3580 6180
rect 3500 6120 3520 6160
rect 3560 6120 3580 6160
rect 3500 6100 3580 6120
rect 3720 6160 3800 6180
rect 3720 6120 3740 6160
rect 3780 6120 3800 6160
rect 3720 6100 3800 6120
rect 3950 6160 4010 6180
rect 8600 6170 8690 6290
rect 3950 6120 3960 6160
rect 4000 6120 4010 6160
rect 3950 6100 4010 6120
rect 8210 6150 8690 6170
rect 8210 6110 8230 6150
rect 8270 6110 8630 6150
rect 8670 6110 8690 6150
rect 2880 6040 3020 6100
rect 8210 6090 8690 6110
rect 2880 6000 2890 6040
rect 2930 6000 2970 6040
rect 3010 6000 3020 6040
rect 2880 5940 3020 6000
rect 2880 5900 2890 5940
rect 2930 5900 2970 5940
rect 3010 5900 3020 5940
rect 2880 5840 3020 5900
rect 3420 6040 3570 6060
rect 3420 6000 3430 6040
rect 3470 6000 3520 6040
rect 3560 6000 3570 6040
rect 3420 5940 3570 6000
rect 3420 5900 3430 5940
rect 3470 5900 3520 5940
rect 3560 5900 3570 5940
rect 3420 5880 3570 5900
rect 3620 6040 3680 6060
rect 3620 6000 3630 6040
rect 3670 6000 3680 6040
rect 3620 5940 3680 6000
rect 3620 5900 3630 5940
rect 3670 5900 3680 5940
rect 3620 5880 3680 5900
rect 3730 6040 3790 6060
rect 3730 6000 3740 6040
rect 3780 6000 3790 6040
rect 3730 5940 3790 6000
rect 3730 5900 3740 5940
rect 3780 5900 3790 5940
rect 3730 5880 3790 5900
rect 3840 6040 3900 6060
rect 3840 6000 3850 6040
rect 3890 6000 3900 6040
rect 3840 5940 3900 6000
rect 3840 5900 3850 5940
rect 3890 5900 3900 5940
rect 3840 5880 3900 5900
rect 3950 6040 4090 6060
rect 8230 6050 8270 6090
rect 8630 6050 8670 6090
rect 3950 6000 3960 6040
rect 4000 6000 4040 6040
rect 4080 6000 4090 6040
rect 3950 5940 4090 6000
rect 3950 5900 3960 5940
rect 4000 5900 4040 5940
rect 4080 5900 4090 5940
rect 3950 5880 4090 5900
rect 7310 6030 7490 6050
rect 7310 5980 7330 6030
rect 7370 5980 7430 6030
rect 7470 5980 7490 6030
rect 7310 5890 7490 5980
rect 7310 5840 7330 5890
rect 7370 5840 7430 5890
rect 7470 5840 7490 5890
rect 2880 5800 2890 5840
rect 2930 5800 2970 5840
rect 3010 5800 3020 5840
rect 2880 5740 3020 5800
rect 3600 5820 3680 5840
rect 3600 5780 3620 5820
rect 3660 5780 3680 5820
rect 3600 5760 3680 5780
rect 3720 5820 3800 5840
rect 3720 5780 3740 5820
rect 3780 5780 3800 5820
rect 3720 5760 3800 5780
rect 3840 5820 3920 5840
rect 7310 5820 7490 5840
rect 7610 6030 7690 6050
rect 7610 5980 7630 6030
rect 7670 5980 7690 6030
rect 7610 5890 7690 5980
rect 7610 5840 7630 5890
rect 7670 5840 7690 5890
rect 7610 5820 7690 5840
rect 7810 6030 7890 6050
rect 7810 5980 7830 6030
rect 7870 5980 7890 6030
rect 7810 5890 7890 5980
rect 7810 5840 7830 5890
rect 7870 5840 7890 5890
rect 7810 5820 7890 5840
rect 8010 6030 8090 6050
rect 8010 5980 8030 6030
rect 8070 5980 8090 6030
rect 8010 5890 8090 5980
rect 8010 5840 8030 5890
rect 8070 5840 8090 5890
rect 8010 5820 8090 5840
rect 8210 6030 8290 6050
rect 8210 5980 8230 6030
rect 8270 5980 8290 6030
rect 8210 5890 8290 5980
rect 8210 5840 8230 5890
rect 8270 5840 8290 5890
rect 8210 5820 8290 5840
rect 8410 6030 8490 6050
rect 8410 5980 8430 6030
rect 8470 5980 8490 6030
rect 8410 5890 8490 5980
rect 8410 5840 8430 5890
rect 8470 5840 8490 5890
rect 8410 5820 8490 5840
rect 8610 6030 8690 6050
rect 8610 5980 8630 6030
rect 8670 5980 8690 6030
rect 8610 5890 8690 5980
rect 8610 5840 8630 5890
rect 8670 5840 8690 5890
rect 8610 5820 8690 5840
rect 8810 6030 8890 6050
rect 8810 5980 8830 6030
rect 8870 5980 8890 6030
rect 8810 5890 8890 5980
rect 8810 5840 8830 5890
rect 8870 5840 8890 5890
rect 8810 5820 8890 5840
rect 9010 6030 9090 6050
rect 9010 5980 9030 6030
rect 9070 5980 9090 6030
rect 9010 5890 9090 5980
rect 9010 5840 9030 5890
rect 9070 5840 9090 5890
rect 9010 5820 9090 5840
rect 9210 6030 9290 6050
rect 9210 5980 9230 6030
rect 9270 5980 9290 6030
rect 9210 5890 9290 5980
rect 9210 5840 9230 5890
rect 9270 5840 9290 5890
rect 9210 5820 9290 5840
rect 9410 6030 9590 6050
rect 9410 5980 9430 6030
rect 9470 5980 9530 6030
rect 9570 5980 9590 6030
rect 9410 5890 9590 5980
rect 9410 5840 9430 5890
rect 9470 5840 9530 5890
rect 9570 5840 9590 5890
rect 9410 5820 9590 5840
rect 3840 5780 3860 5820
rect 3900 5780 3920 5820
rect 7430 5780 7470 5820
rect 7830 5780 7870 5820
rect 9030 5780 9070 5820
rect 9430 5780 9470 5820
rect 3840 5760 3920 5780
rect 7410 5760 7490 5780
rect 2880 5700 2890 5740
rect 2930 5700 2970 5740
rect 3010 5700 3020 5740
rect 7410 5720 7430 5760
rect 7470 5720 7490 5760
rect 7830 5740 9070 5780
rect 7410 5700 7490 5720
rect 8990 5720 9070 5740
rect 2880 5680 3020 5700
rect 8990 5680 9010 5720
rect 9050 5680 9070 5720
rect 9410 5760 9490 5780
rect 9410 5720 9430 5760
rect 9470 5720 9490 5760
rect 9410 5700 9490 5720
rect 8990 5660 9070 5680
rect 11077 6670 11100 6690
rect -90 5620 -20 5640
rect -90 5580 -80 5620
rect -40 5580 -20 5620
rect -90 5560 -20 5580
rect 80 5620 160 5640
rect 80 5580 100 5620
rect 140 5580 160 5620
rect 80 5560 160 5580
rect 260 5620 340 5640
rect 260 5580 280 5620
rect 320 5580 340 5620
rect 260 5560 340 5580
rect 440 5620 520 5640
rect 440 5580 460 5620
rect 500 5580 520 5620
rect 440 5560 520 5580
rect 620 5620 700 5640
rect 620 5580 640 5620
rect 680 5580 700 5620
rect 620 5560 700 5580
rect 800 5620 880 5640
rect 800 5580 820 5620
rect 860 5580 880 5620
rect 800 5560 880 5580
rect 980 5620 1060 5640
rect 980 5580 1000 5620
rect 1040 5580 1060 5620
rect 980 5560 1060 5580
rect 1160 5620 1230 5640
rect 1160 5580 1180 5620
rect 1220 5580 1230 5620
rect 1160 5560 1230 5580
rect 1350 5620 1420 5640
rect 1350 5580 1360 5620
rect 1400 5580 1420 5620
rect 1350 5560 1420 5580
rect 1520 5620 1600 5640
rect 1520 5580 1540 5620
rect 1580 5580 1600 5620
rect 1520 5560 1600 5580
rect 1700 5620 1780 5640
rect 1700 5580 1720 5620
rect 1760 5580 1780 5620
rect 1700 5560 1780 5580
rect 1880 5620 1960 5640
rect 1880 5580 1900 5620
rect 1940 5580 1960 5620
rect 1880 5560 1960 5580
rect 2060 5620 2140 5640
rect 2060 5580 2080 5620
rect 2120 5580 2140 5620
rect 2060 5560 2140 5580
rect 2240 5620 2320 5640
rect 2240 5580 2260 5620
rect 2300 5580 2320 5620
rect 2240 5560 2320 5580
rect 2420 5620 2500 5640
rect 2420 5580 2440 5620
rect 2480 5580 2500 5620
rect 2420 5560 2500 5580
rect 2600 5620 2670 5640
rect 2600 5580 2620 5620
rect 2660 5580 2670 5620
rect 2600 5560 2670 5580
rect 7850 5610 7930 5630
rect 7850 5570 7870 5610
rect 7910 5570 7930 5610
rect 7850 5550 7930 5570
rect 10130 5610 10210 5630
rect 10130 5570 10150 5610
rect 10190 5570 10210 5610
rect 10130 5550 10210 5570
rect 11043 5597 11077 5659
rect 11461 5597 11495 5659
rect 11043 5563 11139 5597
rect 11399 5563 11495 5597
rect 7520 5470 7610 5490
rect 7520 5440 7540 5470
rect 7480 5420 7540 5440
rect 7590 5440 7610 5470
rect 7870 5440 7910 5550
rect 8990 5500 9070 5520
rect 8170 5470 8260 5490
rect 8170 5440 8190 5470
rect 7590 5420 8190 5440
rect 8240 5440 8260 5470
rect 8660 5460 8740 5480
rect 8660 5440 8680 5460
rect 8240 5420 8300 5440
rect 7480 5400 8300 5420
rect 7480 5360 7520 5400
rect 7610 5360 7650 5400
rect 7870 5360 7910 5400
rect 8130 5360 8170 5400
rect 8260 5360 8300 5400
rect 8620 5420 8680 5440
rect 8720 5440 8740 5460
rect 8990 5460 9010 5500
rect 9050 5460 9070 5500
rect 8990 5440 9070 5460
rect 9320 5460 9400 5480
rect 9320 5440 9340 5460
rect 8720 5420 9340 5440
rect 9380 5440 9400 5460
rect 9800 5460 9880 5480
rect 9800 5450 9820 5460
rect 9380 5420 9440 5440
rect 8620 5400 9440 5420
rect 8620 5360 8660 5400
rect 8750 5360 8790 5400
rect 9010 5360 9050 5400
rect 9270 5360 9310 5400
rect 9400 5360 9440 5400
rect 9760 5420 9820 5450
rect 9860 5450 9880 5460
rect 10150 5450 10190 5550
rect 10460 5460 10540 5480
rect 10460 5450 10480 5460
rect 9860 5420 10480 5450
rect 10520 5450 10540 5460
rect 10520 5420 10580 5450
rect 9760 5400 10580 5420
rect 9760 5360 9800 5400
rect 9890 5360 9930 5400
rect 10150 5360 10190 5400
rect 10410 5360 10450 5400
rect 10540 5360 10580 5400
rect 7360 5340 7540 5360
rect 7360 5300 7380 5340
rect 7420 5300 7480 5340
rect 7520 5300 7540 5340
rect 7360 5280 7540 5300
rect 7590 5340 7670 5360
rect 7590 5300 7610 5340
rect 7650 5300 7670 5340
rect 7590 5280 7670 5300
rect 7720 5340 7800 5360
rect 7720 5300 7740 5340
rect 7780 5300 7800 5340
rect 7720 5280 7800 5300
rect 7850 5340 7930 5360
rect 7850 5300 7870 5340
rect 7910 5300 7930 5340
rect 7850 5280 7930 5300
rect 7980 5340 8060 5360
rect 7980 5300 8000 5340
rect 8040 5300 8060 5340
rect 7980 5280 8060 5300
rect 8110 5340 8190 5360
rect 8110 5300 8130 5340
rect 8170 5300 8190 5340
rect 8110 5280 8190 5300
rect 8240 5340 8420 5360
rect 8240 5300 8260 5340
rect 8300 5300 8360 5340
rect 8400 5300 8420 5340
rect 8240 5280 8420 5300
rect 8600 5340 8680 5360
rect 8600 5300 8620 5340
rect 8660 5300 8680 5340
rect 8600 5280 8680 5300
rect 8730 5340 8810 5360
rect 8730 5300 8750 5340
rect 8790 5300 8810 5340
rect 8730 5280 8810 5300
rect 8860 5340 8940 5360
rect 8860 5300 8880 5340
rect 8920 5300 8940 5340
rect 8860 5280 8940 5300
rect 8990 5340 9070 5360
rect 8990 5300 9010 5340
rect 9050 5300 9070 5340
rect 8990 5280 9070 5300
rect 9120 5340 9200 5360
rect 9120 5300 9140 5340
rect 9180 5300 9200 5340
rect 9120 5280 9200 5300
rect 9250 5340 9330 5360
rect 9250 5300 9270 5340
rect 9310 5300 9330 5340
rect 9250 5280 9330 5300
rect 9380 5340 9460 5360
rect 9380 5300 9400 5340
rect 9440 5300 9460 5340
rect 9380 5280 9460 5300
rect 9640 5340 9820 5360
rect 9640 5300 9660 5340
rect 9700 5300 9760 5340
rect 9800 5300 9820 5340
rect 9640 5280 9820 5300
rect 9870 5340 9950 5360
rect 9870 5300 9890 5340
rect 9930 5300 9950 5340
rect 9870 5280 9950 5300
rect 10000 5340 10080 5360
rect 10000 5300 10020 5340
rect 10060 5300 10080 5340
rect 10000 5280 10080 5300
rect 10130 5340 10210 5360
rect 10130 5300 10150 5340
rect 10190 5300 10210 5340
rect 10130 5280 10210 5300
rect 10260 5340 10340 5360
rect 10260 5300 10280 5340
rect 10320 5300 10340 5340
rect 10260 5280 10340 5300
rect 10390 5340 10470 5360
rect 10390 5300 10410 5340
rect 10450 5300 10470 5340
rect 10390 5280 10470 5300
rect 10520 5340 10700 5360
rect 10520 5300 10540 5340
rect 10580 5300 10640 5340
rect 10680 5300 10700 5340
rect 10520 5280 10700 5300
rect 11450 5330 11560 5350
rect 7720 5220 7800 5240
rect 7720 5180 7740 5220
rect 7780 5180 7800 5220
rect 7720 5160 7800 5180
rect 8770 5220 8850 5240
rect 8770 5180 8790 5220
rect 8830 5180 8850 5220
rect 8770 5160 8850 5180
rect 9210 5220 9290 5240
rect 9210 5180 9230 5220
rect 9270 5180 9290 5220
rect 9210 5160 9290 5180
rect 10040 5120 10080 5280
rect 10260 5120 10300 5280
rect 11450 5260 11470 5330
rect 11540 5260 11560 5330
rect 11450 5240 11560 5260
rect 10750 5220 10830 5240
rect 10750 5180 10770 5220
rect 10810 5180 10830 5220
rect 10750 5160 10830 5180
rect 11450 5120 11490 5240
rect 9910 5100 9990 5120
rect 9910 5060 9930 5100
rect 9970 5060 9990 5100
rect 10040 5080 11660 5120
rect 9910 5040 9990 5060
rect 11620 5070 11660 5080
rect 11620 5050 11700 5070
rect 11620 5010 11640 5050
rect 11680 5010 11700 5050
rect 11620 4990 11700 5010
rect 11620 4980 11660 4990
rect 10040 4940 11660 4980
rect 7630 4880 7710 4900
rect 7630 4840 7650 4880
rect 7690 4840 7710 4880
rect 7630 4820 7710 4840
rect 8070 4880 8150 4900
rect 8070 4840 8090 4880
rect 8130 4840 8150 4880
rect 8070 4820 8150 4840
rect 8860 4890 8940 4910
rect 8860 4850 8880 4890
rect 8920 4850 8940 4890
rect 8860 4830 8940 4850
rect 9910 4880 9990 4900
rect 9910 4840 9930 4880
rect 9970 4840 9990 4880
rect 9910 4820 9990 4840
rect -1460 4800 -1400 4820
rect -1460 4760 -1450 4800
rect -1410 4760 -1400 4800
rect -1460 4740 -1400 4760
rect 940 4800 1000 4820
rect 940 4760 950 4800
rect 990 4760 1000 4800
rect 940 4740 1000 4760
rect 1580 4800 1640 4820
rect 1580 4760 1590 4800
rect 1630 4760 1640 4800
rect 1580 4740 1640 4760
rect 3980 4800 4040 4820
rect 3980 4760 3990 4800
rect 4030 4760 4040 4800
rect 10040 4780 10080 4940
rect 10260 4780 10300 4940
rect 10750 4880 10830 4900
rect 10750 4840 10770 4880
rect 10810 4840 10830 4880
rect 10750 4820 10830 4840
rect 11450 4840 11490 4940
rect 11450 4820 11560 4840
rect 3980 4740 4040 4760
rect 7460 4760 7540 4780
rect 7460 4720 7480 4760
rect 7520 4720 7540 4760
rect -1540 4680 -1400 4700
rect -1540 4640 -1530 4680
rect -1490 4640 -1450 4680
rect -1410 4640 -1400 4680
rect -1540 4580 -1400 4640
rect -1540 4540 -1530 4580
rect -1490 4540 -1450 4580
rect -1410 4540 -1400 4580
rect -1540 4520 -1400 4540
rect -1340 4680 -1280 4700
rect -1340 4640 -1330 4680
rect -1290 4640 -1280 4680
rect -1340 4580 -1280 4640
rect -1340 4540 -1330 4580
rect -1290 4540 -1280 4580
rect -1340 4520 -1280 4540
rect -1220 4680 -1160 4700
rect -1220 4640 -1210 4680
rect -1170 4640 -1160 4680
rect -1220 4580 -1160 4640
rect -1220 4540 -1210 4580
rect -1170 4540 -1160 4580
rect -1220 4520 -1160 4540
rect -1100 4680 -1040 4700
rect -1100 4640 -1090 4680
rect -1050 4640 -1040 4680
rect -1100 4580 -1040 4640
rect -1100 4540 -1090 4580
rect -1050 4540 -1040 4580
rect -1100 4520 -1040 4540
rect -980 4680 -920 4700
rect -980 4640 -970 4680
rect -930 4640 -920 4680
rect -980 4580 -920 4640
rect -980 4540 -970 4580
rect -930 4540 -920 4580
rect -980 4520 -920 4540
rect -860 4680 -800 4700
rect -860 4640 -850 4680
rect -810 4640 -800 4680
rect -860 4580 -800 4640
rect -860 4540 -850 4580
rect -810 4540 -800 4580
rect -860 4520 -800 4540
rect -740 4680 -680 4700
rect -740 4640 -730 4680
rect -690 4640 -680 4680
rect -740 4580 -680 4640
rect -740 4540 -730 4580
rect -690 4540 -680 4580
rect -740 4520 -680 4540
rect -620 4680 -560 4700
rect -620 4640 -610 4680
rect -570 4640 -560 4680
rect -620 4580 -560 4640
rect -620 4540 -610 4580
rect -570 4540 -560 4580
rect -620 4520 -560 4540
rect -500 4680 -440 4700
rect -500 4640 -490 4680
rect -450 4640 -440 4680
rect -500 4580 -440 4640
rect -500 4540 -490 4580
rect -450 4540 -440 4580
rect -500 4520 -440 4540
rect -380 4680 -320 4700
rect -380 4640 -370 4680
rect -330 4640 -320 4680
rect -380 4580 -320 4640
rect -380 4540 -370 4580
rect -330 4540 -320 4580
rect -380 4520 -320 4540
rect -260 4680 -200 4700
rect -260 4640 -250 4680
rect -210 4640 -200 4680
rect -260 4580 -200 4640
rect -260 4540 -250 4580
rect -210 4540 -200 4580
rect -260 4520 -200 4540
rect -140 4680 -80 4700
rect -140 4640 -130 4680
rect -90 4640 -80 4680
rect -140 4580 -80 4640
rect -140 4540 -130 4580
rect -90 4540 -80 4580
rect -140 4520 -80 4540
rect -20 4680 40 4700
rect -20 4640 -10 4680
rect 30 4640 40 4680
rect -20 4580 40 4640
rect -20 4540 -10 4580
rect 30 4540 40 4580
rect -20 4520 40 4540
rect 100 4680 160 4700
rect 100 4640 110 4680
rect 150 4640 160 4680
rect 100 4580 160 4640
rect 100 4540 110 4580
rect 150 4540 160 4580
rect 100 4520 160 4540
rect 220 4680 280 4700
rect 220 4640 230 4680
rect 270 4640 280 4680
rect 220 4580 280 4640
rect 220 4540 230 4580
rect 270 4540 280 4580
rect 220 4520 280 4540
rect 340 4680 400 4700
rect 340 4640 350 4680
rect 390 4640 400 4680
rect 340 4580 400 4640
rect 340 4540 350 4580
rect 390 4540 400 4580
rect 340 4520 400 4540
rect 460 4680 520 4700
rect 460 4640 470 4680
rect 510 4640 520 4680
rect 460 4580 520 4640
rect 460 4540 470 4580
rect 510 4540 520 4580
rect 460 4520 520 4540
rect 580 4680 640 4700
rect 580 4640 590 4680
rect 630 4640 640 4680
rect 580 4580 640 4640
rect 580 4540 590 4580
rect 630 4540 640 4580
rect 580 4520 640 4540
rect 700 4680 760 4700
rect 700 4640 710 4680
rect 750 4640 760 4680
rect 700 4580 760 4640
rect 700 4540 710 4580
rect 750 4540 760 4580
rect 700 4520 760 4540
rect 820 4680 880 4700
rect 820 4640 830 4680
rect 870 4640 880 4680
rect 820 4580 880 4640
rect 820 4540 830 4580
rect 870 4540 880 4580
rect 820 4520 880 4540
rect 940 4680 1080 4700
rect 940 4640 950 4680
rect 990 4640 1030 4680
rect 1070 4640 1080 4680
rect 940 4580 1080 4640
rect 940 4540 950 4580
rect 990 4540 1030 4580
rect 1070 4540 1080 4580
rect 940 4520 1080 4540
rect 1500 4680 1640 4700
rect 1500 4640 1510 4680
rect 1550 4640 1590 4680
rect 1630 4640 1640 4680
rect 1500 4580 1640 4640
rect 1500 4540 1510 4580
rect 1550 4540 1590 4580
rect 1630 4540 1640 4580
rect 1500 4520 1640 4540
rect 1700 4680 1760 4700
rect 1700 4640 1710 4680
rect 1750 4640 1760 4680
rect 1700 4580 1760 4640
rect 1700 4540 1710 4580
rect 1750 4540 1760 4580
rect 1700 4520 1760 4540
rect 1820 4680 1880 4700
rect 1820 4640 1830 4680
rect 1870 4640 1880 4680
rect 1820 4580 1880 4640
rect 1820 4540 1830 4580
rect 1870 4540 1880 4580
rect 1820 4520 1880 4540
rect 1940 4680 2000 4700
rect 1940 4640 1950 4680
rect 1990 4640 2000 4680
rect 1940 4580 2000 4640
rect 1940 4540 1950 4580
rect 1990 4540 2000 4580
rect 1940 4520 2000 4540
rect 2060 4680 2120 4700
rect 2060 4640 2070 4680
rect 2110 4640 2120 4680
rect 2060 4580 2120 4640
rect 2060 4540 2070 4580
rect 2110 4540 2120 4580
rect 2060 4520 2120 4540
rect 2180 4680 2240 4700
rect 2180 4640 2190 4680
rect 2230 4640 2240 4680
rect 2180 4580 2240 4640
rect 2180 4540 2190 4580
rect 2230 4540 2240 4580
rect 2180 4520 2240 4540
rect 2300 4680 2360 4700
rect 2300 4640 2310 4680
rect 2350 4640 2360 4680
rect 2300 4580 2360 4640
rect 2300 4540 2310 4580
rect 2350 4540 2360 4580
rect 2300 4520 2360 4540
rect 2420 4680 2480 4700
rect 2420 4640 2430 4680
rect 2470 4640 2480 4680
rect 2420 4580 2480 4640
rect 2420 4540 2430 4580
rect 2470 4540 2480 4580
rect 2420 4520 2480 4540
rect 2540 4680 2600 4700
rect 2540 4640 2550 4680
rect 2590 4640 2600 4680
rect 2540 4580 2600 4640
rect 2540 4540 2550 4580
rect 2590 4540 2600 4580
rect 2540 4520 2600 4540
rect 2660 4680 2720 4700
rect 2660 4640 2670 4680
rect 2710 4640 2720 4680
rect 2660 4580 2720 4640
rect 2660 4540 2670 4580
rect 2710 4540 2720 4580
rect 2660 4520 2720 4540
rect 2780 4680 2840 4700
rect 2780 4640 2790 4680
rect 2830 4640 2840 4680
rect 2780 4580 2840 4640
rect 2780 4540 2790 4580
rect 2830 4540 2840 4580
rect 2780 4520 2840 4540
rect 2900 4680 2960 4700
rect 2900 4640 2910 4680
rect 2950 4640 2960 4680
rect 2900 4580 2960 4640
rect 2900 4540 2910 4580
rect 2950 4540 2960 4580
rect 2900 4520 2960 4540
rect 3020 4680 3080 4700
rect 3020 4640 3030 4680
rect 3070 4640 3080 4680
rect 3020 4580 3080 4640
rect 3020 4540 3030 4580
rect 3070 4540 3080 4580
rect 3020 4520 3080 4540
rect 3140 4680 3200 4700
rect 3140 4640 3150 4680
rect 3190 4640 3200 4680
rect 3140 4580 3200 4640
rect 3140 4540 3150 4580
rect 3190 4540 3200 4580
rect 3140 4520 3200 4540
rect 3260 4680 3320 4700
rect 3260 4640 3270 4680
rect 3310 4640 3320 4680
rect 3260 4580 3320 4640
rect 3260 4540 3270 4580
rect 3310 4540 3320 4580
rect 3260 4520 3320 4540
rect 3380 4680 3440 4700
rect 3380 4640 3390 4680
rect 3430 4640 3440 4680
rect 3380 4580 3440 4640
rect 3380 4540 3390 4580
rect 3430 4540 3440 4580
rect 3380 4520 3440 4540
rect 3500 4680 3560 4700
rect 3500 4640 3510 4680
rect 3550 4640 3560 4680
rect 3500 4580 3560 4640
rect 3500 4540 3510 4580
rect 3550 4540 3560 4580
rect 3500 4520 3560 4540
rect 3620 4680 3680 4700
rect 3620 4640 3630 4680
rect 3670 4640 3680 4680
rect 3620 4580 3680 4640
rect 3620 4540 3630 4580
rect 3670 4540 3680 4580
rect 3620 4520 3680 4540
rect 3740 4680 3800 4700
rect 3740 4640 3750 4680
rect 3790 4640 3800 4680
rect 3740 4580 3800 4640
rect 3740 4540 3750 4580
rect 3790 4540 3800 4580
rect 3740 4520 3800 4540
rect 3860 4680 3920 4700
rect 3860 4640 3870 4680
rect 3910 4640 3920 4680
rect 3860 4580 3920 4640
rect 3860 4540 3870 4580
rect 3910 4540 3920 4580
rect 3860 4520 3920 4540
rect 3980 4680 4120 4700
rect 3980 4640 3990 4680
rect 4030 4640 4070 4680
rect 4110 4640 4120 4680
rect 3980 4580 4120 4640
rect 7460 4660 7540 4720
rect 7460 4620 7480 4660
rect 7520 4620 7540 4660
rect 7460 4600 7540 4620
rect 7590 4760 7670 4780
rect 7590 4720 7610 4760
rect 7650 4720 7670 4760
rect 7590 4660 7670 4720
rect 7590 4620 7610 4660
rect 7650 4620 7670 4660
rect 7590 4600 7670 4620
rect 7720 4760 7800 4780
rect 7720 4720 7740 4760
rect 7780 4720 7800 4760
rect 7720 4660 7800 4720
rect 7720 4620 7740 4660
rect 7780 4620 7800 4660
rect 7720 4600 7800 4620
rect 7850 4760 7930 4780
rect 7850 4720 7870 4760
rect 7910 4720 7930 4760
rect 7850 4660 7930 4720
rect 7850 4620 7870 4660
rect 7910 4620 7930 4660
rect 7850 4600 7930 4620
rect 7980 4760 8060 4780
rect 7980 4720 8000 4760
rect 8040 4720 8060 4760
rect 7980 4660 8060 4720
rect 7980 4620 8000 4660
rect 8040 4620 8060 4660
rect 7980 4600 8060 4620
rect 8110 4760 8200 4780
rect 8110 4720 8130 4760
rect 8170 4720 8200 4760
rect 8110 4660 8200 4720
rect 8110 4620 8130 4660
rect 8170 4620 8200 4660
rect 8110 4600 8200 4620
rect 8240 4760 8320 4780
rect 8240 4720 8260 4760
rect 8300 4720 8320 4760
rect 8240 4660 8320 4720
rect 8240 4620 8260 4660
rect 8300 4620 8320 4660
rect 8240 4600 8320 4620
rect 8500 4760 8680 4780
rect 8500 4720 8520 4760
rect 8560 4720 8620 4760
rect 8660 4720 8680 4760
rect 8500 4660 8680 4720
rect 8500 4620 8520 4660
rect 8560 4620 8620 4660
rect 8660 4620 8680 4660
rect 8500 4600 8680 4620
rect 8730 4760 8810 4780
rect 8730 4720 8750 4760
rect 8790 4720 8810 4760
rect 8730 4660 8810 4720
rect 8730 4620 8750 4660
rect 8790 4620 8810 4660
rect 8730 4600 8810 4620
rect 8860 4760 8940 4780
rect 8860 4720 8880 4760
rect 8920 4720 8940 4760
rect 8860 4660 8940 4720
rect 8860 4620 8880 4660
rect 8920 4620 8940 4660
rect 8860 4600 8940 4620
rect 8990 4760 9070 4780
rect 8990 4720 9010 4760
rect 9050 4720 9070 4760
rect 8990 4660 9070 4720
rect 8990 4620 9010 4660
rect 9050 4620 9070 4660
rect 8990 4600 9070 4620
rect 9120 4760 9200 4780
rect 9120 4720 9140 4760
rect 9180 4720 9200 4760
rect 9120 4660 9200 4720
rect 9120 4620 9140 4660
rect 9180 4620 9200 4660
rect 9120 4600 9200 4620
rect 9250 4760 9330 4780
rect 9250 4720 9270 4760
rect 9310 4720 9330 4760
rect 9250 4660 9330 4720
rect 9250 4620 9270 4660
rect 9310 4620 9330 4660
rect 9250 4600 9330 4620
rect 9380 4760 9560 4780
rect 9380 4720 9400 4760
rect 9440 4720 9500 4760
rect 9540 4720 9560 4760
rect 9380 4660 9560 4720
rect 9380 4620 9400 4660
rect 9440 4620 9500 4660
rect 9540 4620 9560 4660
rect 9380 4600 9560 4620
rect 9640 4760 9820 4780
rect 9640 4720 9660 4760
rect 9700 4720 9760 4760
rect 9800 4720 9820 4760
rect 9640 4660 9820 4720
rect 9640 4620 9660 4660
rect 9700 4620 9760 4660
rect 9800 4620 9820 4660
rect 9640 4600 9820 4620
rect 9870 4760 9950 4780
rect 9870 4720 9890 4760
rect 9930 4720 9950 4760
rect 9870 4660 9950 4720
rect 9870 4620 9890 4660
rect 9930 4620 9950 4660
rect 9870 4600 9950 4620
rect 10000 4760 10080 4780
rect 10000 4720 10020 4760
rect 10060 4720 10080 4760
rect 10000 4660 10080 4720
rect 10000 4620 10020 4660
rect 10060 4620 10080 4660
rect 10000 4600 10080 4620
rect 10130 4760 10210 4780
rect 10130 4720 10150 4760
rect 10190 4720 10210 4760
rect 10130 4660 10210 4720
rect 10130 4620 10150 4660
rect 10190 4620 10210 4660
rect 10130 4600 10210 4620
rect 10260 4760 10340 4780
rect 10260 4720 10280 4760
rect 10320 4720 10340 4760
rect 10260 4660 10340 4720
rect 10260 4620 10280 4660
rect 10320 4620 10340 4660
rect 10260 4600 10340 4620
rect 10390 4760 10470 4780
rect 10390 4720 10410 4760
rect 10450 4720 10470 4760
rect 10390 4660 10470 4720
rect 10390 4620 10410 4660
rect 10450 4620 10470 4660
rect 10390 4600 10470 4620
rect 10520 4760 10700 4780
rect 10520 4720 10540 4760
rect 10580 4720 10640 4760
rect 10680 4720 10700 4760
rect 11450 4750 11470 4820
rect 11540 4750 11560 4820
rect 11450 4730 11560 4750
rect 10520 4660 10700 4720
rect 10520 4620 10540 4660
rect 10580 4620 10640 4660
rect 10680 4620 10700 4660
rect 10520 4600 10700 4620
rect 3980 4540 3990 4580
rect 4030 4540 4070 4580
rect 4110 4540 4120 4580
rect 3980 4520 4120 4540
rect 7480 4560 7520 4600
rect 7610 4560 7650 4600
rect 7870 4560 7910 4600
rect 8130 4560 8170 4600
rect 8260 4560 8300 4600
rect 7480 4540 8300 4560
rect 7480 4520 7540 4540
rect 7520 4500 7540 4520
rect 7580 4520 8200 4540
rect 7580 4500 7600 4520
rect 7520 4480 7600 4500
rect 7930 4500 8010 4520
rect -1280 4450 -1220 4470
rect -1280 4410 -1270 4450
rect -1230 4410 -1220 4450
rect -1280 4390 -1220 4410
rect -1110 4460 -1030 4480
rect -1110 4420 -1090 4460
rect -1050 4420 -1030 4460
rect -1110 4400 -1030 4420
rect -620 4460 -560 4480
rect -620 4420 -610 4460
rect -570 4420 -560 4460
rect -620 4400 -560 4420
rect -390 4460 -310 4480
rect -390 4420 -370 4460
rect -330 4420 -310 4460
rect -390 4400 -310 4420
rect 100 4460 160 4480
rect 100 4420 110 4460
rect 150 4420 160 4460
rect 100 4400 160 4420
rect 330 4460 410 4480
rect 330 4420 350 4460
rect 390 4420 410 4460
rect 330 4400 410 4420
rect 760 4460 820 4480
rect 760 4420 770 4460
rect 810 4420 820 4460
rect 760 4400 820 4420
rect 1760 4460 1820 4480
rect 1760 4420 1770 4460
rect 1810 4420 1820 4460
rect 1760 4400 1820 4420
rect 2170 4460 2250 4480
rect 2170 4420 2190 4460
rect 2230 4420 2250 4460
rect 2170 4400 2250 4420
rect 2420 4460 2480 4480
rect 2420 4420 2430 4460
rect 2470 4420 2480 4460
rect 2420 4400 2480 4420
rect 2890 4460 2970 4480
rect 2890 4420 2910 4460
rect 2950 4420 2970 4460
rect 2890 4400 2970 4420
rect 3140 4460 3200 4480
rect 3140 4420 3150 4460
rect 3190 4420 3200 4460
rect 3140 4400 3200 4420
rect 3610 4460 3690 4480
rect 3610 4420 3630 4460
rect 3670 4420 3690 4460
rect 3610 4400 3690 4420
rect 3800 4450 3860 4470
rect 3800 4410 3810 4450
rect 3850 4410 3860 4450
rect 7930 4460 7950 4500
rect 7990 4460 8010 4500
rect 8180 4500 8200 4520
rect 8240 4520 8300 4540
rect 8620 4560 8660 4600
rect 8750 4560 8790 4600
rect 9010 4560 9050 4600
rect 9270 4560 9310 4600
rect 9400 4560 9440 4600
rect 8620 4540 9440 4560
rect 8620 4520 8680 4540
rect 8240 4500 8260 4520
rect 8180 4480 8260 4500
rect 8660 4500 8680 4520
rect 8720 4520 9340 4540
rect 8720 4500 8740 4520
rect 8660 4480 8740 4500
rect 7930 4440 8010 4460
rect 3800 4390 3860 4410
rect 9010 4410 9050 4520
rect 9320 4500 9340 4520
rect 9380 4520 9440 4540
rect 9760 4560 9800 4600
rect 9890 4560 9930 4600
rect 10150 4560 10190 4600
rect 10410 4560 10450 4600
rect 10540 4560 10580 4600
rect 9760 4540 10580 4560
rect 9760 4520 9820 4540
rect 9380 4500 9400 4520
rect 9320 4480 9400 4500
rect 9800 4500 9820 4520
rect 9860 4520 10480 4540
rect 9860 4500 9880 4520
rect 9800 4480 9880 4500
rect 10150 4410 10190 4520
rect 10460 4500 10480 4520
rect 10520 4520 10580 4540
rect 10520 4500 10540 4520
rect 10460 4480 10540 4500
rect 9010 4390 9090 4410
rect 9010 4350 9030 4390
rect 9070 4350 9090 4390
rect 9010 4330 9090 4350
rect 10130 4390 10210 4410
rect 10130 4350 10150 4390
rect 10190 4350 10210 4390
rect 10130 4330 10210 4350
rect 11043 4347 11139 4381
rect 11399 4347 11495 4381
rect 11043 4285 11077 4347
rect 7530 4230 7610 4250
rect 7530 4190 7550 4230
rect 7590 4190 7610 4230
rect 7530 4130 7610 4190
rect 9530 4230 9610 4250
rect 9530 4190 9550 4230
rect 9590 4190 9610 4230
rect 9530 4170 9610 4190
rect 7430 4110 7610 4130
rect 7430 4070 7450 4110
rect 7490 4070 7550 4110
rect 7590 4070 7610 4110
rect 7430 4010 7610 4070
rect 7430 3970 7450 4010
rect 7490 3970 7550 4010
rect 7590 3970 7610 4010
rect 7430 3910 7610 3970
rect 7430 3870 7450 3910
rect 7490 3870 7550 3910
rect 7590 3870 7610 3910
rect -458 3852 -400 3870
rect -458 3818 -446 3852
rect -412 3818 -400 3852
rect -458 3800 -400 3818
rect -300 3852 -242 3870
rect -300 3818 -288 3852
rect -254 3818 -242 3852
rect -300 3800 -242 3818
rect 24 3852 82 3870
rect 24 3818 36 3852
rect 70 3818 82 3852
rect 24 3800 82 3818
rect 178 3852 236 3870
rect 178 3818 190 3852
rect 224 3818 236 3852
rect 178 3800 236 3818
rect 502 3852 560 3870
rect 502 3818 514 3852
rect 548 3818 560 3852
rect 2020 3852 2078 3870
rect 502 3800 560 3818
rect 810 3810 890 3830
rect 810 3770 830 3810
rect 870 3770 890 3810
rect -620 3740 -560 3760
rect -620 3700 -610 3740
rect -570 3700 -560 3740
rect -620 3680 -560 3700
rect -500 3740 -440 3760
rect -500 3700 -490 3740
rect -450 3700 -440 3740
rect -500 3680 -440 3700
rect -380 3740 -320 3760
rect -380 3700 -370 3740
rect -330 3700 -320 3740
rect -380 3680 -320 3700
rect -260 3740 -200 3760
rect -260 3700 -250 3740
rect -210 3700 -200 3740
rect -260 3680 -200 3700
rect -140 3740 -80 3760
rect -140 3700 -130 3740
rect -90 3700 -80 3740
rect -140 3680 -80 3700
rect -20 3740 40 3760
rect -20 3700 -10 3740
rect 30 3700 40 3740
rect -20 3680 40 3700
rect 100 3740 160 3760
rect 100 3700 110 3740
rect 150 3700 160 3740
rect 100 3680 160 3700
rect 220 3740 280 3760
rect 220 3700 230 3740
rect 270 3700 280 3740
rect 220 3680 280 3700
rect 340 3740 400 3760
rect 340 3700 350 3740
rect 390 3700 400 3740
rect 340 3680 400 3700
rect 460 3740 520 3760
rect 460 3700 470 3740
rect 510 3700 520 3740
rect 460 3680 520 3700
rect 580 3740 640 3760
rect 580 3700 590 3740
rect 630 3700 640 3740
rect 580 3680 640 3700
rect 810 3730 890 3770
rect 810 3690 830 3730
rect 870 3690 890 3730
rect 810 3650 890 3690
rect -559 3622 -501 3640
rect -559 3588 -547 3622
rect -513 3588 -501 3622
rect -559 3570 -501 3588
rect -199 3622 -141 3640
rect -199 3588 -187 3622
rect -153 3588 -141 3622
rect -199 3570 -141 3588
rect -79 3622 -21 3640
rect -79 3588 -67 3622
rect -33 3588 -21 3622
rect -79 3570 -21 3588
rect 281 3622 339 3640
rect 281 3588 293 3622
rect 327 3588 339 3622
rect 281 3570 339 3588
rect 401 3622 459 3640
rect 401 3588 413 3622
rect 447 3588 459 3622
rect 810 3610 830 3650
rect 870 3610 890 3650
rect 810 3590 890 3610
rect 1690 3810 1770 3830
rect 1690 3770 1710 3810
rect 1750 3770 1770 3810
rect 2020 3818 2032 3852
rect 2066 3818 2078 3852
rect 2020 3800 2078 3818
rect 2344 3852 2402 3870
rect 2344 3818 2356 3852
rect 2390 3818 2402 3852
rect 2344 3800 2402 3818
rect 2498 3852 2556 3870
rect 2498 3818 2510 3852
rect 2544 3818 2556 3852
rect 2498 3800 2556 3818
rect 2822 3852 2880 3870
rect 2822 3818 2834 3852
rect 2868 3818 2880 3852
rect 2822 3800 2880 3818
rect 2980 3852 3038 3870
rect 2980 3818 2992 3852
rect 3026 3818 3038 3852
rect 2980 3800 3038 3818
rect 7430 3810 7610 3870
rect 1690 3730 1770 3770
rect 7430 3770 7450 3810
rect 7490 3770 7550 3810
rect 7590 3770 7610 3810
rect 1690 3690 1710 3730
rect 1750 3690 1770 3730
rect 1690 3650 1770 3690
rect 1940 3740 2000 3760
rect 1940 3700 1950 3740
rect 1990 3700 2000 3740
rect 1940 3680 2000 3700
rect 2060 3740 2120 3760
rect 2060 3700 2070 3740
rect 2110 3700 2120 3740
rect 2060 3680 2120 3700
rect 2180 3740 2240 3760
rect 2180 3700 2190 3740
rect 2230 3700 2240 3740
rect 2180 3680 2240 3700
rect 2300 3740 2360 3760
rect 2300 3700 2310 3740
rect 2350 3700 2360 3740
rect 2300 3680 2360 3700
rect 2420 3740 2480 3760
rect 2420 3700 2430 3740
rect 2470 3700 2480 3740
rect 2420 3680 2480 3700
rect 2540 3740 2600 3760
rect 2540 3700 2550 3740
rect 2590 3700 2600 3740
rect 2540 3680 2600 3700
rect 2660 3740 2720 3760
rect 2660 3700 2670 3740
rect 2710 3700 2720 3740
rect 2660 3680 2720 3700
rect 2780 3740 2840 3760
rect 2780 3700 2790 3740
rect 2830 3700 2840 3740
rect 2780 3680 2840 3700
rect 2900 3740 2960 3760
rect 2900 3700 2910 3740
rect 2950 3700 2960 3740
rect 2900 3680 2960 3700
rect 3020 3740 3080 3760
rect 3020 3700 3030 3740
rect 3070 3700 3080 3740
rect 3020 3680 3080 3700
rect 3140 3740 3200 3760
rect 3140 3700 3150 3740
rect 3190 3700 3200 3740
rect 3140 3680 3200 3700
rect 7430 3710 7610 3770
rect 7430 3670 7450 3710
rect 7490 3670 7550 3710
rect 7590 3670 7610 3710
rect 7430 3650 7610 3670
rect 7730 4110 7810 4130
rect 7730 4070 7750 4110
rect 7790 4070 7810 4110
rect 7730 4010 7810 4070
rect 7730 3970 7750 4010
rect 7790 3970 7810 4010
rect 7730 3910 7810 3970
rect 7730 3870 7750 3910
rect 7790 3870 7810 3910
rect 7730 3810 7810 3870
rect 7730 3770 7750 3810
rect 7790 3770 7810 3810
rect 7730 3710 7810 3770
rect 7730 3670 7750 3710
rect 7790 3670 7810 3710
rect 7730 3650 7810 3670
rect 7930 4110 8010 4130
rect 7930 4070 7950 4110
rect 7990 4070 8010 4110
rect 7930 4010 8010 4070
rect 7930 3970 7950 4010
rect 7990 3970 8010 4010
rect 7930 3910 8010 3970
rect 7930 3870 7950 3910
rect 7990 3870 8010 3910
rect 7930 3810 8010 3870
rect 7930 3770 7950 3810
rect 7990 3770 8010 3810
rect 7930 3710 8010 3770
rect 7930 3670 7950 3710
rect 7990 3670 8010 3710
rect 7930 3650 8010 3670
rect 8130 4110 8210 4130
rect 8130 4070 8150 4110
rect 8190 4070 8210 4110
rect 8130 4010 8210 4070
rect 8130 3970 8150 4010
rect 8190 3970 8210 4010
rect 8130 3910 8210 3970
rect 8130 3870 8150 3910
rect 8190 3870 8210 3910
rect 8130 3810 8210 3870
rect 8130 3770 8150 3810
rect 8190 3770 8210 3810
rect 8130 3710 8210 3770
rect 8130 3670 8150 3710
rect 8190 3670 8210 3710
rect 8130 3650 8210 3670
rect 8330 4110 8410 4130
rect 8330 4070 8350 4110
rect 8390 4070 8410 4110
rect 8330 4010 8410 4070
rect 8330 3970 8350 4010
rect 8390 3970 8410 4010
rect 8330 3910 8410 3970
rect 8330 3870 8350 3910
rect 8390 3870 8410 3910
rect 8330 3810 8410 3870
rect 8330 3770 8350 3810
rect 8390 3770 8410 3810
rect 8330 3710 8410 3770
rect 8330 3670 8350 3710
rect 8390 3670 8410 3710
rect 8330 3650 8410 3670
rect 8530 4110 8610 4130
rect 8530 4070 8550 4110
rect 8590 4070 8610 4110
rect 8530 4010 8610 4070
rect 8530 3970 8550 4010
rect 8590 3970 8610 4010
rect 8530 3910 8610 3970
rect 8530 3870 8550 3910
rect 8590 3870 8610 3910
rect 8530 3810 8610 3870
rect 8530 3770 8550 3810
rect 8590 3770 8610 3810
rect 8530 3710 8610 3770
rect 8530 3670 8550 3710
rect 8590 3670 8610 3710
rect 8530 3650 8610 3670
rect 8730 4110 8810 4130
rect 8730 4070 8750 4110
rect 8790 4070 8810 4110
rect 8730 4010 8810 4070
rect 8730 3970 8750 4010
rect 8790 3970 8810 4010
rect 8730 3910 8810 3970
rect 8730 3870 8750 3910
rect 8790 3870 8810 3910
rect 8730 3810 8810 3870
rect 8730 3770 8750 3810
rect 8790 3770 8810 3810
rect 8730 3710 8810 3770
rect 8730 3670 8750 3710
rect 8790 3670 8810 3710
rect 8730 3650 8810 3670
rect 8930 4110 9010 4130
rect 8930 4070 8950 4110
rect 8990 4070 9010 4110
rect 8930 4010 9010 4070
rect 8930 3970 8950 4010
rect 8990 3970 9010 4010
rect 8930 3910 9010 3970
rect 8930 3870 8950 3910
rect 8990 3870 9010 3910
rect 8930 3810 9010 3870
rect 8930 3770 8950 3810
rect 8990 3770 9010 3810
rect 8930 3710 9010 3770
rect 8930 3670 8950 3710
rect 8990 3670 9010 3710
rect 8930 3650 9010 3670
rect 9130 4110 9210 4130
rect 9130 4070 9150 4110
rect 9190 4070 9210 4110
rect 9130 4010 9210 4070
rect 9130 3970 9150 4010
rect 9190 3970 9210 4010
rect 9130 3910 9210 3970
rect 9130 3870 9150 3910
rect 9190 3870 9210 3910
rect 9130 3810 9210 3870
rect 9130 3770 9150 3810
rect 9190 3770 9210 3810
rect 9130 3710 9210 3770
rect 9130 3670 9150 3710
rect 9190 3670 9210 3710
rect 9130 3650 9210 3670
rect 9330 4110 9410 4130
rect 9330 4070 9350 4110
rect 9390 4070 9410 4110
rect 9330 4010 9410 4070
rect 9330 3970 9350 4010
rect 9390 3970 9410 4010
rect 9330 3910 9410 3970
rect 9330 3870 9350 3910
rect 9390 3870 9410 3910
rect 9330 3810 9410 3870
rect 9330 3770 9350 3810
rect 9390 3770 9410 3810
rect 9330 3710 9410 3770
rect 9330 3670 9350 3710
rect 9390 3670 9410 3710
rect 9330 3650 9410 3670
rect 9530 4110 9710 4130
rect 9530 4070 9550 4110
rect 9590 4070 9650 4110
rect 9690 4070 9710 4110
rect 9530 4010 9710 4070
rect 9530 3970 9550 4010
rect 9590 3970 9650 4010
rect 9690 3970 9710 4010
rect 9530 3910 9710 3970
rect 9530 3870 9550 3910
rect 9590 3870 9650 3910
rect 9690 3870 9710 3910
rect 9530 3810 9710 3870
rect 9530 3770 9550 3810
rect 9590 3770 9650 3810
rect 9690 3770 9710 3810
rect 9530 3710 9710 3770
rect 9530 3670 9550 3710
rect 9590 3670 9650 3710
rect 9690 3670 9710 3710
rect 9530 3650 9710 3670
rect 1690 3610 1710 3650
rect 1750 3610 1770 3650
rect 1690 3590 1770 3610
rect 2121 3622 2179 3640
rect 401 3570 459 3588
rect 2121 3588 2133 3622
rect 2167 3588 2179 3622
rect 2121 3570 2179 3588
rect 2241 3622 2299 3640
rect 2241 3588 2253 3622
rect 2287 3588 2299 3622
rect 2241 3570 2299 3588
rect 2601 3622 2659 3640
rect 2601 3588 2613 3622
rect 2647 3588 2659 3622
rect 2601 3570 2659 3588
rect 2721 3622 2779 3640
rect 2721 3588 2733 3622
rect 2767 3588 2779 3622
rect 2721 3570 2779 3588
rect 3081 3622 3139 3640
rect 3081 3588 3093 3622
rect 3127 3588 3139 3622
rect 3081 3570 3139 3588
rect 8330 3590 8410 3610
rect 8330 3550 8350 3590
rect 8390 3550 8410 3590
rect 8330 3530 8410 3550
rect 8730 3590 8810 3610
rect 8730 3550 8750 3590
rect 8790 3550 8810 3590
rect 8730 3530 8810 3550
rect -1070 3250 -990 3270
rect -1250 3210 -1170 3230
rect -1250 3170 -1230 3210
rect -1190 3170 -1170 3210
rect -1070 3210 -1050 3250
rect -1010 3210 -990 3250
rect -1070 3190 -990 3210
rect -830 3250 -750 3270
rect -830 3210 -810 3250
rect -770 3210 -750 3250
rect -830 3190 -750 3210
rect -590 3250 -510 3270
rect -590 3210 -570 3250
rect -530 3210 -510 3250
rect -590 3190 -510 3210
rect -350 3250 -270 3270
rect -350 3210 -330 3250
rect -290 3210 -270 3250
rect -350 3190 -270 3210
rect 290 3250 370 3270
rect 290 3210 310 3250
rect 350 3210 370 3250
rect 290 3190 370 3210
rect 530 3250 610 3270
rect 530 3210 550 3250
rect 590 3210 610 3250
rect 530 3190 610 3210
rect 770 3250 850 3270
rect 770 3210 790 3250
rect 830 3210 850 3250
rect 1730 3250 1810 3270
rect 770 3190 850 3210
rect 1080 3220 1140 3240
rect -1250 3150 -1170 3170
rect 1080 3180 1090 3220
rect 1130 3180 1140 3220
rect -1240 3130 -1180 3150
rect -1240 3090 -1230 3130
rect -1190 3090 -1180 3130
rect -1240 3030 -1180 3090
rect -1240 2990 -1230 3030
rect -1190 2990 -1180 3030
rect -1240 2930 -1180 2990
rect -1240 2890 -1230 2930
rect -1190 2890 -1180 2930
rect -1240 2830 -1180 2890
rect -1240 2790 -1230 2830
rect -1190 2790 -1180 2830
rect -1240 2730 -1180 2790
rect -1240 2690 -1230 2730
rect -1190 2690 -1180 2730
rect -1240 2670 -1180 2690
rect -160 3130 60 3150
rect -160 3090 -150 3130
rect -110 3090 -70 3130
rect -30 3090 10 3130
rect 50 3090 60 3130
rect -160 3030 60 3090
rect -160 2990 -150 3030
rect -110 2990 -70 3030
rect -30 2990 10 3030
rect 50 2990 60 3030
rect -160 2930 60 2990
rect -160 2890 -150 2930
rect -110 2890 -70 2930
rect -30 2890 10 2930
rect 50 2890 60 2930
rect -160 2830 60 2890
rect -160 2790 -150 2830
rect -110 2790 -70 2830
rect -30 2790 10 2830
rect 50 2790 60 2830
rect -160 2730 60 2790
rect -160 2690 -150 2730
rect -110 2690 -70 2730
rect -30 2690 10 2730
rect 50 2690 60 2730
rect -160 2670 60 2690
rect 1080 3130 1140 3180
rect 1080 3090 1090 3130
rect 1130 3090 1140 3130
rect 1080 3030 1140 3090
rect 1080 2990 1090 3030
rect 1130 2990 1140 3030
rect 1080 2930 1140 2990
rect 1080 2890 1090 2930
rect 1130 2890 1140 2930
rect 1080 2830 1140 2890
rect 1080 2790 1090 2830
rect 1130 2790 1140 2830
rect 1080 2730 1140 2790
rect 1080 2690 1090 2730
rect 1130 2690 1140 2730
rect 1080 2670 1140 2690
rect 1440 3220 1500 3240
rect 1440 3180 1450 3220
rect 1490 3180 1500 3220
rect 1730 3210 1750 3250
rect 1790 3210 1810 3250
rect 1730 3190 1810 3210
rect 1970 3250 2050 3270
rect 1970 3210 1990 3250
rect 2030 3210 2050 3250
rect 1970 3190 2050 3210
rect 2210 3250 2290 3270
rect 2210 3210 2230 3250
rect 2270 3210 2290 3250
rect 2210 3190 2290 3210
rect 2850 3250 2930 3270
rect 2850 3210 2870 3250
rect 2910 3210 2930 3250
rect 2850 3190 2930 3210
rect 3090 3250 3170 3270
rect 3090 3210 3110 3250
rect 3150 3210 3170 3250
rect 3090 3190 3170 3210
rect 3330 3250 3410 3270
rect 3330 3210 3350 3250
rect 3390 3210 3410 3250
rect 3330 3190 3410 3210
rect 3570 3250 3650 3270
rect 3570 3210 3590 3250
rect 3630 3210 3650 3250
rect 3570 3190 3650 3210
rect 11020 3200 11043 3220
rect 11461 4285 11495 4347
rect 11077 3200 11100 3220
rect 1440 3130 1500 3180
rect 11020 3160 11040 3200
rect 11080 3160 11100 3200
rect 1440 3090 1450 3130
rect 1490 3090 1500 3130
rect 1440 3030 1500 3090
rect 1440 2990 1450 3030
rect 1490 2990 1500 3030
rect 1440 2930 1500 2990
rect 1440 2890 1450 2930
rect 1490 2890 1500 2930
rect 1440 2830 1500 2890
rect 1440 2790 1450 2830
rect 1490 2790 1500 2830
rect 1440 2730 1500 2790
rect 1440 2690 1450 2730
rect 1490 2690 1500 2730
rect 1440 2670 1500 2690
rect 2520 3130 2740 3150
rect 2520 3090 2530 3130
rect 2570 3090 2610 3130
rect 2650 3090 2690 3130
rect 2730 3090 2740 3130
rect 2520 3030 2740 3090
rect 2520 2990 2530 3030
rect 2570 2990 2610 3030
rect 2650 2990 2690 3030
rect 2730 2990 2740 3030
rect 2520 2930 2740 2990
rect 2520 2890 2530 2930
rect 2570 2890 2610 2930
rect 2650 2890 2690 2930
rect 2730 2890 2740 2930
rect 2520 2830 2740 2890
rect 2520 2790 2530 2830
rect 2570 2790 2610 2830
rect 2650 2790 2690 2830
rect 2730 2790 2740 2830
rect 2520 2730 2740 2790
rect 2520 2690 2530 2730
rect 2570 2690 2610 2730
rect 2650 2690 2690 2730
rect 2730 2690 2740 2730
rect 2520 2670 2740 2690
rect 3760 3130 3820 3150
rect 11020 3140 11043 3160
rect 3760 3090 3770 3130
rect 3810 3090 3820 3130
rect 3760 3030 3820 3090
rect 11077 3140 11100 3160
rect 11043 3077 11077 3139
rect 11461 3077 11495 3139
rect 11043 3043 11139 3077
rect 11399 3043 11495 3077
rect 3760 2990 3770 3030
rect 3810 2990 3820 3030
rect 3760 2930 3820 2990
rect 3760 2890 3770 2930
rect 3810 2890 3820 2930
rect 3760 2830 3820 2890
rect 3760 2790 3770 2830
rect 3810 2790 3820 2830
rect 11220 2880 11320 2900
rect 11220 2820 11240 2880
rect 11300 2820 11320 2880
rect 11220 2800 11320 2820
rect 3760 2730 3820 2790
rect 3760 2690 3770 2730
rect 3810 2690 3820 2730
rect 3760 2670 3820 2690
rect -70 2630 -30 2670
rect 2610 2630 2650 2670
rect -90 2610 -10 2630
rect -90 2570 -70 2610
rect -30 2570 -10 2610
rect -90 2550 -10 2570
rect 2590 2610 2670 2630
rect 2590 2570 2610 2610
rect 2650 2570 2670 2610
rect 2590 2550 2670 2570
rect -830 2340 -750 2360
rect -830 2300 -810 2340
rect -770 2300 -750 2340
rect -830 2280 -750 2300
rect -670 2340 -590 2360
rect -670 2300 -650 2340
rect -610 2300 -590 2340
rect -670 2280 -590 2300
rect -510 2340 -430 2360
rect -510 2300 -490 2340
rect -450 2300 -430 2340
rect -510 2280 -430 2300
rect -350 2340 -270 2360
rect -350 2300 -330 2340
rect -290 2300 -270 2340
rect -350 2280 -270 2300
rect -190 2340 -110 2360
rect -190 2300 -170 2340
rect -130 2300 -110 2340
rect -190 2280 -110 2300
rect -30 2340 50 2360
rect -30 2300 -10 2340
rect 30 2300 50 2340
rect -30 2280 50 2300
rect 130 2340 210 2360
rect 130 2300 150 2340
rect 190 2300 210 2340
rect 130 2280 210 2300
rect 290 2340 370 2360
rect 290 2300 310 2340
rect 350 2300 370 2340
rect 290 2280 370 2300
rect 450 2340 530 2360
rect 450 2300 470 2340
rect 510 2300 530 2340
rect 450 2280 530 2300
rect 610 2340 690 2360
rect 610 2300 630 2340
rect 670 2300 690 2340
rect 610 2280 690 2300
rect 770 2340 850 2360
rect 770 2300 790 2340
rect 830 2300 850 2340
rect 770 2280 850 2300
rect 930 2340 1010 2360
rect 930 2300 950 2340
rect 990 2300 1010 2340
rect 930 2280 1010 2300
rect 1090 2340 1170 2360
rect 1090 2300 1110 2340
rect 1150 2300 1170 2340
rect 1090 2280 1170 2300
rect 1250 2340 1330 2360
rect 1250 2300 1270 2340
rect 1310 2300 1330 2340
rect 1250 2280 1330 2300
rect 1410 2340 1490 2360
rect 1410 2300 1430 2340
rect 1470 2300 1490 2340
rect 1410 2280 1490 2300
rect 1570 2340 1650 2360
rect 1570 2300 1590 2340
rect 1630 2300 1650 2340
rect 1570 2280 1650 2300
rect 1730 2340 1810 2360
rect 1730 2300 1750 2340
rect 1790 2300 1810 2340
rect 1730 2280 1810 2300
rect 1890 2340 1970 2360
rect 1890 2300 1910 2340
rect 1950 2300 1970 2340
rect 1890 2280 1970 2300
rect 2050 2340 2130 2360
rect 2050 2300 2070 2340
rect 2110 2300 2130 2340
rect 2050 2280 2130 2300
rect 2210 2340 2290 2360
rect 2210 2300 2230 2340
rect 2270 2300 2290 2340
rect 2210 2280 2290 2300
rect 2370 2340 2450 2360
rect 2370 2300 2390 2340
rect 2430 2300 2450 2340
rect 2370 2280 2450 2300
rect 2530 2340 2610 2360
rect 2530 2300 2550 2340
rect 2590 2300 2610 2340
rect 2530 2280 2610 2300
rect 2690 2340 2770 2360
rect 2690 2300 2710 2340
rect 2750 2300 2770 2340
rect 2690 2280 2770 2300
rect 2850 2340 2930 2360
rect 2850 2300 2870 2340
rect 2910 2300 2930 2340
rect 2850 2280 2930 2300
rect 3010 2340 3090 2360
rect 3010 2300 3030 2340
rect 3070 2300 3090 2340
rect 3010 2280 3090 2300
rect 3170 2340 3250 2360
rect 3170 2300 3190 2340
rect 3230 2300 3250 2340
rect 3170 2280 3250 2300
rect -810 2240 -770 2280
rect 1270 2240 1310 2280
rect -820 2220 -760 2240
rect -820 2190 -810 2220
rect -910 2180 -810 2190
rect -770 2180 -760 2220
rect -910 2170 -760 2180
rect -910 2130 -890 2170
rect -850 2130 -760 2170
rect -910 2120 -760 2130
rect -910 2110 -810 2120
rect -820 2080 -810 2110
rect -770 2080 -760 2120
rect -820 2060 -760 2080
rect 1260 2220 1320 2240
rect 1260 2180 1270 2220
rect 1310 2180 1320 2220
rect 1260 2120 1320 2180
rect 1260 2080 1270 2120
rect 1310 2080 1320 2120
rect 1260 2060 1320 2080
rect 3340 2230 3480 2240
rect 3340 2220 3560 2230
rect 3340 2180 3350 2220
rect 3390 2180 3430 2220
rect 3470 2210 3560 2220
rect 3470 2180 3500 2210
rect 3340 2170 3500 2180
rect 3540 2170 3560 2210
rect 3340 2130 3560 2170
rect 3340 2120 3500 2130
rect 3340 2080 3350 2120
rect 3390 2080 3430 2120
rect 3470 2090 3500 2120
rect 3540 2090 3560 2130
rect 3470 2080 3560 2090
rect 3340 2070 3560 2080
rect 3340 2060 3480 2070
rect 552 1780 642 1790
rect 552 1730 572 1780
rect 622 1730 642 1780
rect 552 1720 642 1730
rect 1950 1780 2040 1790
rect 1950 1730 1970 1780
rect 2020 1730 2040 1780
rect 1950 1720 2040 1730
rect -720 1519 3300 1560
rect -720 1496 -580 1519
rect -720 1462 -681 1496
rect -647 1485 -580 1496
rect -546 1485 -490 1519
rect -456 1485 -400 1519
rect -366 1485 -310 1519
rect -276 1485 -220 1519
rect -186 1485 -130 1519
rect -96 1485 -40 1519
rect -6 1485 50 1519
rect 84 1485 140 1519
rect 174 1485 230 1519
rect 264 1485 320 1519
rect 354 1485 410 1519
rect 444 1496 780 1519
rect 444 1485 506 1496
rect -647 1462 506 1485
rect 540 1462 679 1496
rect 713 1485 780 1496
rect 814 1485 870 1519
rect 904 1485 960 1519
rect 994 1485 1050 1519
rect 1084 1485 1140 1519
rect 1174 1485 1230 1519
rect 1264 1485 1320 1519
rect 1354 1485 1410 1519
rect 1444 1485 1500 1519
rect 1534 1485 1590 1519
rect 1624 1485 1680 1519
rect 1714 1485 1770 1519
rect 1804 1496 2140 1519
rect 1804 1485 1866 1496
rect 713 1462 1866 1485
rect 1900 1462 2039 1496
rect 2073 1485 2140 1496
rect 2174 1485 2230 1519
rect 2264 1485 2320 1519
rect 2354 1485 2410 1519
rect 2444 1485 2500 1519
rect 2534 1485 2590 1519
rect 2624 1485 2680 1519
rect 2714 1485 2770 1519
rect 2804 1485 2860 1519
rect 2894 1485 2950 1519
rect 2984 1485 3040 1519
rect 3074 1485 3130 1519
rect 3164 1496 3300 1519
rect 3164 1485 3226 1496
rect 2073 1462 3226 1485
rect 3260 1462 3300 1496
rect -720 1406 3300 1462
rect -720 1372 -681 1406
rect -647 1372 506 1406
rect 540 1372 679 1406
rect 713 1372 1866 1406
rect 1900 1372 2039 1406
rect 2073 1372 3226 1406
rect 3260 1372 3300 1406
rect -720 1338 -474 1372
rect -440 1338 -384 1372
rect -350 1338 -294 1372
rect -260 1338 -204 1372
rect -170 1338 -114 1372
rect -80 1338 -24 1372
rect 10 1338 66 1372
rect 100 1338 156 1372
rect 190 1338 246 1372
rect 280 1338 886 1372
rect 920 1338 976 1372
rect 1010 1338 1066 1372
rect 1100 1338 1156 1372
rect 1190 1338 1246 1372
rect 1280 1338 1336 1372
rect 1370 1338 1426 1372
rect 1460 1338 1516 1372
rect 1550 1338 1606 1372
rect 1640 1338 2246 1372
rect 2280 1338 2336 1372
rect 2370 1338 2426 1372
rect 2460 1338 2516 1372
rect 2550 1338 2606 1372
rect 2640 1338 2696 1372
rect 2730 1338 2786 1372
rect 2820 1338 2876 1372
rect 2910 1338 2966 1372
rect 3000 1338 3300 1372
rect -720 1316 3300 1338
rect -720 1310 -681 1316
rect -714 1282 -681 1310
rect -647 1315 506 1316
rect -647 1310 358 1315
rect -647 1282 -615 1310
rect -714 1226 -615 1282
rect -714 1192 -681 1226
rect -647 1192 -615 1226
rect -714 1136 -615 1192
rect -714 1102 -681 1136
rect -647 1102 -615 1136
rect -714 1046 -615 1102
rect -714 1012 -681 1046
rect -647 1012 -615 1046
rect -714 956 -615 1012
rect -714 922 -681 956
rect -647 922 -615 956
rect -714 866 -615 922
rect -714 832 -681 866
rect -647 832 -615 866
rect -714 776 -615 832
rect -714 742 -681 776
rect -647 742 -615 776
rect -714 686 -615 742
rect -714 652 -681 686
rect -647 652 -615 686
rect -714 596 -615 652
rect -714 562 -681 596
rect -647 562 -615 596
rect -714 506 -615 562
rect -714 472 -681 506
rect -647 472 -615 506
rect -714 416 -615 472
rect -551 1296 -479 1310
rect -551 1262 -532 1296
rect -498 1262 -479 1296
rect -551 1206 -479 1262
rect 339 1281 358 1310
rect 392 1310 506 1315
rect 392 1281 411 1310
rect -551 1172 -532 1206
rect -498 1172 -479 1206
rect -551 1116 -479 1172
rect -551 1082 -532 1116
rect -498 1082 -479 1116
rect -551 1026 -479 1082
rect -551 992 -532 1026
rect -498 992 -479 1026
rect -551 936 -479 992
rect -551 902 -532 936
rect -498 902 -479 936
rect -551 846 -479 902
rect -551 812 -532 846
rect -498 812 -479 846
rect -551 756 -479 812
rect -551 722 -532 756
rect -498 722 -479 756
rect -551 666 -479 722
rect -551 632 -532 666
rect -498 632 -479 666
rect -551 576 -479 632
rect -551 542 -532 576
rect -498 542 -479 576
rect -417 1198 277 1257
rect -417 1164 -358 1198
rect -324 1170 -268 1198
rect -296 1164 -268 1170
rect -234 1170 -178 1198
rect -234 1164 -230 1170
rect -417 1136 -330 1164
rect -296 1136 -230 1164
rect -196 1164 -178 1170
rect -144 1170 -88 1198
rect -144 1164 -130 1170
rect -196 1136 -130 1164
rect -96 1164 -88 1170
rect -54 1170 2 1198
rect 36 1170 92 1198
rect 126 1170 182 1198
rect -54 1164 -30 1170
rect 36 1164 70 1170
rect 126 1164 170 1170
rect 216 1164 277 1198
rect -96 1136 -30 1164
rect 4 1136 70 1164
rect 104 1136 170 1164
rect 204 1136 277 1164
rect -417 1108 277 1136
rect -417 1074 -358 1108
rect -324 1074 -268 1108
rect -234 1074 -178 1108
rect -144 1074 -88 1108
rect -54 1074 2 1108
rect 36 1074 92 1108
rect 126 1074 182 1108
rect 216 1074 277 1108
rect -417 1070 277 1074
rect -417 1036 -330 1070
rect -296 1036 -230 1070
rect -196 1036 -130 1070
rect -96 1036 -30 1070
rect 4 1036 70 1070
rect 104 1036 170 1070
rect 204 1036 277 1070
rect -417 1018 277 1036
rect -417 984 -358 1018
rect -324 984 -268 1018
rect -234 984 -178 1018
rect -144 984 -88 1018
rect -54 984 2 1018
rect 36 984 92 1018
rect 126 984 182 1018
rect 216 984 277 1018
rect -417 970 277 984
rect -417 936 -330 970
rect -296 936 -230 970
rect -196 936 -130 970
rect -96 936 -30 970
rect 4 936 70 970
rect 104 936 170 970
rect 204 936 277 970
rect -417 928 277 936
rect -417 894 -358 928
rect -324 894 -268 928
rect -234 894 -178 928
rect -144 894 -88 928
rect -54 894 2 928
rect 36 894 92 928
rect 126 894 182 928
rect 216 894 277 928
rect -417 870 277 894
rect -417 838 -330 870
rect -296 838 -230 870
rect -417 804 -358 838
rect -296 836 -268 838
rect -324 804 -268 836
rect -234 836 -230 838
rect -196 838 -130 870
rect -196 836 -178 838
rect -234 804 -178 836
rect -144 836 -130 838
rect -96 838 -30 870
rect 4 838 70 870
rect 104 838 170 870
rect 204 838 277 870
rect -96 836 -88 838
rect -144 804 -88 836
rect -54 836 -30 838
rect 36 836 70 838
rect 126 836 170 838
rect -54 804 2 836
rect 36 804 92 836
rect 126 804 182 836
rect 216 804 277 838
rect -417 770 277 804
rect -417 748 -330 770
rect -296 748 -230 770
rect -417 714 -358 748
rect -296 736 -268 748
rect -324 714 -268 736
rect -234 736 -230 748
rect -196 748 -130 770
rect -196 736 -178 748
rect -234 714 -178 736
rect -144 736 -130 748
rect -96 748 -30 770
rect 4 748 70 770
rect 104 748 170 770
rect 204 748 277 770
rect -96 736 -88 748
rect -144 714 -88 736
rect -54 736 -30 748
rect 36 736 70 748
rect 126 736 170 748
rect -54 714 2 736
rect 36 714 92 736
rect 126 714 182 736
rect 216 714 277 748
rect -417 670 277 714
rect -417 658 -330 670
rect -296 658 -230 670
rect -417 624 -358 658
rect -296 636 -268 658
rect -324 624 -268 636
rect -234 636 -230 658
rect -196 658 -130 670
rect -196 636 -178 658
rect -234 624 -178 636
rect -144 636 -130 658
rect -96 658 -30 670
rect 4 658 70 670
rect 104 658 170 670
rect 204 658 277 670
rect -96 636 -88 658
rect -144 624 -88 636
rect -54 636 -30 658
rect 36 636 70 658
rect 126 636 170 658
rect -54 624 2 636
rect 36 624 92 636
rect 126 624 182 636
rect 216 624 277 658
rect -417 563 277 624
rect 339 1225 411 1281
rect 339 1191 358 1225
rect 392 1191 411 1225
rect 339 1135 411 1191
rect 339 1101 358 1135
rect 392 1101 411 1135
rect 339 1045 411 1101
rect 339 1011 358 1045
rect 392 1011 411 1045
rect 339 955 411 1011
rect 339 921 358 955
rect 392 921 411 955
rect 339 865 411 921
rect 339 831 358 865
rect 392 831 411 865
rect 339 775 411 831
rect 339 741 358 775
rect 392 741 411 775
rect 339 685 411 741
rect 339 651 358 685
rect 392 651 411 685
rect 339 595 411 651
rect -551 501 -479 542
rect 339 561 358 595
rect 392 561 411 595
rect 339 501 411 561
rect -551 482 411 501
rect -551 448 -440 482
rect -406 448 -350 482
rect -316 448 -260 482
rect -226 448 -170 482
rect -136 448 -80 482
rect -46 448 10 482
rect 44 448 100 482
rect 134 448 190 482
rect 224 448 280 482
rect 314 448 411 482
rect -551 429 411 448
rect 475 1282 506 1310
rect 540 1282 679 1316
rect 713 1315 1866 1316
rect 713 1310 1718 1315
rect 713 1282 745 1310
rect 475 1226 745 1282
rect 475 1192 506 1226
rect 540 1192 679 1226
rect 713 1192 745 1226
rect 475 1136 745 1192
rect 475 1102 506 1136
rect 540 1102 679 1136
rect 713 1102 745 1136
rect 475 1046 745 1102
rect 475 1012 506 1046
rect 540 1012 679 1046
rect 713 1012 745 1046
rect 475 956 745 1012
rect 475 922 506 956
rect 540 922 679 956
rect 713 922 745 956
rect 475 866 745 922
rect 475 832 506 866
rect 540 832 679 866
rect 713 832 745 866
rect 475 776 745 832
rect 475 742 506 776
rect 540 742 679 776
rect 713 742 745 776
rect 475 686 745 742
rect 475 652 506 686
rect 540 652 679 686
rect 713 652 745 686
rect 475 596 745 652
rect 475 562 506 596
rect 540 562 679 596
rect 713 562 745 596
rect 475 506 745 562
rect 475 472 506 506
rect 540 472 679 506
rect 713 472 745 506
rect -714 382 -681 416
rect -647 382 -615 416
rect -714 365 -615 382
rect 475 416 745 472
rect 809 1296 881 1310
rect 809 1262 828 1296
rect 862 1262 881 1296
rect 809 1206 881 1262
rect 1699 1281 1718 1310
rect 1752 1310 1866 1315
rect 1752 1281 1771 1310
rect 809 1172 828 1206
rect 862 1172 881 1206
rect 809 1116 881 1172
rect 809 1082 828 1116
rect 862 1082 881 1116
rect 809 1026 881 1082
rect 809 992 828 1026
rect 862 992 881 1026
rect 809 936 881 992
rect 809 902 828 936
rect 862 902 881 936
rect 809 846 881 902
rect 809 812 828 846
rect 862 812 881 846
rect 809 756 881 812
rect 809 722 828 756
rect 862 722 881 756
rect 809 666 881 722
rect 809 632 828 666
rect 862 632 881 666
rect 809 576 881 632
rect 809 542 828 576
rect 862 542 881 576
rect 943 1198 1637 1257
rect 943 1164 1002 1198
rect 1036 1170 1092 1198
rect 1064 1164 1092 1170
rect 1126 1170 1182 1198
rect 1126 1164 1130 1170
rect 943 1136 1030 1164
rect 1064 1136 1130 1164
rect 1164 1164 1182 1170
rect 1216 1170 1272 1198
rect 1216 1164 1230 1170
rect 1164 1136 1230 1164
rect 1264 1164 1272 1170
rect 1306 1170 1362 1198
rect 1396 1170 1452 1198
rect 1486 1170 1542 1198
rect 1306 1164 1330 1170
rect 1396 1164 1430 1170
rect 1486 1164 1530 1170
rect 1576 1164 1637 1198
rect 1264 1136 1330 1164
rect 1364 1136 1430 1164
rect 1464 1136 1530 1164
rect 1564 1136 1637 1164
rect 943 1108 1637 1136
rect 943 1074 1002 1108
rect 1036 1074 1092 1108
rect 1126 1074 1182 1108
rect 1216 1074 1272 1108
rect 1306 1074 1362 1108
rect 1396 1074 1452 1108
rect 1486 1074 1542 1108
rect 1576 1074 1637 1108
rect 943 1070 1637 1074
rect 943 1036 1030 1070
rect 1064 1036 1130 1070
rect 1164 1036 1230 1070
rect 1264 1036 1330 1070
rect 1364 1036 1430 1070
rect 1464 1036 1530 1070
rect 1564 1036 1637 1070
rect 943 1018 1637 1036
rect 943 984 1002 1018
rect 1036 984 1092 1018
rect 1126 984 1182 1018
rect 1216 984 1272 1018
rect 1306 984 1362 1018
rect 1396 984 1452 1018
rect 1486 984 1542 1018
rect 1576 984 1637 1018
rect 943 970 1637 984
rect 943 936 1030 970
rect 1064 936 1130 970
rect 1164 936 1230 970
rect 1264 936 1330 970
rect 1364 936 1430 970
rect 1464 936 1530 970
rect 1564 936 1637 970
rect 943 928 1637 936
rect 943 894 1002 928
rect 1036 894 1092 928
rect 1126 894 1182 928
rect 1216 894 1272 928
rect 1306 894 1362 928
rect 1396 894 1452 928
rect 1486 894 1542 928
rect 1576 894 1637 928
rect 943 870 1637 894
rect 943 838 1030 870
rect 1064 838 1130 870
rect 943 804 1002 838
rect 1064 836 1092 838
rect 1036 804 1092 836
rect 1126 836 1130 838
rect 1164 838 1230 870
rect 1164 836 1182 838
rect 1126 804 1182 836
rect 1216 836 1230 838
rect 1264 838 1330 870
rect 1364 838 1430 870
rect 1464 838 1530 870
rect 1564 838 1637 870
rect 1264 836 1272 838
rect 1216 804 1272 836
rect 1306 836 1330 838
rect 1396 836 1430 838
rect 1486 836 1530 838
rect 1306 804 1362 836
rect 1396 804 1452 836
rect 1486 804 1542 836
rect 1576 804 1637 838
rect 943 770 1637 804
rect 943 748 1030 770
rect 1064 748 1130 770
rect 943 714 1002 748
rect 1064 736 1092 748
rect 1036 714 1092 736
rect 1126 736 1130 748
rect 1164 748 1230 770
rect 1164 736 1182 748
rect 1126 714 1182 736
rect 1216 736 1230 748
rect 1264 748 1330 770
rect 1364 748 1430 770
rect 1464 748 1530 770
rect 1564 748 1637 770
rect 1264 736 1272 748
rect 1216 714 1272 736
rect 1306 736 1330 748
rect 1396 736 1430 748
rect 1486 736 1530 748
rect 1306 714 1362 736
rect 1396 714 1452 736
rect 1486 714 1542 736
rect 1576 714 1637 748
rect 943 670 1637 714
rect 943 658 1030 670
rect 1064 658 1130 670
rect 943 624 1002 658
rect 1064 636 1092 658
rect 1036 624 1092 636
rect 1126 636 1130 658
rect 1164 658 1230 670
rect 1164 636 1182 658
rect 1126 624 1182 636
rect 1216 636 1230 658
rect 1264 658 1330 670
rect 1364 658 1430 670
rect 1464 658 1530 670
rect 1564 658 1637 670
rect 1264 636 1272 658
rect 1216 624 1272 636
rect 1306 636 1330 658
rect 1396 636 1430 658
rect 1486 636 1530 658
rect 1306 624 1362 636
rect 1396 624 1452 636
rect 1486 624 1542 636
rect 1576 624 1637 658
rect 943 563 1637 624
rect 1699 1225 1771 1281
rect 1699 1191 1718 1225
rect 1752 1191 1771 1225
rect 1699 1135 1771 1191
rect 1699 1101 1718 1135
rect 1752 1101 1771 1135
rect 1699 1045 1771 1101
rect 1699 1011 1718 1045
rect 1752 1011 1771 1045
rect 1699 955 1771 1011
rect 1699 921 1718 955
rect 1752 921 1771 955
rect 1699 865 1771 921
rect 1699 831 1718 865
rect 1752 831 1771 865
rect 1699 775 1771 831
rect 1699 741 1718 775
rect 1752 741 1771 775
rect 1699 685 1771 741
rect 1699 651 1718 685
rect 1752 651 1771 685
rect 1699 595 1771 651
rect 809 501 881 542
rect 1699 561 1718 595
rect 1752 561 1771 595
rect 1699 501 1771 561
rect 809 482 1771 501
rect 809 448 920 482
rect 954 448 1010 482
rect 1044 448 1100 482
rect 1134 448 1190 482
rect 1224 448 1280 482
rect 1314 448 1370 482
rect 1404 448 1460 482
rect 1494 448 1550 482
rect 1584 448 1640 482
rect 1674 448 1771 482
rect 809 429 1771 448
rect 1835 1282 1866 1310
rect 1900 1282 2039 1316
rect 2073 1315 3226 1316
rect 2073 1310 3078 1315
rect 2073 1282 2105 1310
rect 1835 1226 2105 1282
rect 1835 1192 1866 1226
rect 1900 1192 2039 1226
rect 2073 1192 2105 1226
rect 1835 1136 2105 1192
rect 1835 1102 1866 1136
rect 1900 1102 2039 1136
rect 2073 1102 2105 1136
rect 1835 1046 2105 1102
rect 1835 1012 1866 1046
rect 1900 1012 2039 1046
rect 2073 1012 2105 1046
rect 1835 956 2105 1012
rect 1835 922 1866 956
rect 1900 922 2039 956
rect 2073 922 2105 956
rect 1835 866 2105 922
rect 1835 832 1866 866
rect 1900 832 2039 866
rect 2073 832 2105 866
rect 1835 776 2105 832
rect 1835 742 1866 776
rect 1900 742 2039 776
rect 2073 742 2105 776
rect 1835 686 2105 742
rect 1835 652 1866 686
rect 1900 652 2039 686
rect 2073 652 2105 686
rect 1835 596 2105 652
rect 1835 562 1866 596
rect 1900 562 2039 596
rect 2073 562 2105 596
rect 1835 506 2105 562
rect 1835 472 1866 506
rect 1900 472 2039 506
rect 2073 472 2105 506
rect 475 382 506 416
rect 540 382 679 416
rect 713 382 745 416
rect 475 365 745 382
rect 1835 416 2105 472
rect 2169 1296 2241 1310
rect 2169 1262 2188 1296
rect 2222 1262 2241 1296
rect 2169 1206 2241 1262
rect 3059 1281 3078 1310
rect 3112 1310 3226 1315
rect 3112 1281 3131 1310
rect 2169 1172 2188 1206
rect 2222 1172 2241 1206
rect 2169 1116 2241 1172
rect 2169 1082 2188 1116
rect 2222 1082 2241 1116
rect 2169 1026 2241 1082
rect 2169 992 2188 1026
rect 2222 992 2241 1026
rect 2169 936 2241 992
rect 2169 902 2188 936
rect 2222 902 2241 936
rect 2169 846 2241 902
rect 2169 812 2188 846
rect 2222 812 2241 846
rect 2169 756 2241 812
rect 2169 722 2188 756
rect 2222 722 2241 756
rect 2169 666 2241 722
rect 2169 632 2188 666
rect 2222 632 2241 666
rect 2169 576 2241 632
rect 2169 542 2188 576
rect 2222 542 2241 576
rect 2303 1198 2997 1257
rect 2303 1164 2362 1198
rect 2396 1170 2452 1198
rect 2424 1164 2452 1170
rect 2486 1170 2542 1198
rect 2486 1164 2490 1170
rect 2303 1136 2390 1164
rect 2424 1136 2490 1164
rect 2524 1164 2542 1170
rect 2576 1170 2632 1198
rect 2576 1164 2590 1170
rect 2524 1136 2590 1164
rect 2624 1164 2632 1170
rect 2666 1170 2722 1198
rect 2756 1170 2812 1198
rect 2846 1170 2902 1198
rect 2666 1164 2690 1170
rect 2756 1164 2790 1170
rect 2846 1164 2890 1170
rect 2936 1164 2997 1198
rect 2624 1136 2690 1164
rect 2724 1136 2790 1164
rect 2824 1136 2890 1164
rect 2924 1136 2997 1164
rect 2303 1108 2997 1136
rect 2303 1074 2362 1108
rect 2396 1074 2452 1108
rect 2486 1074 2542 1108
rect 2576 1074 2632 1108
rect 2666 1074 2722 1108
rect 2756 1074 2812 1108
rect 2846 1074 2902 1108
rect 2936 1074 2997 1108
rect 2303 1070 2997 1074
rect 2303 1036 2390 1070
rect 2424 1036 2490 1070
rect 2524 1036 2590 1070
rect 2624 1036 2690 1070
rect 2724 1036 2790 1070
rect 2824 1036 2890 1070
rect 2924 1036 2997 1070
rect 2303 1018 2997 1036
rect 2303 984 2362 1018
rect 2396 984 2452 1018
rect 2486 984 2542 1018
rect 2576 984 2632 1018
rect 2666 984 2722 1018
rect 2756 984 2812 1018
rect 2846 984 2902 1018
rect 2936 984 2997 1018
rect 2303 970 2997 984
rect 2303 936 2390 970
rect 2424 936 2490 970
rect 2524 936 2590 970
rect 2624 936 2690 970
rect 2724 936 2790 970
rect 2824 936 2890 970
rect 2924 936 2997 970
rect 2303 928 2997 936
rect 2303 894 2362 928
rect 2396 894 2452 928
rect 2486 894 2542 928
rect 2576 894 2632 928
rect 2666 894 2722 928
rect 2756 894 2812 928
rect 2846 894 2902 928
rect 2936 894 2997 928
rect 2303 870 2997 894
rect 2303 838 2390 870
rect 2424 838 2490 870
rect 2303 804 2362 838
rect 2424 836 2452 838
rect 2396 804 2452 836
rect 2486 836 2490 838
rect 2524 838 2590 870
rect 2524 836 2542 838
rect 2486 804 2542 836
rect 2576 836 2590 838
rect 2624 838 2690 870
rect 2724 838 2790 870
rect 2824 838 2890 870
rect 2924 838 2997 870
rect 2624 836 2632 838
rect 2576 804 2632 836
rect 2666 836 2690 838
rect 2756 836 2790 838
rect 2846 836 2890 838
rect 2666 804 2722 836
rect 2756 804 2812 836
rect 2846 804 2902 836
rect 2936 804 2997 838
rect 2303 770 2997 804
rect 2303 748 2390 770
rect 2424 748 2490 770
rect 2303 714 2362 748
rect 2424 736 2452 748
rect 2396 714 2452 736
rect 2486 736 2490 748
rect 2524 748 2590 770
rect 2524 736 2542 748
rect 2486 714 2542 736
rect 2576 736 2590 748
rect 2624 748 2690 770
rect 2724 748 2790 770
rect 2824 748 2890 770
rect 2924 748 2997 770
rect 2624 736 2632 748
rect 2576 714 2632 736
rect 2666 736 2690 748
rect 2756 736 2790 748
rect 2846 736 2890 748
rect 2666 714 2722 736
rect 2756 714 2812 736
rect 2846 714 2902 736
rect 2936 714 2997 748
rect 2303 670 2997 714
rect 2303 658 2390 670
rect 2424 658 2490 670
rect 2303 624 2362 658
rect 2424 636 2452 658
rect 2396 624 2452 636
rect 2486 636 2490 658
rect 2524 658 2590 670
rect 2524 636 2542 658
rect 2486 624 2542 636
rect 2576 636 2590 658
rect 2624 658 2690 670
rect 2724 658 2790 670
rect 2824 658 2890 670
rect 2924 658 2997 670
rect 2624 636 2632 658
rect 2576 624 2632 636
rect 2666 636 2690 658
rect 2756 636 2790 658
rect 2846 636 2890 658
rect 2666 624 2722 636
rect 2756 624 2812 636
rect 2846 624 2902 636
rect 2936 624 2997 658
rect 2303 563 2997 624
rect 3059 1225 3131 1281
rect 3059 1191 3078 1225
rect 3112 1191 3131 1225
rect 3059 1135 3131 1191
rect 3059 1101 3078 1135
rect 3112 1101 3131 1135
rect 3059 1045 3131 1101
rect 3059 1011 3078 1045
rect 3112 1011 3131 1045
rect 3059 955 3131 1011
rect 3059 921 3078 955
rect 3112 921 3131 955
rect 3059 865 3131 921
rect 3059 831 3078 865
rect 3112 831 3131 865
rect 3059 775 3131 831
rect 3059 741 3078 775
rect 3112 741 3131 775
rect 3059 685 3131 741
rect 3059 651 3078 685
rect 3112 651 3131 685
rect 3059 595 3131 651
rect 2169 501 2241 542
rect 3059 561 3078 595
rect 3112 561 3131 595
rect 3059 501 3131 561
rect 2169 482 3131 501
rect 2169 448 2280 482
rect 2314 448 2370 482
rect 2404 448 2460 482
rect 2494 448 2550 482
rect 2584 448 2640 482
rect 2674 448 2730 482
rect 2764 448 2820 482
rect 2854 448 2910 482
rect 2944 448 3000 482
rect 3034 448 3131 482
rect 2169 429 3131 448
rect 3195 1282 3226 1310
rect 3260 1310 3300 1316
rect 3260 1282 3294 1310
rect 3195 1226 3294 1282
rect 3195 1192 3226 1226
rect 3260 1192 3294 1226
rect 3195 1136 3294 1192
rect 3195 1102 3226 1136
rect 3260 1102 3294 1136
rect 3195 1046 3294 1102
rect 3195 1012 3226 1046
rect 3260 1012 3294 1046
rect 3195 956 3294 1012
rect 3195 922 3226 956
rect 3260 922 3294 956
rect 3195 866 3294 922
rect 3195 832 3226 866
rect 3260 832 3294 866
rect 3195 776 3294 832
rect 3195 742 3226 776
rect 3260 742 3294 776
rect 3195 686 3294 742
rect 3195 652 3226 686
rect 3260 652 3294 686
rect 3195 596 3294 652
rect 3195 562 3226 596
rect 3260 562 3294 596
rect 3195 506 3294 562
rect 3195 472 3226 506
rect 3260 472 3294 506
rect 1835 382 1866 416
rect 1900 382 2039 416
rect 2073 382 2105 416
rect 1835 365 2105 382
rect 3195 416 3294 472
rect 3195 382 3226 416
rect 3260 382 3294 416
rect 3195 365 3294 382
rect -714 332 3294 365
rect -714 298 -580 332
rect -546 298 -490 332
rect -456 298 -400 332
rect -366 298 -310 332
rect -276 298 -220 332
rect -186 298 -130 332
rect -96 298 -40 332
rect -6 298 50 332
rect 84 298 140 332
rect 174 298 230 332
rect 264 298 320 332
rect 354 298 410 332
rect 444 298 780 332
rect 814 298 870 332
rect 904 298 960 332
rect 994 298 1050 332
rect 1084 298 1140 332
rect 1174 298 1230 332
rect 1264 298 1320 332
rect 1354 298 1410 332
rect 1444 298 1500 332
rect 1534 298 1590 332
rect 1624 298 1680 332
rect 1714 298 1770 332
rect 1804 298 2140 332
rect 2174 298 2230 332
rect 2264 298 2320 332
rect 2354 298 2410 332
rect 2444 298 2500 332
rect 2534 298 2590 332
rect 2624 298 2680 332
rect 2714 298 2770 332
rect 2804 298 2860 332
rect 2894 298 2950 332
rect 2984 298 3040 332
rect 3074 298 3130 332
rect 3164 298 3294 332
rect -714 266 3294 298
rect 570 200 650 266
rect 1930 200 2010 266
rect -1827 149 -1731 183
rect -1139 149 -1043 183
rect -1827 87 -1793 149
rect -2940 -382 -2844 -348
rect -2252 -382 -2156 -348
rect -2940 -444 -2906 -382
rect -3727 -781 -3631 -747
rect -3371 -781 -3275 -747
rect -3727 -843 -3693 -781
rect -3309 -843 -3275 -781
rect -3727 -2233 -3693 -2171
rect -3540 -2233 -3460 -2220
rect -3309 -2233 -3275 -2171
rect -3727 -2267 -3631 -2233
rect -3371 -2267 -3275 -2233
rect -2190 -444 -2156 -382
rect -2940 -2236 -2906 -2174
rect -2750 -2236 -2670 -2220
rect -2190 -2236 -2156 -2174
rect -3540 -2280 -3520 -2267
rect -3480 -2280 -3460 -2267
rect -2940 -2270 -2844 -2236
rect -2252 -2270 -2156 -2236
rect -1077 87 -1043 149
rect -1827 -2233 -1793 -2171
rect -720 159 3300 200
rect -720 136 -580 159
rect -720 102 -681 136
rect -647 125 -580 136
rect -546 125 -490 159
rect -456 125 -400 159
rect -366 125 -310 159
rect -276 125 -220 159
rect -186 125 -130 159
rect -96 125 -40 159
rect -6 125 50 159
rect 84 125 140 159
rect 174 125 230 159
rect 264 125 320 159
rect 354 125 410 159
rect 444 136 780 159
rect 444 125 506 136
rect -647 102 506 125
rect 540 102 679 136
rect 713 125 780 136
rect 814 125 870 159
rect 904 125 960 159
rect 994 125 1050 159
rect 1084 125 1140 159
rect 1174 125 1230 159
rect 1264 125 1320 159
rect 1354 125 1410 159
rect 1444 125 1500 159
rect 1534 125 1590 159
rect 1624 125 1680 159
rect 1714 125 1770 159
rect 1804 136 2140 159
rect 1804 125 1866 136
rect 713 102 1866 125
rect 1900 102 2039 136
rect 2073 125 2140 136
rect 2174 125 2230 159
rect 2264 125 2320 159
rect 2354 125 2410 159
rect 2444 125 2500 159
rect 2534 125 2590 159
rect 2624 125 2680 159
rect 2714 125 2770 159
rect 2804 125 2860 159
rect 2894 125 2950 159
rect 2984 125 3040 159
rect 3074 125 3130 159
rect 3164 136 3300 159
rect 3164 125 3226 136
rect 2073 102 3226 125
rect 3260 102 3300 136
rect -720 46 3300 102
rect -720 12 -681 46
rect -647 12 506 46
rect 540 12 679 46
rect 713 12 1866 46
rect 1900 12 2039 46
rect 2073 12 3226 46
rect 3260 12 3300 46
rect -720 -22 -474 12
rect -440 -22 -384 12
rect -350 -22 -294 12
rect -260 -22 -204 12
rect -170 -22 -114 12
rect -80 -22 -24 12
rect 10 -22 66 12
rect 100 -22 156 12
rect 190 -22 246 12
rect 280 -22 886 12
rect 920 -22 976 12
rect 1010 -22 1066 12
rect 1100 -22 1156 12
rect 1190 -22 1246 12
rect 1280 -22 1336 12
rect 1370 -22 1426 12
rect 1460 -22 1516 12
rect 1550 -22 1606 12
rect 1640 -22 2246 12
rect 2280 -22 2336 12
rect 2370 -22 2426 12
rect 2460 -22 2516 12
rect 2550 -22 2606 12
rect 2640 -22 2696 12
rect 2730 -22 2786 12
rect 2820 -22 2876 12
rect 2910 -22 2966 12
rect 3000 -22 3300 12
rect -720 -44 3300 -22
rect -720 -50 -681 -44
rect -714 -78 -681 -50
rect -647 -45 506 -44
rect -647 -50 358 -45
rect -647 -78 -615 -50
rect -714 -134 -615 -78
rect -714 -168 -681 -134
rect -647 -168 -615 -134
rect -714 -224 -615 -168
rect -714 -258 -681 -224
rect -647 -258 -615 -224
rect -714 -314 -615 -258
rect -714 -348 -681 -314
rect -647 -348 -615 -314
rect -714 -404 -615 -348
rect -714 -438 -681 -404
rect -647 -438 -615 -404
rect -714 -494 -615 -438
rect -714 -528 -681 -494
rect -647 -528 -615 -494
rect -714 -584 -615 -528
rect -714 -618 -681 -584
rect -647 -618 -615 -584
rect -714 -674 -615 -618
rect -714 -708 -681 -674
rect -647 -708 -615 -674
rect -714 -764 -615 -708
rect -714 -798 -681 -764
rect -647 -798 -615 -764
rect -714 -854 -615 -798
rect -714 -888 -681 -854
rect -647 -888 -615 -854
rect -714 -944 -615 -888
rect -551 -64 -479 -50
rect -551 -98 -532 -64
rect -498 -98 -479 -64
rect -551 -154 -479 -98
rect 339 -79 358 -50
rect 392 -50 506 -45
rect 392 -79 411 -50
rect -551 -188 -532 -154
rect -498 -188 -479 -154
rect -551 -244 -479 -188
rect -551 -278 -532 -244
rect -498 -278 -479 -244
rect -551 -334 -479 -278
rect -551 -368 -532 -334
rect -498 -368 -479 -334
rect -551 -424 -479 -368
rect -551 -458 -532 -424
rect -498 -458 -479 -424
rect -551 -514 -479 -458
rect -551 -548 -532 -514
rect -498 -548 -479 -514
rect -551 -604 -479 -548
rect -551 -638 -532 -604
rect -498 -638 -479 -604
rect -551 -694 -479 -638
rect -551 -728 -532 -694
rect -498 -728 -479 -694
rect -551 -784 -479 -728
rect -551 -818 -532 -784
rect -498 -818 -479 -784
rect -417 -162 277 -103
rect -417 -196 -358 -162
rect -324 -190 -268 -162
rect -296 -196 -268 -190
rect -234 -190 -178 -162
rect -234 -196 -230 -190
rect -417 -224 -330 -196
rect -296 -224 -230 -196
rect -196 -196 -178 -190
rect -144 -190 -88 -162
rect -144 -196 -130 -190
rect -196 -224 -130 -196
rect -96 -196 -88 -190
rect -54 -190 2 -162
rect 36 -190 92 -162
rect 126 -190 182 -162
rect -54 -196 -30 -190
rect 36 -196 70 -190
rect 126 -196 170 -190
rect 216 -196 277 -162
rect -96 -224 -30 -196
rect 4 -224 70 -196
rect 104 -224 170 -196
rect 204 -224 277 -196
rect -417 -252 277 -224
rect -417 -286 -358 -252
rect -324 -286 -268 -252
rect -234 -286 -178 -252
rect -144 -286 -88 -252
rect -54 -286 2 -252
rect 36 -286 92 -252
rect 126 -286 182 -252
rect 216 -286 277 -252
rect -417 -290 277 -286
rect -417 -324 -330 -290
rect -296 -324 -230 -290
rect -196 -324 -130 -290
rect -96 -324 -30 -290
rect 4 -324 70 -290
rect 104 -324 170 -290
rect 204 -324 277 -290
rect -417 -342 277 -324
rect -417 -376 -358 -342
rect -324 -376 -268 -342
rect -234 -376 -178 -342
rect -144 -376 -88 -342
rect -54 -376 2 -342
rect 36 -376 92 -342
rect 126 -376 182 -342
rect 216 -376 277 -342
rect -417 -390 277 -376
rect -417 -424 -330 -390
rect -296 -424 -230 -390
rect -196 -424 -130 -390
rect -96 -424 -30 -390
rect 4 -424 70 -390
rect 104 -424 170 -390
rect 204 -424 277 -390
rect -417 -432 277 -424
rect -417 -466 -358 -432
rect -324 -466 -268 -432
rect -234 -466 -178 -432
rect -144 -466 -88 -432
rect -54 -466 2 -432
rect 36 -466 92 -432
rect 126 -466 182 -432
rect 216 -466 277 -432
rect -417 -490 277 -466
rect -417 -522 -330 -490
rect -296 -522 -230 -490
rect -417 -556 -358 -522
rect -296 -524 -268 -522
rect -324 -556 -268 -524
rect -234 -524 -230 -522
rect -196 -522 -130 -490
rect -196 -524 -178 -522
rect -234 -556 -178 -524
rect -144 -524 -130 -522
rect -96 -522 -30 -490
rect 4 -522 70 -490
rect 104 -522 170 -490
rect 204 -522 277 -490
rect -96 -524 -88 -522
rect -144 -556 -88 -524
rect -54 -524 -30 -522
rect 36 -524 70 -522
rect 126 -524 170 -522
rect -54 -556 2 -524
rect 36 -556 92 -524
rect 126 -556 182 -524
rect 216 -556 277 -522
rect -417 -590 277 -556
rect -417 -612 -330 -590
rect -296 -612 -230 -590
rect -417 -646 -358 -612
rect -296 -624 -268 -612
rect -324 -646 -268 -624
rect -234 -624 -230 -612
rect -196 -612 -130 -590
rect -196 -624 -178 -612
rect -234 -646 -178 -624
rect -144 -624 -130 -612
rect -96 -612 -30 -590
rect 4 -612 70 -590
rect 104 -612 170 -590
rect 204 -612 277 -590
rect -96 -624 -88 -612
rect -144 -646 -88 -624
rect -54 -624 -30 -612
rect 36 -624 70 -612
rect 126 -624 170 -612
rect -54 -646 2 -624
rect 36 -646 92 -624
rect 126 -646 182 -624
rect 216 -646 277 -612
rect -417 -690 277 -646
rect -417 -702 -330 -690
rect -296 -702 -230 -690
rect -417 -736 -358 -702
rect -296 -724 -268 -702
rect -324 -736 -268 -724
rect -234 -724 -230 -702
rect -196 -702 -130 -690
rect -196 -724 -178 -702
rect -234 -736 -178 -724
rect -144 -724 -130 -702
rect -96 -702 -30 -690
rect 4 -702 70 -690
rect 104 -702 170 -690
rect 204 -702 277 -690
rect -96 -724 -88 -702
rect -144 -736 -88 -724
rect -54 -724 -30 -702
rect 36 -724 70 -702
rect 126 -724 170 -702
rect -54 -736 2 -724
rect 36 -736 92 -724
rect 126 -736 182 -724
rect 216 -736 277 -702
rect -417 -797 277 -736
rect 339 -135 411 -79
rect 339 -169 358 -135
rect 392 -169 411 -135
rect 339 -225 411 -169
rect 339 -259 358 -225
rect 392 -259 411 -225
rect 339 -315 411 -259
rect 339 -349 358 -315
rect 392 -349 411 -315
rect 339 -405 411 -349
rect 339 -439 358 -405
rect 392 -439 411 -405
rect 339 -495 411 -439
rect 339 -529 358 -495
rect 392 -529 411 -495
rect 339 -585 411 -529
rect 339 -619 358 -585
rect 392 -619 411 -585
rect 339 -675 411 -619
rect 339 -709 358 -675
rect 392 -709 411 -675
rect 339 -765 411 -709
rect -551 -859 -479 -818
rect 339 -799 358 -765
rect 392 -799 411 -765
rect 339 -859 411 -799
rect -551 -878 411 -859
rect -551 -912 -440 -878
rect -406 -912 -350 -878
rect -316 -912 -260 -878
rect -226 -912 -170 -878
rect -136 -912 -80 -878
rect -46 -912 10 -878
rect 44 -912 100 -878
rect 134 -912 190 -878
rect 224 -912 280 -878
rect 314 -912 411 -878
rect -551 -931 411 -912
rect 475 -78 506 -50
rect 540 -78 679 -44
rect 713 -45 1866 -44
rect 713 -50 1718 -45
rect 713 -78 745 -50
rect 475 -134 745 -78
rect 475 -168 506 -134
rect 540 -168 679 -134
rect 713 -168 745 -134
rect 475 -224 745 -168
rect 475 -258 506 -224
rect 540 -258 679 -224
rect 713 -258 745 -224
rect 475 -314 745 -258
rect 475 -348 506 -314
rect 540 -348 679 -314
rect 713 -348 745 -314
rect 475 -404 745 -348
rect 475 -438 506 -404
rect 540 -438 679 -404
rect 713 -438 745 -404
rect 475 -494 745 -438
rect 475 -528 506 -494
rect 540 -528 679 -494
rect 713 -528 745 -494
rect 475 -584 745 -528
rect 475 -618 506 -584
rect 540 -618 679 -584
rect 713 -618 745 -584
rect 475 -674 745 -618
rect 475 -708 506 -674
rect 540 -708 679 -674
rect 713 -708 745 -674
rect 475 -764 745 -708
rect 475 -798 506 -764
rect 540 -798 679 -764
rect 713 -798 745 -764
rect 475 -854 745 -798
rect 475 -888 506 -854
rect 540 -888 679 -854
rect 713 -888 745 -854
rect -714 -978 -681 -944
rect -647 -978 -615 -944
rect -714 -995 -615 -978
rect 475 -944 745 -888
rect 809 -64 881 -50
rect 809 -98 828 -64
rect 862 -98 881 -64
rect 809 -154 881 -98
rect 1699 -79 1718 -50
rect 1752 -50 1866 -45
rect 1752 -79 1771 -50
rect 809 -188 828 -154
rect 862 -188 881 -154
rect 809 -244 881 -188
rect 809 -278 828 -244
rect 862 -278 881 -244
rect 809 -334 881 -278
rect 809 -368 828 -334
rect 862 -368 881 -334
rect 809 -424 881 -368
rect 809 -458 828 -424
rect 862 -458 881 -424
rect 809 -514 881 -458
rect 809 -548 828 -514
rect 862 -548 881 -514
rect 809 -604 881 -548
rect 809 -638 828 -604
rect 862 -638 881 -604
rect 809 -694 881 -638
rect 809 -728 828 -694
rect 862 -728 881 -694
rect 809 -784 881 -728
rect 809 -818 828 -784
rect 862 -818 881 -784
rect 943 -162 1637 -103
rect 943 -196 1002 -162
rect 1036 -190 1092 -162
rect 1064 -196 1092 -190
rect 1126 -190 1182 -162
rect 1126 -196 1130 -190
rect 943 -224 1030 -196
rect 1064 -224 1130 -196
rect 1164 -196 1182 -190
rect 1216 -190 1272 -162
rect 1216 -196 1230 -190
rect 1164 -224 1230 -196
rect 1264 -196 1272 -190
rect 1306 -190 1362 -162
rect 1396 -190 1452 -162
rect 1486 -190 1542 -162
rect 1306 -196 1330 -190
rect 1396 -196 1430 -190
rect 1486 -196 1530 -190
rect 1576 -196 1637 -162
rect 1264 -224 1330 -196
rect 1364 -224 1430 -196
rect 1464 -224 1530 -196
rect 1564 -224 1637 -196
rect 943 -252 1637 -224
rect 943 -286 1002 -252
rect 1036 -286 1092 -252
rect 1126 -286 1182 -252
rect 1216 -286 1272 -252
rect 1306 -286 1362 -252
rect 1396 -286 1452 -252
rect 1486 -286 1542 -252
rect 1576 -286 1637 -252
rect 943 -290 1637 -286
rect 943 -324 1030 -290
rect 1064 -324 1130 -290
rect 1164 -324 1230 -290
rect 1264 -324 1330 -290
rect 1364 -324 1430 -290
rect 1464 -324 1530 -290
rect 1564 -324 1637 -290
rect 943 -342 1637 -324
rect 943 -376 1002 -342
rect 1036 -376 1092 -342
rect 1126 -376 1182 -342
rect 1216 -376 1272 -342
rect 1306 -376 1362 -342
rect 1396 -376 1452 -342
rect 1486 -376 1542 -342
rect 1576 -376 1637 -342
rect 943 -390 1637 -376
rect 943 -424 1030 -390
rect 1064 -424 1130 -390
rect 1164 -424 1230 -390
rect 1264 -424 1330 -390
rect 1364 -424 1430 -390
rect 1464 -424 1530 -390
rect 1564 -424 1637 -390
rect 943 -432 1637 -424
rect 943 -466 1002 -432
rect 1036 -466 1092 -432
rect 1126 -466 1182 -432
rect 1216 -466 1272 -432
rect 1306 -466 1362 -432
rect 1396 -466 1452 -432
rect 1486 -466 1542 -432
rect 1576 -466 1637 -432
rect 943 -490 1637 -466
rect 943 -522 1030 -490
rect 1064 -522 1130 -490
rect 943 -556 1002 -522
rect 1064 -524 1092 -522
rect 1036 -556 1092 -524
rect 1126 -524 1130 -522
rect 1164 -522 1230 -490
rect 1164 -524 1182 -522
rect 1126 -556 1182 -524
rect 1216 -524 1230 -522
rect 1264 -522 1330 -490
rect 1364 -522 1430 -490
rect 1464 -522 1530 -490
rect 1564 -522 1637 -490
rect 1264 -524 1272 -522
rect 1216 -556 1272 -524
rect 1306 -524 1330 -522
rect 1396 -524 1430 -522
rect 1486 -524 1530 -522
rect 1306 -556 1362 -524
rect 1396 -556 1452 -524
rect 1486 -556 1542 -524
rect 1576 -556 1637 -522
rect 943 -590 1637 -556
rect 943 -612 1030 -590
rect 1064 -612 1130 -590
rect 943 -646 1002 -612
rect 1064 -624 1092 -612
rect 1036 -646 1092 -624
rect 1126 -624 1130 -612
rect 1164 -612 1230 -590
rect 1164 -624 1182 -612
rect 1126 -646 1182 -624
rect 1216 -624 1230 -612
rect 1264 -612 1330 -590
rect 1364 -612 1430 -590
rect 1464 -612 1530 -590
rect 1564 -612 1637 -590
rect 1264 -624 1272 -612
rect 1216 -646 1272 -624
rect 1306 -624 1330 -612
rect 1396 -624 1430 -612
rect 1486 -624 1530 -612
rect 1306 -646 1362 -624
rect 1396 -646 1452 -624
rect 1486 -646 1542 -624
rect 1576 -646 1637 -612
rect 943 -690 1637 -646
rect 943 -702 1030 -690
rect 1064 -702 1130 -690
rect 943 -736 1002 -702
rect 1064 -724 1092 -702
rect 1036 -736 1092 -724
rect 1126 -724 1130 -702
rect 1164 -702 1230 -690
rect 1164 -724 1182 -702
rect 1126 -736 1182 -724
rect 1216 -724 1230 -702
rect 1264 -702 1330 -690
rect 1364 -702 1430 -690
rect 1464 -702 1530 -690
rect 1564 -702 1637 -690
rect 1264 -724 1272 -702
rect 1216 -736 1272 -724
rect 1306 -724 1330 -702
rect 1396 -724 1430 -702
rect 1486 -724 1530 -702
rect 1306 -736 1362 -724
rect 1396 -736 1452 -724
rect 1486 -736 1542 -724
rect 1576 -736 1637 -702
rect 943 -797 1637 -736
rect 1699 -135 1771 -79
rect 1699 -169 1718 -135
rect 1752 -169 1771 -135
rect 1699 -225 1771 -169
rect 1699 -259 1718 -225
rect 1752 -259 1771 -225
rect 1699 -315 1771 -259
rect 1699 -349 1718 -315
rect 1752 -349 1771 -315
rect 1699 -405 1771 -349
rect 1699 -439 1718 -405
rect 1752 -439 1771 -405
rect 1699 -495 1771 -439
rect 1699 -529 1718 -495
rect 1752 -529 1771 -495
rect 1699 -585 1771 -529
rect 1699 -619 1718 -585
rect 1752 -619 1771 -585
rect 1699 -675 1771 -619
rect 1699 -709 1718 -675
rect 1752 -709 1771 -675
rect 1699 -765 1771 -709
rect 809 -859 881 -818
rect 1699 -799 1718 -765
rect 1752 -799 1771 -765
rect 1699 -859 1771 -799
rect 809 -878 1771 -859
rect 809 -912 920 -878
rect 954 -912 1010 -878
rect 1044 -912 1100 -878
rect 1134 -912 1190 -878
rect 1224 -912 1280 -878
rect 1314 -912 1370 -878
rect 1404 -912 1460 -878
rect 1494 -912 1550 -878
rect 1584 -912 1640 -878
rect 1674 -912 1771 -878
rect 809 -931 1771 -912
rect 1835 -78 1866 -50
rect 1900 -78 2039 -44
rect 2073 -45 3226 -44
rect 2073 -50 3078 -45
rect 2073 -78 2105 -50
rect 1835 -134 2105 -78
rect 1835 -168 1866 -134
rect 1900 -168 2039 -134
rect 2073 -168 2105 -134
rect 1835 -224 2105 -168
rect 1835 -258 1866 -224
rect 1900 -258 2039 -224
rect 2073 -258 2105 -224
rect 1835 -314 2105 -258
rect 1835 -348 1866 -314
rect 1900 -348 2039 -314
rect 2073 -348 2105 -314
rect 1835 -404 2105 -348
rect 1835 -438 1866 -404
rect 1900 -438 2039 -404
rect 2073 -438 2105 -404
rect 1835 -494 2105 -438
rect 1835 -528 1866 -494
rect 1900 -528 2039 -494
rect 2073 -528 2105 -494
rect 1835 -584 2105 -528
rect 1835 -618 1866 -584
rect 1900 -618 2039 -584
rect 2073 -618 2105 -584
rect 1835 -674 2105 -618
rect 1835 -708 1866 -674
rect 1900 -708 2039 -674
rect 2073 -708 2105 -674
rect 1835 -764 2105 -708
rect 1835 -798 1866 -764
rect 1900 -798 2039 -764
rect 2073 -798 2105 -764
rect 1835 -854 2105 -798
rect 1835 -888 1866 -854
rect 1900 -888 2039 -854
rect 2073 -888 2105 -854
rect 475 -978 506 -944
rect 540 -978 679 -944
rect 713 -978 745 -944
rect 475 -995 745 -978
rect 1835 -944 2105 -888
rect 2169 -64 2241 -50
rect 2169 -98 2188 -64
rect 2222 -98 2241 -64
rect 2169 -154 2241 -98
rect 3059 -79 3078 -50
rect 3112 -50 3226 -45
rect 3112 -79 3131 -50
rect 2169 -188 2188 -154
rect 2222 -188 2241 -154
rect 2169 -244 2241 -188
rect 2169 -278 2188 -244
rect 2222 -278 2241 -244
rect 2169 -334 2241 -278
rect 2169 -368 2188 -334
rect 2222 -368 2241 -334
rect 2169 -424 2241 -368
rect 2169 -458 2188 -424
rect 2222 -458 2241 -424
rect 2169 -514 2241 -458
rect 2169 -548 2188 -514
rect 2222 -548 2241 -514
rect 2169 -604 2241 -548
rect 2169 -638 2188 -604
rect 2222 -638 2241 -604
rect 2169 -694 2241 -638
rect 2169 -728 2188 -694
rect 2222 -728 2241 -694
rect 2169 -784 2241 -728
rect 2169 -818 2188 -784
rect 2222 -818 2241 -784
rect 2303 -162 2997 -103
rect 2303 -196 2362 -162
rect 2396 -190 2452 -162
rect 2424 -196 2452 -190
rect 2486 -190 2542 -162
rect 2486 -196 2490 -190
rect 2303 -224 2390 -196
rect 2424 -224 2490 -196
rect 2524 -196 2542 -190
rect 2576 -190 2632 -162
rect 2576 -196 2590 -190
rect 2524 -224 2590 -196
rect 2624 -196 2632 -190
rect 2666 -190 2722 -162
rect 2756 -190 2812 -162
rect 2846 -190 2902 -162
rect 2666 -196 2690 -190
rect 2756 -196 2790 -190
rect 2846 -196 2890 -190
rect 2936 -196 2997 -162
rect 2624 -224 2690 -196
rect 2724 -224 2790 -196
rect 2824 -224 2890 -196
rect 2924 -224 2997 -196
rect 2303 -252 2997 -224
rect 2303 -286 2362 -252
rect 2396 -286 2452 -252
rect 2486 -286 2542 -252
rect 2576 -286 2632 -252
rect 2666 -286 2722 -252
rect 2756 -286 2812 -252
rect 2846 -286 2902 -252
rect 2936 -286 2997 -252
rect 2303 -290 2997 -286
rect 2303 -324 2390 -290
rect 2424 -324 2490 -290
rect 2524 -324 2590 -290
rect 2624 -324 2690 -290
rect 2724 -324 2790 -290
rect 2824 -324 2890 -290
rect 2924 -324 2997 -290
rect 2303 -342 2997 -324
rect 2303 -376 2362 -342
rect 2396 -376 2452 -342
rect 2486 -376 2542 -342
rect 2576 -376 2632 -342
rect 2666 -376 2722 -342
rect 2756 -376 2812 -342
rect 2846 -376 2902 -342
rect 2936 -376 2997 -342
rect 2303 -390 2997 -376
rect 2303 -424 2390 -390
rect 2424 -424 2490 -390
rect 2524 -424 2590 -390
rect 2624 -424 2690 -390
rect 2724 -424 2790 -390
rect 2824 -424 2890 -390
rect 2924 -424 2997 -390
rect 2303 -432 2997 -424
rect 2303 -466 2362 -432
rect 2396 -466 2452 -432
rect 2486 -466 2542 -432
rect 2576 -466 2632 -432
rect 2666 -466 2722 -432
rect 2756 -466 2812 -432
rect 2846 -466 2902 -432
rect 2936 -466 2997 -432
rect 2303 -490 2997 -466
rect 2303 -522 2390 -490
rect 2424 -522 2490 -490
rect 2303 -556 2362 -522
rect 2424 -524 2452 -522
rect 2396 -556 2452 -524
rect 2486 -524 2490 -522
rect 2524 -522 2590 -490
rect 2524 -524 2542 -522
rect 2486 -556 2542 -524
rect 2576 -524 2590 -522
rect 2624 -522 2690 -490
rect 2724 -522 2790 -490
rect 2824 -522 2890 -490
rect 2924 -522 2997 -490
rect 2624 -524 2632 -522
rect 2576 -556 2632 -524
rect 2666 -524 2690 -522
rect 2756 -524 2790 -522
rect 2846 -524 2890 -522
rect 2666 -556 2722 -524
rect 2756 -556 2812 -524
rect 2846 -556 2902 -524
rect 2936 -556 2997 -522
rect 2303 -590 2997 -556
rect 2303 -612 2390 -590
rect 2424 -612 2490 -590
rect 2303 -646 2362 -612
rect 2424 -624 2452 -612
rect 2396 -646 2452 -624
rect 2486 -624 2490 -612
rect 2524 -612 2590 -590
rect 2524 -624 2542 -612
rect 2486 -646 2542 -624
rect 2576 -624 2590 -612
rect 2624 -612 2690 -590
rect 2724 -612 2790 -590
rect 2824 -612 2890 -590
rect 2924 -612 2997 -590
rect 2624 -624 2632 -612
rect 2576 -646 2632 -624
rect 2666 -624 2690 -612
rect 2756 -624 2790 -612
rect 2846 -624 2890 -612
rect 2666 -646 2722 -624
rect 2756 -646 2812 -624
rect 2846 -646 2902 -624
rect 2936 -646 2997 -612
rect 2303 -690 2997 -646
rect 2303 -702 2390 -690
rect 2424 -702 2490 -690
rect 2303 -736 2362 -702
rect 2424 -724 2452 -702
rect 2396 -736 2452 -724
rect 2486 -724 2490 -702
rect 2524 -702 2590 -690
rect 2524 -724 2542 -702
rect 2486 -736 2542 -724
rect 2576 -724 2590 -702
rect 2624 -702 2690 -690
rect 2724 -702 2790 -690
rect 2824 -702 2890 -690
rect 2924 -702 2997 -690
rect 2624 -724 2632 -702
rect 2576 -736 2632 -724
rect 2666 -724 2690 -702
rect 2756 -724 2790 -702
rect 2846 -724 2890 -702
rect 2666 -736 2722 -724
rect 2756 -736 2812 -724
rect 2846 -736 2902 -724
rect 2936 -736 2997 -702
rect 2303 -797 2997 -736
rect 3059 -135 3131 -79
rect 3059 -169 3078 -135
rect 3112 -169 3131 -135
rect 3059 -225 3131 -169
rect 3059 -259 3078 -225
rect 3112 -259 3131 -225
rect 3059 -315 3131 -259
rect 3059 -349 3078 -315
rect 3112 -349 3131 -315
rect 3059 -405 3131 -349
rect 3059 -439 3078 -405
rect 3112 -439 3131 -405
rect 3059 -495 3131 -439
rect 3059 -529 3078 -495
rect 3112 -529 3131 -495
rect 3059 -585 3131 -529
rect 3059 -619 3078 -585
rect 3112 -619 3131 -585
rect 3059 -675 3131 -619
rect 3059 -709 3078 -675
rect 3112 -709 3131 -675
rect 3059 -765 3131 -709
rect 2169 -859 2241 -818
rect 3059 -799 3078 -765
rect 3112 -799 3131 -765
rect 3059 -859 3131 -799
rect 2169 -878 3131 -859
rect 2169 -912 2280 -878
rect 2314 -912 2370 -878
rect 2404 -912 2460 -878
rect 2494 -912 2550 -878
rect 2584 -912 2640 -878
rect 2674 -912 2730 -878
rect 2764 -912 2820 -878
rect 2854 -912 2910 -878
rect 2944 -912 3000 -878
rect 3034 -912 3131 -878
rect 2169 -931 3131 -912
rect 3195 -78 3226 -50
rect 3260 -50 3300 -44
rect 3493 149 3589 183
rect 4181 149 4277 183
rect 3493 87 3527 149
rect 3260 -78 3294 -50
rect 3195 -134 3294 -78
rect 3195 -168 3226 -134
rect 3260 -168 3294 -134
rect 3195 -224 3294 -168
rect 3195 -258 3226 -224
rect 3260 -258 3294 -224
rect 3195 -314 3294 -258
rect 3195 -348 3226 -314
rect 3260 -348 3294 -314
rect 3195 -404 3294 -348
rect 3195 -438 3226 -404
rect 3260 -438 3294 -404
rect 3195 -494 3294 -438
rect 3195 -528 3226 -494
rect 3260 -528 3294 -494
rect 3195 -584 3294 -528
rect 3195 -618 3226 -584
rect 3260 -618 3294 -584
rect 3195 -674 3294 -618
rect 3195 -708 3226 -674
rect 3260 -708 3294 -674
rect 3195 -764 3294 -708
rect 3195 -798 3226 -764
rect 3260 -798 3294 -764
rect 3195 -854 3294 -798
rect 3195 -888 3226 -854
rect 3260 -888 3294 -854
rect 1835 -978 1866 -944
rect 1900 -978 2039 -944
rect 2073 -978 2105 -944
rect 1835 -995 2105 -978
rect 3195 -944 3294 -888
rect 3195 -978 3226 -944
rect 3260 -978 3294 -944
rect 3195 -995 3294 -978
rect -714 -1028 3294 -995
rect -714 -1062 -580 -1028
rect -546 -1062 -490 -1028
rect -456 -1062 -400 -1028
rect -366 -1062 -310 -1028
rect -276 -1062 -220 -1028
rect -186 -1062 -130 -1028
rect -96 -1062 -40 -1028
rect -6 -1062 50 -1028
rect 84 -1062 140 -1028
rect 174 -1062 230 -1028
rect 264 -1062 320 -1028
rect 354 -1062 410 -1028
rect 444 -1062 780 -1028
rect 814 -1062 870 -1028
rect 904 -1062 960 -1028
rect 994 -1062 1050 -1028
rect 1084 -1062 1140 -1028
rect 1174 -1062 1230 -1028
rect 1264 -1062 1320 -1028
rect 1354 -1062 1410 -1028
rect 1444 -1062 1500 -1028
rect 1534 -1062 1590 -1028
rect 1624 -1062 1680 -1028
rect 1714 -1062 1770 -1028
rect 1804 -1062 2140 -1028
rect 2174 -1062 2230 -1028
rect 2264 -1062 2320 -1028
rect 2354 -1062 2410 -1028
rect 2444 -1062 2500 -1028
rect 2534 -1062 2590 -1028
rect 2624 -1062 2680 -1028
rect 2714 -1062 2770 -1028
rect 2804 -1062 2860 -1028
rect 2894 -1062 2950 -1028
rect 2984 -1062 3040 -1028
rect 3074 -1062 3130 -1028
rect 3164 -1062 3294 -1028
rect -714 -1094 3294 -1062
rect 570 -1160 650 -1094
rect 1930 -1160 2010 -1094
rect -720 -1201 3300 -1160
rect -720 -1224 -580 -1201
rect -720 -1258 -681 -1224
rect -647 -1235 -580 -1224
rect -546 -1235 -490 -1201
rect -456 -1235 -400 -1201
rect -366 -1235 -310 -1201
rect -276 -1235 -220 -1201
rect -186 -1235 -130 -1201
rect -96 -1235 -40 -1201
rect -6 -1235 50 -1201
rect 84 -1235 140 -1201
rect 174 -1235 230 -1201
rect 264 -1235 320 -1201
rect 354 -1235 410 -1201
rect 444 -1224 780 -1201
rect 444 -1235 506 -1224
rect -647 -1258 506 -1235
rect 540 -1258 679 -1224
rect 713 -1235 780 -1224
rect 814 -1235 870 -1201
rect 904 -1235 960 -1201
rect 994 -1235 1050 -1201
rect 1084 -1235 1140 -1201
rect 1174 -1235 1230 -1201
rect 1264 -1235 1320 -1201
rect 1354 -1235 1410 -1201
rect 1444 -1235 1500 -1201
rect 1534 -1235 1590 -1201
rect 1624 -1235 1680 -1201
rect 1714 -1235 1770 -1201
rect 1804 -1224 2140 -1201
rect 1804 -1235 1866 -1224
rect 713 -1258 1866 -1235
rect 1900 -1258 2039 -1224
rect 2073 -1235 2140 -1224
rect 2174 -1235 2230 -1201
rect 2264 -1235 2320 -1201
rect 2354 -1235 2410 -1201
rect 2444 -1235 2500 -1201
rect 2534 -1235 2590 -1201
rect 2624 -1235 2680 -1201
rect 2714 -1235 2770 -1201
rect 2804 -1235 2860 -1201
rect 2894 -1235 2950 -1201
rect 2984 -1235 3040 -1201
rect 3074 -1235 3130 -1201
rect 3164 -1224 3300 -1201
rect 3164 -1235 3226 -1224
rect 2073 -1258 3226 -1235
rect 3260 -1258 3300 -1224
rect -720 -1314 3300 -1258
rect -720 -1348 -681 -1314
rect -647 -1348 506 -1314
rect 540 -1348 679 -1314
rect 713 -1348 1866 -1314
rect 1900 -1348 2039 -1314
rect 2073 -1348 3226 -1314
rect 3260 -1348 3300 -1314
rect -720 -1382 -474 -1348
rect -440 -1382 -384 -1348
rect -350 -1382 -294 -1348
rect -260 -1382 -204 -1348
rect -170 -1382 -114 -1348
rect -80 -1382 -24 -1348
rect 10 -1382 66 -1348
rect 100 -1382 156 -1348
rect 190 -1382 246 -1348
rect 280 -1382 886 -1348
rect 920 -1382 976 -1348
rect 1010 -1382 1066 -1348
rect 1100 -1382 1156 -1348
rect 1190 -1382 1246 -1348
rect 1280 -1382 1336 -1348
rect 1370 -1382 1426 -1348
rect 1460 -1382 1516 -1348
rect 1550 -1382 1606 -1348
rect 1640 -1382 2246 -1348
rect 2280 -1382 2336 -1348
rect 2370 -1382 2426 -1348
rect 2460 -1382 2516 -1348
rect 2550 -1382 2606 -1348
rect 2640 -1382 2696 -1348
rect 2730 -1382 2786 -1348
rect 2820 -1382 2876 -1348
rect 2910 -1382 2966 -1348
rect 3000 -1382 3300 -1348
rect -720 -1404 3300 -1382
rect -720 -1410 -681 -1404
rect -1310 -2233 -1230 -2220
rect -1077 -2233 -1043 -2171
rect -1827 -2267 -1731 -2233
rect -1139 -2267 -1043 -2233
rect -714 -1438 -681 -1410
rect -647 -1405 506 -1404
rect -647 -1410 358 -1405
rect -647 -1438 -615 -1410
rect -714 -1494 -615 -1438
rect -714 -1528 -681 -1494
rect -647 -1528 -615 -1494
rect -714 -1584 -615 -1528
rect -714 -1618 -681 -1584
rect -647 -1618 -615 -1584
rect -714 -1674 -615 -1618
rect -714 -1708 -681 -1674
rect -647 -1708 -615 -1674
rect -714 -1764 -615 -1708
rect -714 -1798 -681 -1764
rect -647 -1798 -615 -1764
rect -714 -1854 -615 -1798
rect -714 -1888 -681 -1854
rect -647 -1888 -615 -1854
rect -714 -1944 -615 -1888
rect -714 -1978 -681 -1944
rect -647 -1978 -615 -1944
rect -714 -2034 -615 -1978
rect -714 -2068 -681 -2034
rect -647 -2068 -615 -2034
rect -714 -2124 -615 -2068
rect -714 -2158 -681 -2124
rect -647 -2158 -615 -2124
rect -714 -2214 -615 -2158
rect -714 -2248 -681 -2214
rect -647 -2248 -615 -2214
rect -3540 -2300 -3460 -2280
rect -2750 -2280 -2730 -2270
rect -2690 -2280 -2670 -2270
rect -2750 -2300 -2670 -2280
rect -1310 -2280 -1290 -2267
rect -1250 -2280 -1230 -2267
rect -1310 -2300 -1230 -2280
rect -714 -2304 -615 -2248
rect -551 -1424 -479 -1410
rect -551 -1458 -532 -1424
rect -498 -1458 -479 -1424
rect -551 -1514 -479 -1458
rect 339 -1439 358 -1410
rect 392 -1410 506 -1405
rect 392 -1439 411 -1410
rect -551 -1548 -532 -1514
rect -498 -1548 -479 -1514
rect -551 -1604 -479 -1548
rect -551 -1638 -532 -1604
rect -498 -1638 -479 -1604
rect -551 -1694 -479 -1638
rect -551 -1728 -532 -1694
rect -498 -1728 -479 -1694
rect -551 -1784 -479 -1728
rect -551 -1818 -532 -1784
rect -498 -1818 -479 -1784
rect -551 -1874 -479 -1818
rect -551 -1908 -532 -1874
rect -498 -1908 -479 -1874
rect -551 -1964 -479 -1908
rect -551 -1998 -532 -1964
rect -498 -1998 -479 -1964
rect -551 -2054 -479 -1998
rect -551 -2088 -532 -2054
rect -498 -2088 -479 -2054
rect -551 -2144 -479 -2088
rect -551 -2178 -532 -2144
rect -498 -2178 -479 -2144
rect -417 -1522 277 -1463
rect -417 -1556 -358 -1522
rect -324 -1550 -268 -1522
rect -296 -1556 -268 -1550
rect -234 -1550 -178 -1522
rect -234 -1556 -230 -1550
rect -417 -1584 -330 -1556
rect -296 -1584 -230 -1556
rect -196 -1556 -178 -1550
rect -144 -1550 -88 -1522
rect -144 -1556 -130 -1550
rect -196 -1584 -130 -1556
rect -96 -1556 -88 -1550
rect -54 -1550 2 -1522
rect 36 -1550 92 -1522
rect 126 -1550 182 -1522
rect -54 -1556 -30 -1550
rect 36 -1556 70 -1550
rect 126 -1556 170 -1550
rect 216 -1556 277 -1522
rect -96 -1584 -30 -1556
rect 4 -1584 70 -1556
rect 104 -1584 170 -1556
rect 204 -1584 277 -1556
rect -417 -1612 277 -1584
rect -417 -1646 -358 -1612
rect -324 -1646 -268 -1612
rect -234 -1646 -178 -1612
rect -144 -1646 -88 -1612
rect -54 -1646 2 -1612
rect 36 -1646 92 -1612
rect 126 -1646 182 -1612
rect 216 -1646 277 -1612
rect -417 -1650 277 -1646
rect -417 -1684 -330 -1650
rect -296 -1684 -230 -1650
rect -196 -1684 -130 -1650
rect -96 -1684 -30 -1650
rect 4 -1684 70 -1650
rect 104 -1684 170 -1650
rect 204 -1684 277 -1650
rect -417 -1702 277 -1684
rect -417 -1736 -358 -1702
rect -324 -1736 -268 -1702
rect -234 -1736 -178 -1702
rect -144 -1736 -88 -1702
rect -54 -1736 2 -1702
rect 36 -1736 92 -1702
rect 126 -1736 182 -1702
rect 216 -1736 277 -1702
rect -417 -1750 277 -1736
rect -417 -1784 -330 -1750
rect -296 -1784 -230 -1750
rect -196 -1784 -130 -1750
rect -96 -1784 -30 -1750
rect 4 -1784 70 -1750
rect 104 -1784 170 -1750
rect 204 -1784 277 -1750
rect -417 -1792 277 -1784
rect -417 -1826 -358 -1792
rect -324 -1826 -268 -1792
rect -234 -1826 -178 -1792
rect -144 -1826 -88 -1792
rect -54 -1826 2 -1792
rect 36 -1826 92 -1792
rect 126 -1826 182 -1792
rect 216 -1826 277 -1792
rect -417 -1850 277 -1826
rect -417 -1882 -330 -1850
rect -296 -1882 -230 -1850
rect -417 -1916 -358 -1882
rect -296 -1884 -268 -1882
rect -324 -1916 -268 -1884
rect -234 -1884 -230 -1882
rect -196 -1882 -130 -1850
rect -196 -1884 -178 -1882
rect -234 -1916 -178 -1884
rect -144 -1884 -130 -1882
rect -96 -1882 -30 -1850
rect 4 -1882 70 -1850
rect 104 -1882 170 -1850
rect 204 -1882 277 -1850
rect -96 -1884 -88 -1882
rect -144 -1916 -88 -1884
rect -54 -1884 -30 -1882
rect 36 -1884 70 -1882
rect 126 -1884 170 -1882
rect -54 -1916 2 -1884
rect 36 -1916 92 -1884
rect 126 -1916 182 -1884
rect 216 -1916 277 -1882
rect -417 -1950 277 -1916
rect -417 -1972 -330 -1950
rect -296 -1972 -230 -1950
rect -417 -2006 -358 -1972
rect -296 -1984 -268 -1972
rect -324 -2006 -268 -1984
rect -234 -1984 -230 -1972
rect -196 -1972 -130 -1950
rect -196 -1984 -178 -1972
rect -234 -2006 -178 -1984
rect -144 -1984 -130 -1972
rect -96 -1972 -30 -1950
rect 4 -1972 70 -1950
rect 104 -1972 170 -1950
rect 204 -1972 277 -1950
rect -96 -1984 -88 -1972
rect -144 -2006 -88 -1984
rect -54 -1984 -30 -1972
rect 36 -1984 70 -1972
rect 126 -1984 170 -1972
rect -54 -2006 2 -1984
rect 36 -2006 92 -1984
rect 126 -2006 182 -1984
rect 216 -2006 277 -1972
rect -417 -2050 277 -2006
rect -417 -2062 -330 -2050
rect -296 -2062 -230 -2050
rect -417 -2096 -358 -2062
rect -296 -2084 -268 -2062
rect -324 -2096 -268 -2084
rect -234 -2084 -230 -2062
rect -196 -2062 -130 -2050
rect -196 -2084 -178 -2062
rect -234 -2096 -178 -2084
rect -144 -2084 -130 -2062
rect -96 -2062 -30 -2050
rect 4 -2062 70 -2050
rect 104 -2062 170 -2050
rect 204 -2062 277 -2050
rect -96 -2084 -88 -2062
rect -144 -2096 -88 -2084
rect -54 -2084 -30 -2062
rect 36 -2084 70 -2062
rect 126 -2084 170 -2062
rect -54 -2096 2 -2084
rect 36 -2096 92 -2084
rect 126 -2096 182 -2084
rect 216 -2096 277 -2062
rect -417 -2157 277 -2096
rect 339 -1495 411 -1439
rect 339 -1529 358 -1495
rect 392 -1529 411 -1495
rect 339 -1585 411 -1529
rect 339 -1619 358 -1585
rect 392 -1619 411 -1585
rect 339 -1675 411 -1619
rect 339 -1709 358 -1675
rect 392 -1709 411 -1675
rect 339 -1765 411 -1709
rect 339 -1799 358 -1765
rect 392 -1799 411 -1765
rect 339 -1855 411 -1799
rect 339 -1889 358 -1855
rect 392 -1889 411 -1855
rect 339 -1945 411 -1889
rect 339 -1979 358 -1945
rect 392 -1979 411 -1945
rect 339 -2035 411 -1979
rect 339 -2069 358 -2035
rect 392 -2069 411 -2035
rect 339 -2125 411 -2069
rect -551 -2219 -479 -2178
rect 339 -2159 358 -2125
rect 392 -2159 411 -2125
rect 339 -2219 411 -2159
rect -551 -2238 411 -2219
rect -551 -2272 -440 -2238
rect -406 -2272 -350 -2238
rect -316 -2272 -260 -2238
rect -226 -2272 -170 -2238
rect -136 -2272 -80 -2238
rect -46 -2272 10 -2238
rect 44 -2272 100 -2238
rect 134 -2272 190 -2238
rect 224 -2272 280 -2238
rect 314 -2272 411 -2238
rect -551 -2291 411 -2272
rect 475 -1438 506 -1410
rect 540 -1438 679 -1404
rect 713 -1405 1866 -1404
rect 713 -1410 1718 -1405
rect 713 -1438 745 -1410
rect 475 -1494 745 -1438
rect 475 -1528 506 -1494
rect 540 -1528 679 -1494
rect 713 -1528 745 -1494
rect 475 -1584 745 -1528
rect 475 -1618 506 -1584
rect 540 -1618 679 -1584
rect 713 -1618 745 -1584
rect 475 -1674 745 -1618
rect 475 -1708 506 -1674
rect 540 -1708 679 -1674
rect 713 -1708 745 -1674
rect 475 -1764 745 -1708
rect 475 -1798 506 -1764
rect 540 -1798 679 -1764
rect 713 -1798 745 -1764
rect 475 -1854 745 -1798
rect 475 -1888 506 -1854
rect 540 -1888 679 -1854
rect 713 -1888 745 -1854
rect 475 -1944 745 -1888
rect 475 -1978 506 -1944
rect 540 -1978 679 -1944
rect 713 -1978 745 -1944
rect 475 -2034 745 -1978
rect 475 -2068 506 -2034
rect 540 -2068 679 -2034
rect 713 -2068 745 -2034
rect 475 -2124 745 -2068
rect 475 -2158 506 -2124
rect 540 -2158 679 -2124
rect 713 -2158 745 -2124
rect 475 -2214 745 -2158
rect 475 -2248 506 -2214
rect 540 -2248 679 -2214
rect 713 -2248 745 -2214
rect -714 -2338 -681 -2304
rect -647 -2338 -615 -2304
rect -714 -2355 -615 -2338
rect 475 -2304 745 -2248
rect 809 -1424 881 -1410
rect 809 -1458 828 -1424
rect 862 -1458 881 -1424
rect 809 -1514 881 -1458
rect 1699 -1439 1718 -1410
rect 1752 -1410 1866 -1405
rect 1752 -1439 1771 -1410
rect 809 -1548 828 -1514
rect 862 -1548 881 -1514
rect 809 -1604 881 -1548
rect 809 -1638 828 -1604
rect 862 -1638 881 -1604
rect 809 -1694 881 -1638
rect 809 -1728 828 -1694
rect 862 -1728 881 -1694
rect 809 -1784 881 -1728
rect 809 -1818 828 -1784
rect 862 -1818 881 -1784
rect 809 -1874 881 -1818
rect 809 -1908 828 -1874
rect 862 -1908 881 -1874
rect 809 -1964 881 -1908
rect 809 -1998 828 -1964
rect 862 -1998 881 -1964
rect 809 -2054 881 -1998
rect 809 -2088 828 -2054
rect 862 -2088 881 -2054
rect 809 -2144 881 -2088
rect 809 -2178 828 -2144
rect 862 -2178 881 -2144
rect 943 -1522 1637 -1463
rect 943 -1556 1002 -1522
rect 1036 -1550 1092 -1522
rect 1064 -1556 1092 -1550
rect 1126 -1550 1182 -1522
rect 1126 -1556 1130 -1550
rect 943 -1584 1030 -1556
rect 1064 -1584 1130 -1556
rect 1164 -1556 1182 -1550
rect 1216 -1550 1272 -1522
rect 1216 -1556 1230 -1550
rect 1164 -1584 1230 -1556
rect 1264 -1556 1272 -1550
rect 1306 -1550 1362 -1522
rect 1396 -1550 1452 -1522
rect 1486 -1550 1542 -1522
rect 1306 -1556 1330 -1550
rect 1396 -1556 1430 -1550
rect 1486 -1556 1530 -1550
rect 1576 -1556 1637 -1522
rect 1264 -1584 1330 -1556
rect 1364 -1584 1430 -1556
rect 1464 -1584 1530 -1556
rect 1564 -1584 1637 -1556
rect 943 -1612 1637 -1584
rect 943 -1646 1002 -1612
rect 1036 -1646 1092 -1612
rect 1126 -1646 1182 -1612
rect 1216 -1646 1272 -1612
rect 1306 -1646 1362 -1612
rect 1396 -1646 1452 -1612
rect 1486 -1646 1542 -1612
rect 1576 -1646 1637 -1612
rect 943 -1650 1637 -1646
rect 943 -1684 1030 -1650
rect 1064 -1684 1130 -1650
rect 1164 -1684 1230 -1650
rect 1264 -1684 1330 -1650
rect 1364 -1684 1430 -1650
rect 1464 -1684 1530 -1650
rect 1564 -1684 1637 -1650
rect 943 -1702 1637 -1684
rect 943 -1736 1002 -1702
rect 1036 -1736 1092 -1702
rect 1126 -1736 1182 -1702
rect 1216 -1736 1272 -1702
rect 1306 -1736 1362 -1702
rect 1396 -1736 1452 -1702
rect 1486 -1736 1542 -1702
rect 1576 -1736 1637 -1702
rect 943 -1750 1637 -1736
rect 943 -1784 1030 -1750
rect 1064 -1784 1130 -1750
rect 1164 -1784 1230 -1750
rect 1264 -1784 1330 -1750
rect 1364 -1784 1430 -1750
rect 1464 -1784 1530 -1750
rect 1564 -1784 1637 -1750
rect 943 -1792 1637 -1784
rect 943 -1826 1002 -1792
rect 1036 -1826 1092 -1792
rect 1126 -1826 1182 -1792
rect 1216 -1826 1272 -1792
rect 1306 -1826 1362 -1792
rect 1396 -1826 1452 -1792
rect 1486 -1826 1542 -1792
rect 1576 -1826 1637 -1792
rect 943 -1850 1637 -1826
rect 943 -1882 1030 -1850
rect 1064 -1882 1130 -1850
rect 943 -1916 1002 -1882
rect 1064 -1884 1092 -1882
rect 1036 -1916 1092 -1884
rect 1126 -1884 1130 -1882
rect 1164 -1882 1230 -1850
rect 1164 -1884 1182 -1882
rect 1126 -1916 1182 -1884
rect 1216 -1884 1230 -1882
rect 1264 -1882 1330 -1850
rect 1364 -1882 1430 -1850
rect 1464 -1882 1530 -1850
rect 1564 -1882 1637 -1850
rect 1264 -1884 1272 -1882
rect 1216 -1916 1272 -1884
rect 1306 -1884 1330 -1882
rect 1396 -1884 1430 -1882
rect 1486 -1884 1530 -1882
rect 1306 -1916 1362 -1884
rect 1396 -1916 1452 -1884
rect 1486 -1916 1542 -1884
rect 1576 -1916 1637 -1882
rect 943 -1950 1637 -1916
rect 943 -1972 1030 -1950
rect 1064 -1972 1130 -1950
rect 943 -2006 1002 -1972
rect 1064 -1984 1092 -1972
rect 1036 -2006 1092 -1984
rect 1126 -1984 1130 -1972
rect 1164 -1972 1230 -1950
rect 1164 -1984 1182 -1972
rect 1126 -2006 1182 -1984
rect 1216 -1984 1230 -1972
rect 1264 -1972 1330 -1950
rect 1364 -1972 1430 -1950
rect 1464 -1972 1530 -1950
rect 1564 -1972 1637 -1950
rect 1264 -1984 1272 -1972
rect 1216 -2006 1272 -1984
rect 1306 -1984 1330 -1972
rect 1396 -1984 1430 -1972
rect 1486 -1984 1530 -1972
rect 1306 -2006 1362 -1984
rect 1396 -2006 1452 -1984
rect 1486 -2006 1542 -1984
rect 1576 -2006 1637 -1972
rect 943 -2050 1637 -2006
rect 943 -2062 1030 -2050
rect 1064 -2062 1130 -2050
rect 943 -2096 1002 -2062
rect 1064 -2084 1092 -2062
rect 1036 -2096 1092 -2084
rect 1126 -2084 1130 -2062
rect 1164 -2062 1230 -2050
rect 1164 -2084 1182 -2062
rect 1126 -2096 1182 -2084
rect 1216 -2084 1230 -2062
rect 1264 -2062 1330 -2050
rect 1364 -2062 1430 -2050
rect 1464 -2062 1530 -2050
rect 1564 -2062 1637 -2050
rect 1264 -2084 1272 -2062
rect 1216 -2096 1272 -2084
rect 1306 -2084 1330 -2062
rect 1396 -2084 1430 -2062
rect 1486 -2084 1530 -2062
rect 1306 -2096 1362 -2084
rect 1396 -2096 1452 -2084
rect 1486 -2096 1542 -2084
rect 1576 -2096 1637 -2062
rect 943 -2157 1637 -2096
rect 1699 -1495 1771 -1439
rect 1699 -1529 1718 -1495
rect 1752 -1529 1771 -1495
rect 1699 -1585 1771 -1529
rect 1699 -1619 1718 -1585
rect 1752 -1619 1771 -1585
rect 1699 -1675 1771 -1619
rect 1699 -1709 1718 -1675
rect 1752 -1709 1771 -1675
rect 1699 -1765 1771 -1709
rect 1699 -1799 1718 -1765
rect 1752 -1799 1771 -1765
rect 1699 -1855 1771 -1799
rect 1699 -1889 1718 -1855
rect 1752 -1889 1771 -1855
rect 1699 -1945 1771 -1889
rect 1699 -1979 1718 -1945
rect 1752 -1979 1771 -1945
rect 1699 -2035 1771 -1979
rect 1699 -2069 1718 -2035
rect 1752 -2069 1771 -2035
rect 1699 -2125 1771 -2069
rect 809 -2219 881 -2178
rect 1699 -2159 1718 -2125
rect 1752 -2159 1771 -2125
rect 1699 -2219 1771 -2159
rect 809 -2238 1771 -2219
rect 809 -2272 920 -2238
rect 954 -2272 1010 -2238
rect 1044 -2272 1100 -2238
rect 1134 -2272 1190 -2238
rect 1224 -2272 1280 -2238
rect 1314 -2272 1370 -2238
rect 1404 -2272 1460 -2238
rect 1494 -2272 1550 -2238
rect 1584 -2272 1640 -2238
rect 1674 -2272 1771 -2238
rect 809 -2291 1771 -2272
rect 1835 -1438 1866 -1410
rect 1900 -1438 2039 -1404
rect 2073 -1405 3226 -1404
rect 2073 -1410 3078 -1405
rect 2073 -1438 2105 -1410
rect 1835 -1494 2105 -1438
rect 1835 -1528 1866 -1494
rect 1900 -1528 2039 -1494
rect 2073 -1528 2105 -1494
rect 1835 -1584 2105 -1528
rect 1835 -1618 1866 -1584
rect 1900 -1618 2039 -1584
rect 2073 -1618 2105 -1584
rect 1835 -1674 2105 -1618
rect 1835 -1708 1866 -1674
rect 1900 -1708 2039 -1674
rect 2073 -1708 2105 -1674
rect 1835 -1764 2105 -1708
rect 1835 -1798 1866 -1764
rect 1900 -1798 2039 -1764
rect 2073 -1798 2105 -1764
rect 1835 -1854 2105 -1798
rect 1835 -1888 1866 -1854
rect 1900 -1888 2039 -1854
rect 2073 -1888 2105 -1854
rect 1835 -1944 2105 -1888
rect 1835 -1978 1866 -1944
rect 1900 -1978 2039 -1944
rect 2073 -1978 2105 -1944
rect 1835 -2034 2105 -1978
rect 1835 -2068 1866 -2034
rect 1900 -2068 2039 -2034
rect 2073 -2068 2105 -2034
rect 1835 -2124 2105 -2068
rect 1835 -2158 1866 -2124
rect 1900 -2158 2039 -2124
rect 2073 -2158 2105 -2124
rect 1835 -2214 2105 -2158
rect 1835 -2248 1866 -2214
rect 1900 -2248 2039 -2214
rect 2073 -2248 2105 -2214
rect 475 -2338 506 -2304
rect 540 -2338 679 -2304
rect 713 -2338 745 -2304
rect 475 -2355 745 -2338
rect 1835 -2304 2105 -2248
rect 2169 -1424 2241 -1410
rect 2169 -1458 2188 -1424
rect 2222 -1458 2241 -1424
rect 2169 -1514 2241 -1458
rect 3059 -1439 3078 -1410
rect 3112 -1410 3226 -1405
rect 3112 -1439 3131 -1410
rect 2169 -1548 2188 -1514
rect 2222 -1548 2241 -1514
rect 2169 -1604 2241 -1548
rect 2169 -1638 2188 -1604
rect 2222 -1638 2241 -1604
rect 2169 -1694 2241 -1638
rect 2169 -1728 2188 -1694
rect 2222 -1728 2241 -1694
rect 2169 -1784 2241 -1728
rect 2169 -1818 2188 -1784
rect 2222 -1818 2241 -1784
rect 2169 -1874 2241 -1818
rect 2169 -1908 2188 -1874
rect 2222 -1908 2241 -1874
rect 2169 -1964 2241 -1908
rect 2169 -1998 2188 -1964
rect 2222 -1998 2241 -1964
rect 2169 -2054 2241 -1998
rect 2169 -2088 2188 -2054
rect 2222 -2088 2241 -2054
rect 2169 -2144 2241 -2088
rect 2169 -2178 2188 -2144
rect 2222 -2178 2241 -2144
rect 2303 -1522 2997 -1463
rect 2303 -1556 2362 -1522
rect 2396 -1550 2452 -1522
rect 2424 -1556 2452 -1550
rect 2486 -1550 2542 -1522
rect 2486 -1556 2490 -1550
rect 2303 -1584 2390 -1556
rect 2424 -1584 2490 -1556
rect 2524 -1556 2542 -1550
rect 2576 -1550 2632 -1522
rect 2576 -1556 2590 -1550
rect 2524 -1584 2590 -1556
rect 2624 -1556 2632 -1550
rect 2666 -1550 2722 -1522
rect 2756 -1550 2812 -1522
rect 2846 -1550 2902 -1522
rect 2666 -1556 2690 -1550
rect 2756 -1556 2790 -1550
rect 2846 -1556 2890 -1550
rect 2936 -1556 2997 -1522
rect 2624 -1584 2690 -1556
rect 2724 -1584 2790 -1556
rect 2824 -1584 2890 -1556
rect 2924 -1584 2997 -1556
rect 2303 -1612 2997 -1584
rect 2303 -1646 2362 -1612
rect 2396 -1646 2452 -1612
rect 2486 -1646 2542 -1612
rect 2576 -1646 2632 -1612
rect 2666 -1646 2722 -1612
rect 2756 -1646 2812 -1612
rect 2846 -1646 2902 -1612
rect 2936 -1646 2997 -1612
rect 2303 -1650 2997 -1646
rect 2303 -1684 2390 -1650
rect 2424 -1684 2490 -1650
rect 2524 -1684 2590 -1650
rect 2624 -1684 2690 -1650
rect 2724 -1684 2790 -1650
rect 2824 -1684 2890 -1650
rect 2924 -1684 2997 -1650
rect 2303 -1702 2997 -1684
rect 2303 -1736 2362 -1702
rect 2396 -1736 2452 -1702
rect 2486 -1736 2542 -1702
rect 2576 -1736 2632 -1702
rect 2666 -1736 2722 -1702
rect 2756 -1736 2812 -1702
rect 2846 -1736 2902 -1702
rect 2936 -1736 2997 -1702
rect 2303 -1750 2997 -1736
rect 2303 -1784 2390 -1750
rect 2424 -1784 2490 -1750
rect 2524 -1784 2590 -1750
rect 2624 -1784 2690 -1750
rect 2724 -1784 2790 -1750
rect 2824 -1784 2890 -1750
rect 2924 -1784 2997 -1750
rect 2303 -1792 2997 -1784
rect 2303 -1826 2362 -1792
rect 2396 -1826 2452 -1792
rect 2486 -1826 2542 -1792
rect 2576 -1826 2632 -1792
rect 2666 -1826 2722 -1792
rect 2756 -1826 2812 -1792
rect 2846 -1826 2902 -1792
rect 2936 -1826 2997 -1792
rect 2303 -1850 2997 -1826
rect 2303 -1882 2390 -1850
rect 2424 -1882 2490 -1850
rect 2303 -1916 2362 -1882
rect 2424 -1884 2452 -1882
rect 2396 -1916 2452 -1884
rect 2486 -1884 2490 -1882
rect 2524 -1882 2590 -1850
rect 2524 -1884 2542 -1882
rect 2486 -1916 2542 -1884
rect 2576 -1884 2590 -1882
rect 2624 -1882 2690 -1850
rect 2724 -1882 2790 -1850
rect 2824 -1882 2890 -1850
rect 2924 -1882 2997 -1850
rect 2624 -1884 2632 -1882
rect 2576 -1916 2632 -1884
rect 2666 -1884 2690 -1882
rect 2756 -1884 2790 -1882
rect 2846 -1884 2890 -1882
rect 2666 -1916 2722 -1884
rect 2756 -1916 2812 -1884
rect 2846 -1916 2902 -1884
rect 2936 -1916 2997 -1882
rect 2303 -1950 2997 -1916
rect 2303 -1972 2390 -1950
rect 2424 -1972 2490 -1950
rect 2303 -2006 2362 -1972
rect 2424 -1984 2452 -1972
rect 2396 -2006 2452 -1984
rect 2486 -1984 2490 -1972
rect 2524 -1972 2590 -1950
rect 2524 -1984 2542 -1972
rect 2486 -2006 2542 -1984
rect 2576 -1984 2590 -1972
rect 2624 -1972 2690 -1950
rect 2724 -1972 2790 -1950
rect 2824 -1972 2890 -1950
rect 2924 -1972 2997 -1950
rect 2624 -1984 2632 -1972
rect 2576 -2006 2632 -1984
rect 2666 -1984 2690 -1972
rect 2756 -1984 2790 -1972
rect 2846 -1984 2890 -1972
rect 2666 -2006 2722 -1984
rect 2756 -2006 2812 -1984
rect 2846 -2006 2902 -1984
rect 2936 -2006 2997 -1972
rect 2303 -2050 2997 -2006
rect 2303 -2062 2390 -2050
rect 2424 -2062 2490 -2050
rect 2303 -2096 2362 -2062
rect 2424 -2084 2452 -2062
rect 2396 -2096 2452 -2084
rect 2486 -2084 2490 -2062
rect 2524 -2062 2590 -2050
rect 2524 -2084 2542 -2062
rect 2486 -2096 2542 -2084
rect 2576 -2084 2590 -2062
rect 2624 -2062 2690 -2050
rect 2724 -2062 2790 -2050
rect 2824 -2062 2890 -2050
rect 2924 -2062 2997 -2050
rect 2624 -2084 2632 -2062
rect 2576 -2096 2632 -2084
rect 2666 -2084 2690 -2062
rect 2756 -2084 2790 -2062
rect 2846 -2084 2890 -2062
rect 2666 -2096 2722 -2084
rect 2756 -2096 2812 -2084
rect 2846 -2096 2902 -2084
rect 2936 -2096 2997 -2062
rect 2303 -2157 2997 -2096
rect 3059 -1495 3131 -1439
rect 3059 -1529 3078 -1495
rect 3112 -1529 3131 -1495
rect 3059 -1585 3131 -1529
rect 3059 -1619 3078 -1585
rect 3112 -1619 3131 -1585
rect 3059 -1675 3131 -1619
rect 3059 -1709 3078 -1675
rect 3112 -1709 3131 -1675
rect 3059 -1765 3131 -1709
rect 3059 -1799 3078 -1765
rect 3112 -1799 3131 -1765
rect 3059 -1855 3131 -1799
rect 3059 -1889 3078 -1855
rect 3112 -1889 3131 -1855
rect 3059 -1945 3131 -1889
rect 3059 -1979 3078 -1945
rect 3112 -1979 3131 -1945
rect 3059 -2035 3131 -1979
rect 3059 -2069 3078 -2035
rect 3112 -2069 3131 -2035
rect 3059 -2125 3131 -2069
rect 2169 -2219 2241 -2178
rect 3059 -2159 3078 -2125
rect 3112 -2159 3131 -2125
rect 3059 -2219 3131 -2159
rect 2169 -2238 3131 -2219
rect 2169 -2272 2280 -2238
rect 2314 -2272 2370 -2238
rect 2404 -2272 2460 -2238
rect 2494 -2272 2550 -2238
rect 2584 -2272 2640 -2238
rect 2674 -2272 2730 -2238
rect 2764 -2272 2820 -2238
rect 2854 -2272 2910 -2238
rect 2944 -2272 3000 -2238
rect 3034 -2272 3131 -2238
rect 2169 -2291 3131 -2272
rect 3195 -1438 3226 -1410
rect 3260 -1410 3300 -1404
rect 3260 -1438 3294 -1410
rect 3195 -1494 3294 -1438
rect 3195 -1528 3226 -1494
rect 3260 -1528 3294 -1494
rect 3195 -1584 3294 -1528
rect 3195 -1618 3226 -1584
rect 3260 -1618 3294 -1584
rect 3195 -1674 3294 -1618
rect 3195 -1708 3226 -1674
rect 3260 -1708 3294 -1674
rect 3195 -1764 3294 -1708
rect 3195 -1798 3226 -1764
rect 3260 -1798 3294 -1764
rect 3195 -1854 3294 -1798
rect 3195 -1888 3226 -1854
rect 3260 -1888 3294 -1854
rect 3195 -1944 3294 -1888
rect 3195 -1978 3226 -1944
rect 3260 -1978 3294 -1944
rect 3195 -2034 3294 -1978
rect 3195 -2068 3226 -2034
rect 3260 -2068 3294 -2034
rect 3195 -2124 3294 -2068
rect 3195 -2158 3226 -2124
rect 3260 -2158 3294 -2124
rect 3195 -2214 3294 -2158
rect 3195 -2248 3226 -2214
rect 3260 -2248 3294 -2214
rect 1835 -2338 1866 -2304
rect 1900 -2338 2039 -2304
rect 2073 -2338 2105 -2304
rect 1835 -2355 2105 -2338
rect 3195 -2304 3294 -2248
rect 4243 87 4277 149
rect 3493 -2233 3527 -2171
rect 5393 -781 5489 -747
rect 5749 -781 5845 -747
rect 5393 -843 5427 -781
rect 3680 -2233 3760 -2220
rect 4243 -2233 4277 -2171
rect 3493 -2267 3589 -2233
rect 4181 -2267 4277 -2233
rect 4606 -988 4702 -954
rect 4962 -988 5058 -954
rect 4606 -1050 4640 -988
rect 5024 -1050 5058 -988
rect 4606 -2230 4640 -2168
rect 4790 -2230 4870 -2220
rect 5024 -2230 5058 -2168
rect 4606 -2264 4702 -2230
rect 4962 -2264 5058 -2230
rect 5811 -843 5845 -781
rect 5393 -2233 5427 -2171
rect 5580 -2233 5660 -2220
rect 5811 -2233 5845 -2171
rect 3680 -2280 3700 -2267
rect 3740 -2280 3760 -2267
rect 3680 -2300 3760 -2280
rect 4790 -2280 4810 -2264
rect 4850 -2280 4870 -2264
rect 5393 -2267 5489 -2233
rect 5749 -2267 5845 -2233
rect 4790 -2300 4870 -2280
rect 5580 -2280 5600 -2267
rect 5640 -2280 5660 -2267
rect 5580 -2300 5660 -2280
rect 3195 -2338 3226 -2304
rect 3260 -2338 3294 -2304
rect 3195 -2355 3294 -2338
rect -714 -2388 3294 -2355
rect -714 -2422 -580 -2388
rect -546 -2422 -490 -2388
rect -456 -2422 -400 -2388
rect -366 -2422 -310 -2388
rect -276 -2422 -220 -2388
rect -186 -2422 -130 -2388
rect -96 -2422 -40 -2388
rect -6 -2422 50 -2388
rect 84 -2422 140 -2388
rect 174 -2422 230 -2388
rect 264 -2422 320 -2388
rect 354 -2422 410 -2388
rect 444 -2422 780 -2388
rect 814 -2422 870 -2388
rect 904 -2422 960 -2388
rect 994 -2422 1050 -2388
rect 1084 -2422 1140 -2388
rect 1174 -2422 1230 -2388
rect 1264 -2422 1320 -2388
rect 1354 -2422 1410 -2388
rect 1444 -2422 1500 -2388
rect 1534 -2422 1590 -2388
rect 1624 -2422 1680 -2388
rect 1714 -2422 1770 -2388
rect 1804 -2422 2140 -2388
rect 2174 -2422 2230 -2388
rect 2264 -2422 2320 -2388
rect 2354 -2422 2410 -2388
rect 2444 -2422 2500 -2388
rect 2534 -2422 2590 -2388
rect 2624 -2422 2680 -2388
rect 2714 -2422 2770 -2388
rect 2804 -2422 2860 -2388
rect 2894 -2422 2950 -2388
rect 2984 -2422 3040 -2388
rect 3074 -2422 3130 -2388
rect 3164 -2422 3294 -2388
rect -714 -2454 3294 -2422
rect 570 -2460 650 -2454
rect 1250 -2540 1330 -2454
rect 1930 -2460 2010 -2454
rect 1250 -2580 1270 -2540
rect 1310 -2580 1330 -2540
rect 1250 -2620 1330 -2580
rect 1250 -2660 1270 -2620
rect 1310 -2660 1330 -2620
rect 1250 -2700 1330 -2660
rect 1250 -2740 1270 -2700
rect 1310 -2740 1330 -2700
rect 1250 -2760 1330 -2740
rect 2863 -2949 2959 -2915
rect 5381 -2949 5477 -2915
rect 2863 -3011 2897 -2949
rect 5443 -3011 5477 -2949
rect 2863 -3333 2897 -3271
rect 4130 -3310 4210 -3290
rect 4130 -3333 4150 -3310
rect 4190 -3333 4210 -3310
rect 5443 -3333 5477 -3271
rect 2863 -3367 2959 -3333
rect 5381 -3367 5477 -3333
rect 4130 -3370 4210 -3367
<< viali >>
rect 11340 14410 11380 14450
rect 11860 14410 11900 14450
rect 12380 14410 12420 14450
rect 12870 14410 12910 14450
rect 11230 14280 11270 14320
rect 11230 14180 11270 14220
rect 11340 14280 11380 14320
rect 11340 14180 11380 14220
rect 11750 14280 11790 14320
rect 11750 14180 11790 14220
rect 11860 14280 11900 14320
rect 11860 14180 11900 14220
rect 12270 14280 12310 14320
rect 12270 14180 12310 14220
rect 12380 14280 12420 14320
rect 12380 14180 12420 14220
rect 12870 14280 12910 14320
rect 12870 14180 12910 14220
rect 12980 14280 13020 14320
rect 12980 14180 13020 14220
rect 11288 14068 11322 14102
rect 11808 14068 11842 14102
rect 12328 14068 12362 14102
rect 12896 14068 12930 14102
rect 11230 13900 11270 13940
rect 11230 13800 11270 13840
rect 11230 13700 11270 13740
rect 11340 13900 11380 13940
rect 11340 13800 11380 13840
rect 11340 13700 11380 13740
rect 11750 13900 11790 13940
rect 11750 13800 11790 13840
rect 11750 13700 11790 13740
rect 11860 13900 11900 13940
rect 11860 13800 11900 13840
rect 11860 13700 11900 13740
rect 12270 13900 12310 13940
rect 12270 13800 12310 13840
rect 12270 13700 12310 13740
rect 12380 13900 12420 13940
rect 12380 13800 12420 13840
rect 12380 13700 12420 13740
rect 570 13380 610 13420
rect 790 13380 830 13420
rect 1260 13380 1300 13420
rect 1600 13380 1640 13420
rect 1820 13380 1860 13420
rect 2260 13380 2300 13420
rect 2940 13380 2980 13420
rect 3160 13380 3200 13420
rect 3630 13380 3670 13420
rect 4090 13380 4130 13420
rect 4440 13380 4480 13420
rect 4690 13380 4730 13420
rect 4910 13380 4950 13420
rect 5240 13380 5280 13420
rect 5900 13380 5940 13420
rect 6120 13380 6160 13420
rect 6690 13380 6730 13420
rect 6950 13380 6990 13420
rect 7200 13380 7240 13420
rect 7420 13380 7460 13420
rect 7970 13380 8010 13420
rect 8250 13380 8290 13420
rect 8500 13380 8540 13420
rect 8720 13380 8760 13420
rect 9270 13380 9310 13420
rect 9550 13380 9590 13420
rect 9800 13380 9840 13420
rect 10020 13380 10060 13420
rect 10570 13380 10610 13420
rect 410 13270 450 13310
rect 1360 13250 1400 13290
rect 1490 13260 1530 13300
rect 2430 13260 2470 13300
rect 3990 13260 4030 13300
rect 6594 13270 6634 13310
rect 350 13000 390 13040
rect 2020 13030 2060 13070
rect 2540 13030 2580 13070
rect 2760 12830 2800 12870
rect 4260 13020 4300 13060
rect 11302 13588 11336 13622
rect 11822 13588 11856 13622
rect 12342 13588 12376 13622
rect 11228 13420 11268 13460
rect 11228 13320 11268 13360
rect 11340 13420 11380 13460
rect 11340 13320 11380 13360
rect 11748 13420 11788 13460
rect 11748 13320 11788 13360
rect 11860 13420 11900 13460
rect 11860 13320 11900 13360
rect 12268 13420 12308 13460
rect 12268 13320 12308 13360
rect 12380 13420 12420 13460
rect 12380 13320 12420 13360
rect 11274 13208 11308 13242
rect 11794 13208 11828 13242
rect 12314 13208 12348 13242
rect 10774 13008 10808 13042
rect 1050 12710 1090 12750
rect 1240 12710 1280 12750
rect 1360 12730 1400 12770
rect 2170 12710 2210 12750
rect 2300 12710 2340 12750
rect 3430 12710 3470 12750
rect 3650 12710 3690 12750
rect 4780 12700 4820 12740
rect 5190 12700 5230 12740
rect 7140 12710 7180 12750
rect 7720 12710 7760 12750
rect 8440 12710 8480 12750
rect 9020 12710 9060 12750
rect 9740 12710 9780 12750
rect 10320 12710 10360 12750
rect 730 12600 770 12640
rect 1150 12600 1190 12640
rect 1820 12600 1860 12640
rect 2390 12600 2430 12640
rect 3100 12600 3140 12640
rect 3530 12600 3570 12640
rect 3970 12600 4010 12640
rect 4220 12600 4260 12640
rect 4440 12600 4480 12640
rect 4910 12600 4950 12640
rect 5350 12600 5390 12640
rect 5970 12600 6010 12640
rect 6310 12600 6350 12640
rect 6670 12600 6710 12640
rect 7270 12600 7310 12640
rect 7610 12600 7650 12640
rect 7970 12600 8010 12640
rect 8570 12600 8610 12640
rect 8910 12600 8950 12640
rect 9270 12600 9310 12640
rect 9870 12600 9910 12640
rect 10210 12600 10250 12640
rect 10570 12600 10610 12640
rect 11274 12818 11308 12852
rect 11794 12818 11828 12852
rect 12314 12818 12348 12852
rect 11228 12700 11268 12740
rect 11228 12600 11268 12640
rect 11228 12500 11268 12540
rect 11228 12400 11268 12440
rect 11340 12700 11380 12740
rect 11340 12600 11380 12640
rect 11340 12500 11380 12540
rect 11340 12400 11380 12440
rect 11748 12700 11788 12740
rect 11748 12600 11788 12640
rect 11748 12500 11788 12540
rect 11748 12400 11788 12440
rect 11860 12700 11900 12740
rect 11860 12600 11900 12640
rect 11860 12500 11900 12540
rect 11860 12400 11900 12440
rect 12268 12700 12308 12740
rect 12268 12600 12308 12640
rect 12268 12500 12308 12540
rect 12268 12400 12308 12440
rect 12380 12700 12420 12740
rect 12380 12600 12420 12640
rect 12380 12500 12420 12540
rect 12380 12400 12420 12440
rect 11302 12238 11336 12272
rect 11822 12238 11856 12272
rect 12342 12238 12376 12272
rect 11230 12120 11270 12160
rect 11230 12020 11270 12060
rect 11230 11920 11270 11960
rect 11230 11820 11270 11860
rect 11230 11720 11270 11760
rect 11230 11620 11270 11660
rect 11340 12120 11380 12160
rect 11340 12020 11380 12060
rect 11340 11920 11380 11960
rect 11340 11820 11380 11860
rect 11340 11720 11380 11760
rect 11340 11620 11380 11660
rect 11750 12120 11790 12160
rect 11750 12020 11790 12060
rect 11750 11920 11790 11960
rect 11750 11820 11790 11860
rect 11750 11720 11790 11760
rect 11750 11620 11790 11660
rect 11860 12120 11900 12160
rect 11860 12020 11900 12060
rect 11860 11920 11900 11960
rect 11860 11820 11900 11860
rect 11860 11720 11900 11760
rect 11860 11620 11900 11660
rect 12270 12120 12310 12160
rect 12270 12020 12310 12060
rect 12270 11920 12310 11960
rect 12270 11820 12310 11860
rect 12270 11720 12310 11760
rect 12270 11620 12310 11660
rect 12380 12120 12420 12160
rect 12380 12020 12420 12060
rect 12380 11920 12420 11960
rect 12380 11820 12420 11860
rect 12380 11720 12420 11760
rect 12380 11620 12420 11660
rect 11420 11350 11460 11390
rect 11940 11350 11980 11390
rect 12460 11350 12500 11390
rect 12980 11350 13020 11390
rect 11230 11230 11270 11270
rect 11230 11130 11270 11170
rect 11230 11030 11270 11070
rect 11230 10930 11270 10970
rect 11610 11230 11650 11270
rect 11610 11130 11650 11170
rect 11610 11030 11650 11070
rect 11610 10930 11650 10970
rect 11750 11230 11790 11270
rect 11750 11130 11790 11170
rect 11750 11030 11790 11070
rect 11750 10930 11790 10970
rect 12130 11230 12170 11270
rect 12130 11130 12170 11170
rect 12130 11030 12170 11070
rect 12130 10930 12170 10970
rect 12270 11230 12310 11270
rect 12270 11130 12310 11170
rect 12270 11030 12310 11070
rect 12270 10930 12310 10970
rect 12650 11230 12690 11270
rect 12650 11130 12690 11170
rect 12650 11030 12690 11070
rect 12650 10930 12690 10970
rect 12790 11230 12830 11270
rect 12790 11130 12830 11170
rect 12790 11030 12830 11070
rect 12790 10930 12830 10970
rect 13170 11230 13210 11270
rect 13170 11130 13210 11170
rect 13170 11030 13210 11070
rect 13170 10930 13210 10970
rect 11610 10800 11650 10840
rect 12130 10800 12170 10840
rect 12650 10800 12690 10840
rect 13170 10800 13210 10840
rect 1280 10400 1320 10440
rect 1500 10400 1540 10440
rect 1800 10400 1840 10440
rect 2020 10400 2060 10440
rect 2180 10400 2220 10440
rect 2400 10400 2440 10440
rect 2700 10400 2740 10440
rect 2920 10400 2960 10440
rect 3220 10400 3260 10440
rect 3660 10400 3700 10440
rect 3990 10400 4030 10440
rect 4420 10400 4460 10440
rect 4810 10400 4850 10440
rect 5200 10400 5240 10440
rect 11010 10450 11080 10520
rect 1690 10290 1730 10330
rect 1160 9910 1200 9950
rect 3410 10290 3450 10330
rect 5490 10290 5530 10330
rect 3060 9940 3100 9980
rect 4150 9900 4190 9940
rect 4280 9930 4320 9970
rect 6030 9950 6070 9990
rect 5720 9870 5760 9910
rect 7570 9840 7610 9880
rect 10410 9840 10450 9880
rect 7570 9720 7610 9760
rect 7570 9620 7610 9660
rect 7570 9520 7610 9560
rect 3280 9330 3320 9370
rect 7570 9420 7610 9460
rect 7790 9720 7830 9760
rect 7790 9620 7830 9660
rect 7790 9520 7830 9560
rect 7790 9420 7830 9460
rect 8010 9720 8050 9760
rect 8010 9620 8050 9660
rect 8010 9520 8050 9560
rect 8010 9420 8050 9460
rect 8230 9720 8270 9760
rect 8230 9620 8270 9660
rect 8230 9520 8270 9560
rect 8230 9420 8270 9460
rect 8450 9720 8490 9760
rect 8450 9620 8490 9660
rect 8450 9520 8490 9560
rect 8450 9420 8490 9460
rect 8670 9720 8710 9760
rect 8670 9620 8710 9660
rect 8670 9520 8710 9560
rect 8670 9420 8710 9460
rect 8890 9720 8930 9760
rect 8990 9720 9030 9760
rect 9090 9720 9130 9760
rect 8890 9620 8930 9660
rect 8990 9620 9030 9660
rect 9090 9620 9130 9660
rect 8890 9520 8930 9560
rect 8990 9520 9030 9560
rect 9090 9520 9130 9560
rect 8890 9420 8930 9460
rect 8990 9420 9030 9460
rect 9090 9420 9130 9460
rect 9310 9720 9350 9760
rect 9310 9620 9350 9660
rect 9310 9520 9350 9560
rect 9310 9420 9350 9460
rect 9530 9720 9570 9760
rect 9530 9620 9570 9660
rect 9530 9520 9570 9560
rect 9530 9420 9570 9460
rect 9750 9720 9790 9760
rect 9750 9620 9790 9660
rect 9750 9520 9790 9560
rect 9750 9420 9790 9460
rect 9970 9720 10010 9760
rect 9970 9620 10010 9660
rect 9970 9520 10010 9560
rect 9970 9420 10010 9460
rect 10190 9720 10230 9760
rect 10190 9620 10230 9660
rect 10190 9520 10230 9560
rect 10190 9420 10230 9460
rect 10410 9720 10450 9760
rect 10410 9620 10450 9660
rect 10410 9520 10450 9560
rect 10410 9420 10450 9460
rect 8230 9300 8270 9340
rect 1280 9220 1320 9260
rect 2020 9220 2060 9260
rect 2180 9220 2220 9260
rect 2920 9220 2960 9260
rect 3170 9220 3210 9260
rect 3360 9220 3400 9260
rect 3440 9220 3480 9260
rect 3650 9220 3690 9260
rect 3980 9220 4020 9260
rect 4420 9220 4460 9260
rect 4810 9220 4850 9260
rect 5200 9220 5240 9260
rect 5880 9220 5920 9260
rect 9400 9270 9440 9310
rect 10100 9270 10140 9310
rect 10770 9270 10840 9340
rect 1730 9110 1770 9150
rect 4850 9110 4890 9150
rect 5490 9110 5530 9150
rect 1160 8530 1200 8570
rect 7810 8730 7850 8770
rect 3080 8540 3120 8580
rect 4110 8540 4150 8580
rect 4260 8530 4300 8570
rect 7370 8620 7410 8660
rect 6030 8490 6070 8530
rect 7370 8520 7410 8560
rect 7370 8420 7410 8460
rect 7370 8320 7410 8360
rect 7590 8620 7630 8660
rect 7590 8520 7630 8560
rect 7590 8420 7630 8460
rect 7590 8320 7630 8360
rect 9840 8770 9880 8810
rect 10100 8770 10140 8810
rect 10770 8740 10840 8810
rect 7810 8620 7850 8660
rect 7810 8520 7850 8560
rect 7810 8420 7850 8460
rect 7810 8320 7850 8360
rect 8030 8620 8070 8660
rect 8030 8520 8070 8560
rect 8030 8420 8070 8460
rect 8030 8320 8070 8360
rect 8250 8620 8290 8660
rect 8350 8620 8390 8660
rect 8450 8620 8490 8660
rect 8250 8520 8290 8560
rect 8350 8520 8390 8560
rect 8450 8520 8490 8560
rect 8250 8420 8290 8460
rect 8350 8420 8390 8460
rect 8450 8420 8490 8460
rect 8250 8320 8290 8360
rect 8350 8320 8390 8360
rect 8450 8320 8490 8360
rect 8670 8620 8710 8660
rect 8670 8520 8710 8560
rect 8670 8420 8710 8460
rect 8670 8320 8710 8360
rect 8890 8620 8930 8660
rect 8890 8520 8930 8560
rect 8890 8420 8930 8460
rect 8890 8320 8930 8360
rect 9110 8620 9150 8660
rect 9110 8520 9150 8560
rect 9110 8420 9150 8460
rect 9110 8320 9150 8360
rect 9330 8620 9370 8660
rect 9430 8620 9470 8660
rect 9530 8620 9570 8660
rect 9330 8520 9370 8560
rect 9430 8520 9470 8560
rect 9530 8520 9570 8560
rect 9330 8420 9370 8460
rect 9430 8420 9470 8460
rect 9530 8420 9570 8460
rect 9330 8320 9370 8360
rect 9430 8320 9470 8360
rect 9530 8320 9570 8360
rect 9750 8620 9790 8660
rect 9750 8520 9790 8560
rect 9750 8420 9790 8460
rect 9750 8320 9790 8360
rect 9970 8620 10010 8660
rect 9970 8520 10010 8560
rect 9970 8420 10010 8460
rect 9970 8320 10010 8360
rect 10190 8620 10230 8660
rect 10190 8520 10230 8560
rect 10190 8420 10230 8460
rect 10190 8320 10230 8360
rect 10410 8620 10450 8660
rect 10410 8520 10450 8560
rect 10410 8420 10450 8460
rect 10410 8320 10450 8360
rect 4930 8150 4970 8190
rect 5560 8150 5600 8190
rect 7370 8200 7410 8240
rect 10410 8200 10450 8240
rect 1280 8040 1320 8080
rect 1500 8040 1540 8080
rect 1800 8040 1840 8080
rect 2030 8040 2070 8080
rect 2180 8040 2220 8080
rect 2400 8040 2440 8080
rect 2700 8040 2740 8080
rect 2920 8040 2960 8080
rect 3320 8040 3360 8080
rect 3650 8040 3690 8080
rect 3980 8040 4020 8080
rect 4420 8040 4460 8080
rect 5200 8040 5240 8080
rect 5880 8040 5920 8080
rect 11120 7950 11190 8020
rect 11240 7200 11300 7260
rect -340 6920 -300 6960
rect 980 6920 1020 6960
rect 1560 6920 1600 6960
rect 2880 6920 2920 6960
rect -420 6800 -380 6840
rect -340 6800 -300 6840
rect -420 6700 -380 6740
rect -340 6700 -300 6740
rect -230 6800 -190 6840
rect -230 6700 -190 6740
rect -120 6800 -80 6840
rect -120 6700 -80 6740
rect -10 6800 30 6840
rect -10 6700 30 6740
rect 100 6800 140 6840
rect 100 6700 140 6740
rect 210 6800 250 6840
rect 210 6700 250 6740
rect 320 6800 360 6840
rect 320 6700 360 6740
rect 430 6800 470 6840
rect 430 6700 470 6740
rect 540 6800 580 6840
rect 540 6700 580 6740
rect 650 6800 690 6840
rect 650 6700 690 6740
rect 760 6800 800 6840
rect 760 6700 800 6740
rect 870 6800 910 6840
rect 870 6700 910 6740
rect 980 6800 1020 6840
rect 1060 6800 1100 6840
rect 980 6700 1020 6740
rect 1060 6700 1100 6740
rect 1480 6800 1520 6840
rect 1560 6800 1600 6840
rect 1480 6700 1520 6740
rect 1560 6700 1600 6740
rect 1670 6800 1710 6840
rect 1670 6700 1710 6740
rect 1780 6800 1820 6840
rect 1780 6700 1820 6740
rect 1890 6800 1930 6840
rect 1890 6700 1930 6740
rect 2000 6800 2040 6840
rect 2000 6700 2040 6740
rect 2110 6800 2150 6840
rect 2110 6700 2150 6740
rect 2220 6800 2260 6840
rect 2220 6700 2260 6740
rect 2330 6800 2370 6840
rect 2330 6700 2370 6740
rect 2440 6800 2480 6840
rect 2440 6700 2480 6740
rect 2550 6800 2590 6840
rect 2550 6700 2590 6740
rect 2660 6800 2700 6840
rect 2660 6700 2700 6740
rect 2770 6800 2810 6840
rect 2770 6700 2810 6740
rect 2880 6800 2920 6840
rect 2960 6800 3000 6840
rect 2880 6700 2920 6740
rect 2960 6700 3000 6740
rect 11040 6690 11043 6730
rect 11043 6690 11077 6730
rect 11077 6690 11080 6730
rect -172 6588 -138 6622
rect -62 6588 -28 6622
rect 48 6588 82 6622
rect 158 6588 192 6622
rect 268 6588 302 6622
rect 378 6588 412 6622
rect 488 6588 522 6622
rect 598 6588 632 6622
rect 708 6588 742 6622
rect 818 6588 852 6622
rect 1728 6588 1762 6622
rect 1838 6588 1872 6622
rect 1948 6588 1982 6622
rect 2058 6588 2092 6622
rect 2168 6588 2202 6622
rect 2278 6588 2312 6622
rect 2388 6588 2422 6622
rect 2498 6588 2532 6622
rect 2608 6588 2642 6622
rect 2718 6588 2752 6622
rect -350 6320 -310 6360
rect 10 6320 50 6360
rect 370 6320 410 6360
rect 730 6320 770 6360
rect 1090 6320 1130 6360
rect 1450 6320 1490 6360
rect 1810 6320 1850 6360
rect 2170 6320 2210 6360
rect 2530 6320 2570 6360
rect 2890 6320 2930 6360
rect 7170 6300 7210 6340
rect -350 6200 -310 6240
rect -350 6100 -310 6140
rect -350 6000 -310 6040
rect -350 5900 -310 5940
rect -350 5800 -310 5840
rect -350 5700 -310 5740
rect -170 6200 -130 6240
rect -170 6100 -130 6140
rect -170 6000 -130 6040
rect -170 5900 -130 5940
rect -170 5800 -130 5840
rect -170 5700 -130 5740
rect 10 6200 50 6240
rect 10 6100 50 6140
rect 10 6000 50 6040
rect 10 5900 50 5940
rect 10 5800 50 5840
rect 10 5700 50 5740
rect 190 6200 230 6240
rect 190 6100 230 6140
rect 190 6000 230 6040
rect 190 5900 230 5940
rect 190 5800 230 5840
rect 190 5700 230 5740
rect 370 6200 410 6240
rect 370 6100 410 6140
rect 370 6000 410 6040
rect 370 5900 410 5940
rect 370 5800 410 5840
rect 370 5700 410 5740
rect 550 6200 590 6240
rect 550 6100 590 6140
rect 550 6000 590 6040
rect 550 5900 590 5940
rect 550 5800 590 5840
rect 550 5700 590 5740
rect 730 6200 770 6240
rect 730 6100 770 6140
rect 730 6000 770 6040
rect 730 5900 770 5940
rect 730 5800 770 5840
rect 730 5700 770 5740
rect 910 6200 950 6240
rect 910 6100 950 6140
rect 910 6000 950 6040
rect 910 5900 950 5940
rect 910 5800 950 5840
rect 910 5700 950 5740
rect 1090 6200 1130 6240
rect 1090 6100 1130 6140
rect 1090 6000 1130 6040
rect 1090 5900 1130 5940
rect 1090 5800 1130 5840
rect 1090 5700 1130 5740
rect 1270 6200 1310 6240
rect 1270 6100 1310 6140
rect 1270 6000 1310 6040
rect 1270 5900 1310 5940
rect 1270 5800 1310 5840
rect 1270 5700 1310 5740
rect 1450 6200 1490 6240
rect 1450 6100 1490 6140
rect 1450 6000 1490 6040
rect 1450 5900 1490 5940
rect 1450 5800 1490 5840
rect 1450 5700 1490 5740
rect 1630 6200 1670 6240
rect 1630 6100 1670 6140
rect 1630 6000 1670 6040
rect 1630 5900 1670 5940
rect 1630 5800 1670 5840
rect 1630 5700 1670 5740
rect 1810 6200 1850 6240
rect 1810 6100 1850 6140
rect 1810 6000 1850 6040
rect 1810 5900 1850 5940
rect 1810 5800 1850 5840
rect 1810 5700 1850 5740
rect 1990 6200 2030 6240
rect 1990 6100 2030 6140
rect 1990 6000 2030 6040
rect 1990 5900 2030 5940
rect 1990 5800 2030 5840
rect 1990 5700 2030 5740
rect 2170 6200 2210 6240
rect 2170 6100 2210 6140
rect 2170 6000 2210 6040
rect 2170 5900 2210 5940
rect 2170 5800 2210 5840
rect 2170 5700 2210 5740
rect 2350 6200 2390 6240
rect 2350 6100 2390 6140
rect 2350 6000 2390 6040
rect 2350 5900 2390 5940
rect 2350 5800 2390 5840
rect 2350 5700 2390 5740
rect 2530 6200 2570 6240
rect 2530 6100 2570 6140
rect 2530 6000 2570 6040
rect 2530 5900 2570 5940
rect 2530 5800 2570 5840
rect 2530 5700 2570 5740
rect 2710 6200 2750 6240
rect 2710 6100 2750 6140
rect 2710 6000 2750 6040
rect 2710 5900 2750 5940
rect 2710 5800 2750 5840
rect 2710 5700 2750 5740
rect 2890 6200 2930 6240
rect 2890 6100 2930 6140
rect 3520 6120 3560 6160
rect 3740 6120 3780 6160
rect 3960 6120 4000 6160
rect 2890 6000 2930 6040
rect 2890 5900 2930 5940
rect 3520 6000 3560 6040
rect 3520 5900 3560 5940
rect 3630 6000 3670 6040
rect 3630 5900 3670 5940
rect 3740 6000 3780 6040
rect 3740 5900 3780 5940
rect 3850 6000 3890 6040
rect 3850 5900 3890 5940
rect 3960 6000 4000 6040
rect 3960 5900 4000 5940
rect 2890 5800 2930 5840
rect 3620 5780 3660 5820
rect 3740 5780 3780 5820
rect 7630 5980 7670 6030
rect 7630 5840 7670 5890
rect 8030 5980 8070 6030
rect 8030 5840 8070 5890
rect 8430 5980 8470 6030
rect 8430 5840 8470 5890
rect 8830 5980 8870 6030
rect 8830 5840 8870 5890
rect 9230 5980 9270 6030
rect 9230 5840 9270 5890
rect 3860 5780 3900 5820
rect 2890 5700 2930 5740
rect 7430 5720 7470 5760
rect 9010 5680 9050 5720
rect 9430 5720 9470 5760
rect 11250 6291 11288 6688
rect 11250 5720 11288 6117
rect -80 5580 -40 5620
rect 100 5580 140 5620
rect 280 5580 320 5620
rect 460 5580 500 5620
rect 640 5580 680 5620
rect 820 5580 860 5620
rect 1000 5580 1040 5620
rect 1180 5580 1220 5620
rect 1360 5580 1400 5620
rect 1540 5580 1580 5620
rect 1720 5580 1760 5620
rect 1900 5580 1940 5620
rect 2080 5580 2120 5620
rect 2260 5580 2300 5620
rect 2440 5580 2480 5620
rect 2620 5580 2660 5620
rect 7870 5570 7910 5610
rect 10150 5570 10190 5610
rect 9010 5460 9050 5500
rect 7480 5300 7520 5340
rect 7610 5300 7650 5340
rect 7740 5300 7780 5340
rect 7870 5300 7910 5340
rect 8000 5300 8040 5340
rect 8130 5300 8170 5340
rect 8260 5300 8300 5340
rect 8620 5300 8660 5340
rect 8750 5300 8790 5340
rect 8880 5300 8920 5340
rect 9010 5300 9050 5340
rect 9140 5300 9180 5340
rect 9270 5300 9310 5340
rect 9400 5300 9440 5340
rect 7740 5180 7780 5220
rect 8790 5180 8830 5220
rect 9230 5180 9270 5220
rect 11470 5260 11540 5330
rect 10770 5180 10810 5220
rect 9930 5060 9970 5100
rect 11640 5010 11680 5050
rect 7650 4840 7690 4880
rect 8090 4840 8130 4880
rect 8880 4850 8920 4890
rect 9930 4840 9970 4880
rect -1450 4760 -1410 4800
rect 950 4760 990 4800
rect 1590 4760 1630 4800
rect 3990 4760 4030 4800
rect 10770 4840 10810 4880
rect 7480 4720 7520 4760
rect -1450 4640 -1410 4680
rect -1450 4540 -1410 4580
rect -1330 4640 -1290 4680
rect -1330 4540 -1290 4580
rect -1210 4640 -1170 4680
rect -1210 4540 -1170 4580
rect -1090 4640 -1050 4680
rect -1090 4540 -1050 4580
rect -970 4640 -930 4680
rect -970 4540 -930 4580
rect -850 4640 -810 4680
rect -850 4540 -810 4580
rect -730 4640 -690 4680
rect -730 4540 -690 4580
rect -610 4640 -570 4680
rect -610 4540 -570 4580
rect -490 4640 -450 4680
rect -490 4540 -450 4580
rect -370 4640 -330 4680
rect -370 4540 -330 4580
rect -250 4640 -210 4680
rect -250 4540 -210 4580
rect -130 4640 -90 4680
rect -130 4540 -90 4580
rect -10 4640 30 4680
rect -10 4540 30 4580
rect 110 4640 150 4680
rect 110 4540 150 4580
rect 230 4640 270 4680
rect 230 4540 270 4580
rect 350 4640 390 4680
rect 350 4540 390 4580
rect 470 4640 510 4680
rect 470 4540 510 4580
rect 590 4640 630 4680
rect 590 4540 630 4580
rect 710 4640 750 4680
rect 710 4540 750 4580
rect 830 4640 870 4680
rect 830 4540 870 4580
rect 950 4640 990 4680
rect 950 4540 990 4580
rect 1590 4640 1630 4680
rect 1590 4540 1630 4580
rect 1710 4640 1750 4680
rect 1710 4540 1750 4580
rect 1830 4640 1870 4680
rect 1830 4540 1870 4580
rect 1950 4640 1990 4680
rect 1950 4540 1990 4580
rect 2070 4640 2110 4680
rect 2070 4540 2110 4580
rect 2190 4640 2230 4680
rect 2190 4540 2230 4580
rect 2310 4640 2350 4680
rect 2310 4540 2350 4580
rect 2430 4640 2470 4680
rect 2430 4540 2470 4580
rect 2550 4640 2590 4680
rect 2550 4540 2590 4580
rect 2670 4640 2710 4680
rect 2670 4540 2710 4580
rect 2790 4640 2830 4680
rect 2790 4540 2830 4580
rect 2910 4640 2950 4680
rect 2910 4540 2950 4580
rect 3030 4640 3070 4680
rect 3030 4540 3070 4580
rect 3150 4640 3190 4680
rect 3150 4540 3190 4580
rect 3270 4640 3310 4680
rect 3270 4540 3310 4580
rect 3390 4640 3430 4680
rect 3390 4540 3430 4580
rect 3510 4640 3550 4680
rect 3510 4540 3550 4580
rect 3630 4640 3670 4680
rect 3630 4540 3670 4580
rect 3750 4640 3790 4680
rect 3750 4540 3790 4580
rect 3870 4640 3910 4680
rect 3870 4540 3910 4580
rect 3990 4640 4030 4680
rect 7480 4620 7520 4660
rect 7610 4720 7650 4760
rect 7610 4620 7650 4660
rect 7740 4720 7780 4760
rect 7740 4620 7780 4660
rect 7870 4720 7910 4760
rect 7870 4620 7910 4660
rect 8000 4720 8040 4760
rect 8000 4620 8040 4660
rect 8130 4720 8170 4760
rect 8130 4620 8170 4660
rect 8260 4720 8300 4760
rect 8260 4620 8300 4660
rect 8620 4720 8660 4760
rect 8620 4620 8660 4660
rect 8750 4720 8790 4760
rect 8750 4620 8790 4660
rect 8880 4720 8920 4760
rect 8880 4620 8920 4660
rect 9010 4720 9050 4760
rect 9010 4620 9050 4660
rect 9140 4720 9180 4760
rect 9140 4620 9180 4660
rect 9270 4720 9310 4760
rect 9270 4620 9310 4660
rect 9400 4720 9440 4760
rect 9400 4620 9440 4660
rect 11470 4750 11540 4820
rect 3990 4540 4030 4580
rect -1270 4410 -1230 4450
rect -1090 4420 -1050 4460
rect -610 4420 -570 4460
rect -370 4420 -330 4460
rect 110 4420 150 4460
rect 350 4420 390 4460
rect 770 4420 810 4460
rect 1770 4420 1810 4460
rect 2190 4420 2230 4460
rect 2430 4420 2470 4460
rect 2910 4420 2950 4460
rect 3150 4420 3190 4460
rect 3630 4420 3670 4460
rect 3810 4410 3850 4450
rect 7950 4460 7990 4500
rect 9030 4350 9070 4390
rect 10150 4350 10190 4390
rect 7550 4190 7590 4230
rect 9550 4190 9590 4230
rect 7550 4070 7590 4110
rect 7550 3970 7590 4010
rect 7550 3870 7590 3910
rect -446 3818 -412 3852
rect -288 3818 -254 3852
rect 36 3818 70 3852
rect 190 3818 224 3852
rect 514 3818 548 3852
rect 830 3770 870 3810
rect -610 3700 -570 3740
rect -490 3700 -450 3740
rect -370 3700 -330 3740
rect -250 3700 -210 3740
rect -130 3700 -90 3740
rect -10 3700 30 3740
rect 110 3700 150 3740
rect 230 3700 270 3740
rect 350 3700 390 3740
rect 470 3700 510 3740
rect 590 3700 630 3740
rect 830 3690 870 3730
rect -547 3588 -513 3622
rect -187 3588 -153 3622
rect -67 3588 -33 3622
rect 293 3588 327 3622
rect 413 3588 447 3622
rect 830 3610 870 3650
rect 1710 3770 1750 3810
rect 2032 3818 2066 3852
rect 2356 3818 2390 3852
rect 2510 3818 2544 3852
rect 2834 3818 2868 3852
rect 2992 3818 3026 3852
rect 7550 3770 7590 3810
rect 1710 3690 1750 3730
rect 1950 3700 1990 3740
rect 2070 3700 2110 3740
rect 2190 3700 2230 3740
rect 2310 3700 2350 3740
rect 2430 3700 2470 3740
rect 2550 3700 2590 3740
rect 2670 3700 2710 3740
rect 2790 3700 2830 3740
rect 2910 3700 2950 3740
rect 3030 3700 3070 3740
rect 3150 3700 3190 3740
rect 7550 3670 7590 3710
rect 7750 4070 7790 4110
rect 7750 3970 7790 4010
rect 7750 3870 7790 3910
rect 7750 3770 7790 3810
rect 7750 3670 7790 3710
rect 7950 4070 7990 4110
rect 7950 3970 7990 4010
rect 7950 3870 7990 3910
rect 7950 3770 7990 3810
rect 7950 3670 7990 3710
rect 8150 4070 8190 4110
rect 8150 3970 8190 4010
rect 8150 3870 8190 3910
rect 8150 3770 8190 3810
rect 8150 3670 8190 3710
rect 8350 4070 8390 4110
rect 8350 3970 8390 4010
rect 8350 3870 8390 3910
rect 8350 3770 8390 3810
rect 8350 3670 8390 3710
rect 8550 4070 8590 4110
rect 8550 3970 8590 4010
rect 8550 3870 8590 3910
rect 8550 3770 8590 3810
rect 8550 3670 8590 3710
rect 8750 4070 8790 4110
rect 8750 3970 8790 4010
rect 8750 3870 8790 3910
rect 8750 3770 8790 3810
rect 8750 3670 8790 3710
rect 8950 4070 8990 4110
rect 8950 3970 8990 4010
rect 8950 3870 8990 3910
rect 8950 3770 8990 3810
rect 8950 3670 8990 3710
rect 9150 4070 9190 4110
rect 9150 3970 9190 4010
rect 9150 3870 9190 3910
rect 9150 3770 9190 3810
rect 9150 3670 9190 3710
rect 9350 4070 9390 4110
rect 9350 3970 9390 4010
rect 9350 3870 9390 3910
rect 9350 3770 9390 3810
rect 9350 3670 9390 3710
rect 9550 4070 9590 4110
rect 9550 3970 9590 4010
rect 9550 3870 9590 3910
rect 9550 3770 9590 3810
rect 9550 3670 9590 3710
rect 1710 3610 1750 3650
rect 2133 3588 2167 3622
rect 2253 3588 2287 3622
rect 2613 3588 2647 3622
rect 2733 3588 2767 3622
rect 3093 3588 3127 3622
rect 8350 3550 8390 3590
rect 8750 3550 8790 3590
rect -1230 3170 -1190 3210
rect -1050 3210 -1010 3250
rect -810 3210 -770 3250
rect -570 3210 -530 3250
rect -330 3210 -290 3250
rect 310 3210 350 3250
rect 550 3210 590 3250
rect 790 3210 830 3250
rect 1090 3180 1130 3220
rect 1450 3180 1490 3220
rect 1750 3210 1790 3250
rect 1990 3210 2030 3250
rect 2230 3210 2270 3250
rect 2870 3210 2910 3250
rect 3110 3210 3150 3250
rect 3350 3210 3390 3250
rect 3590 3210 3630 3250
rect 11250 3827 11288 4224
rect 11040 3160 11043 3200
rect 11043 3160 11077 3200
rect 11077 3160 11080 3200
rect 11250 3200 11288 3597
rect 3770 3090 3810 3130
rect 3770 2990 3810 3030
rect 3770 2890 3810 2930
rect 3770 2790 3810 2830
rect 11240 2820 11300 2880
rect 3770 2690 3810 2730
rect -70 2570 -30 2610
rect 2610 2570 2650 2610
rect -810 2300 -770 2340
rect -650 2300 -610 2340
rect -490 2300 -450 2340
rect -330 2300 -290 2340
rect -170 2300 -130 2340
rect -10 2300 30 2340
rect 150 2300 190 2340
rect 310 2300 350 2340
rect 470 2300 510 2340
rect 630 2300 670 2340
rect 790 2300 830 2340
rect 950 2300 990 2340
rect 1110 2300 1150 2340
rect 1270 2300 1310 2340
rect 1430 2300 1470 2340
rect 1590 2300 1630 2340
rect 1750 2300 1790 2340
rect 1910 2300 1950 2340
rect 2070 2300 2110 2340
rect 2230 2300 2270 2340
rect 2390 2300 2430 2340
rect 2550 2300 2590 2340
rect 2710 2300 2750 2340
rect 2870 2300 2910 2340
rect 3030 2300 3070 2340
rect 3190 2300 3230 2340
rect -890 2130 -850 2170
rect 3500 2170 3540 2210
rect 3500 2090 3540 2130
rect 572 1730 622 1780
rect 1970 1730 2020 1780
rect -330 1164 -324 1170
rect -324 1164 -296 1170
rect -330 1136 -296 1164
rect -230 1136 -196 1170
rect -130 1136 -96 1170
rect -30 1164 2 1170
rect 2 1164 4 1170
rect 70 1164 92 1170
rect 92 1164 104 1170
rect 170 1164 182 1170
rect 182 1164 204 1170
rect -30 1136 4 1164
rect 70 1136 104 1164
rect 170 1136 204 1164
rect -330 1036 -296 1070
rect -230 1036 -196 1070
rect -130 1036 -96 1070
rect -30 1036 4 1070
rect 70 1036 104 1070
rect 170 1036 204 1070
rect -330 936 -296 970
rect -230 936 -196 970
rect -130 936 -96 970
rect -30 936 4 970
rect 70 936 104 970
rect 170 936 204 970
rect -330 838 -296 870
rect -330 836 -324 838
rect -324 836 -296 838
rect -230 836 -196 870
rect -130 836 -96 870
rect -30 838 4 870
rect 70 838 104 870
rect 170 838 204 870
rect -30 836 2 838
rect 2 836 4 838
rect 70 836 92 838
rect 92 836 104 838
rect 170 836 182 838
rect 182 836 204 838
rect -330 748 -296 770
rect -330 736 -324 748
rect -324 736 -296 748
rect -230 736 -196 770
rect -130 736 -96 770
rect -30 748 4 770
rect 70 748 104 770
rect 170 748 204 770
rect -30 736 2 748
rect 2 736 4 748
rect 70 736 92 748
rect 92 736 104 748
rect 170 736 182 748
rect 182 736 204 748
rect -330 658 -296 670
rect -330 636 -324 658
rect -324 636 -296 658
rect -230 636 -196 670
rect -130 636 -96 670
rect -30 658 4 670
rect 70 658 104 670
rect 170 658 204 670
rect -30 636 2 658
rect 2 636 4 658
rect 70 636 92 658
rect 92 636 104 658
rect 170 636 182 658
rect 182 636 204 658
rect 1030 1164 1036 1170
rect 1036 1164 1064 1170
rect 1030 1136 1064 1164
rect 1130 1136 1164 1170
rect 1230 1136 1264 1170
rect 1330 1164 1362 1170
rect 1362 1164 1364 1170
rect 1430 1164 1452 1170
rect 1452 1164 1464 1170
rect 1530 1164 1542 1170
rect 1542 1164 1564 1170
rect 1330 1136 1364 1164
rect 1430 1136 1464 1164
rect 1530 1136 1564 1164
rect 1030 1036 1064 1070
rect 1130 1036 1164 1070
rect 1230 1036 1264 1070
rect 1330 1036 1364 1070
rect 1430 1036 1464 1070
rect 1530 1036 1564 1070
rect 1030 936 1064 970
rect 1130 936 1164 970
rect 1230 936 1264 970
rect 1330 936 1364 970
rect 1430 936 1464 970
rect 1530 936 1564 970
rect 1030 838 1064 870
rect 1030 836 1036 838
rect 1036 836 1064 838
rect 1130 836 1164 870
rect 1230 836 1264 870
rect 1330 838 1364 870
rect 1430 838 1464 870
rect 1530 838 1564 870
rect 1330 836 1362 838
rect 1362 836 1364 838
rect 1430 836 1452 838
rect 1452 836 1464 838
rect 1530 836 1542 838
rect 1542 836 1564 838
rect 1030 748 1064 770
rect 1030 736 1036 748
rect 1036 736 1064 748
rect 1130 736 1164 770
rect 1230 736 1264 770
rect 1330 748 1364 770
rect 1430 748 1464 770
rect 1530 748 1564 770
rect 1330 736 1362 748
rect 1362 736 1364 748
rect 1430 736 1452 748
rect 1452 736 1464 748
rect 1530 736 1542 748
rect 1542 736 1564 748
rect 1030 658 1064 670
rect 1030 636 1036 658
rect 1036 636 1064 658
rect 1130 636 1164 670
rect 1230 636 1264 670
rect 1330 658 1364 670
rect 1430 658 1464 670
rect 1530 658 1564 670
rect 1330 636 1362 658
rect 1362 636 1364 658
rect 1430 636 1452 658
rect 1452 636 1464 658
rect 1530 636 1542 658
rect 1542 636 1564 658
rect 2390 1164 2396 1170
rect 2396 1164 2424 1170
rect 2390 1136 2424 1164
rect 2490 1136 2524 1170
rect 2590 1136 2624 1170
rect 2690 1164 2722 1170
rect 2722 1164 2724 1170
rect 2790 1164 2812 1170
rect 2812 1164 2824 1170
rect 2890 1164 2902 1170
rect 2902 1164 2924 1170
rect 2690 1136 2724 1164
rect 2790 1136 2824 1164
rect 2890 1136 2924 1164
rect 2390 1036 2424 1070
rect 2490 1036 2524 1070
rect 2590 1036 2624 1070
rect 2690 1036 2724 1070
rect 2790 1036 2824 1070
rect 2890 1036 2924 1070
rect 2390 936 2424 970
rect 2490 936 2524 970
rect 2590 936 2624 970
rect 2690 936 2724 970
rect 2790 936 2824 970
rect 2890 936 2924 970
rect 2390 838 2424 870
rect 2390 836 2396 838
rect 2396 836 2424 838
rect 2490 836 2524 870
rect 2590 836 2624 870
rect 2690 838 2724 870
rect 2790 838 2824 870
rect 2890 838 2924 870
rect 2690 836 2722 838
rect 2722 836 2724 838
rect 2790 836 2812 838
rect 2812 836 2824 838
rect 2890 836 2902 838
rect 2902 836 2924 838
rect 2390 748 2424 770
rect 2390 736 2396 748
rect 2396 736 2424 748
rect 2490 736 2524 770
rect 2590 736 2624 770
rect 2690 748 2724 770
rect 2790 748 2824 770
rect 2890 748 2924 770
rect 2690 736 2722 748
rect 2722 736 2724 748
rect 2790 736 2812 748
rect 2812 736 2824 748
rect 2890 736 2902 748
rect 2902 736 2924 748
rect 2390 658 2424 670
rect 2390 636 2396 658
rect 2396 636 2424 658
rect 2490 636 2524 670
rect 2590 636 2624 670
rect 2690 658 2724 670
rect 2790 658 2824 670
rect 2890 658 2924 670
rect 2690 636 2722 658
rect 2722 636 2724 658
rect 2790 636 2812 658
rect 2812 636 2824 658
rect 2890 636 2902 658
rect 2902 636 2924 658
rect -3520 -1301 -3482 -904
rect -3520 -2110 -3482 -1713
rect -3520 -2267 -3480 -2240
rect -2400 -896 -2360 -506
rect -2740 -2120 -2700 -1730
rect -3520 -2280 -3480 -2267
rect -2730 -2270 -2690 -2240
rect -1620 -370 -1580 20
rect -1290 -2110 -1250 -1720
rect -330 -196 -324 -190
rect -324 -196 -296 -190
rect -330 -224 -296 -196
rect -230 -224 -196 -190
rect -130 -224 -96 -190
rect -30 -196 2 -190
rect 2 -196 4 -190
rect 70 -196 92 -190
rect 92 -196 104 -190
rect 170 -196 182 -190
rect 182 -196 204 -190
rect -30 -224 4 -196
rect 70 -224 104 -196
rect 170 -224 204 -196
rect -330 -324 -296 -290
rect -230 -324 -196 -290
rect -130 -324 -96 -290
rect -30 -324 4 -290
rect 70 -324 104 -290
rect 170 -324 204 -290
rect -330 -424 -296 -390
rect -230 -424 -196 -390
rect -130 -424 -96 -390
rect -30 -424 4 -390
rect 70 -424 104 -390
rect 170 -424 204 -390
rect -330 -522 -296 -490
rect -330 -524 -324 -522
rect -324 -524 -296 -522
rect -230 -524 -196 -490
rect -130 -524 -96 -490
rect -30 -522 4 -490
rect 70 -522 104 -490
rect 170 -522 204 -490
rect -30 -524 2 -522
rect 2 -524 4 -522
rect 70 -524 92 -522
rect 92 -524 104 -522
rect 170 -524 182 -522
rect 182 -524 204 -522
rect -330 -612 -296 -590
rect -330 -624 -324 -612
rect -324 -624 -296 -612
rect -230 -624 -196 -590
rect -130 -624 -96 -590
rect -30 -612 4 -590
rect 70 -612 104 -590
rect 170 -612 204 -590
rect -30 -624 2 -612
rect 2 -624 4 -612
rect 70 -624 92 -612
rect 92 -624 104 -612
rect 170 -624 182 -612
rect 182 -624 204 -612
rect -330 -702 -296 -690
rect -330 -724 -324 -702
rect -324 -724 -296 -702
rect -230 -724 -196 -690
rect -130 -724 -96 -690
rect -30 -702 4 -690
rect 70 -702 104 -690
rect 170 -702 204 -690
rect -30 -724 2 -702
rect 2 -724 4 -702
rect 70 -724 92 -702
rect 92 -724 104 -702
rect 170 -724 182 -702
rect 182 -724 204 -702
rect 1030 -196 1036 -190
rect 1036 -196 1064 -190
rect 1030 -224 1064 -196
rect 1130 -224 1164 -190
rect 1230 -224 1264 -190
rect 1330 -196 1362 -190
rect 1362 -196 1364 -190
rect 1430 -196 1452 -190
rect 1452 -196 1464 -190
rect 1530 -196 1542 -190
rect 1542 -196 1564 -190
rect 1330 -224 1364 -196
rect 1430 -224 1464 -196
rect 1530 -224 1564 -196
rect 1030 -324 1064 -290
rect 1130 -324 1164 -290
rect 1230 -324 1264 -290
rect 1330 -324 1364 -290
rect 1430 -324 1464 -290
rect 1530 -324 1564 -290
rect 1030 -424 1064 -390
rect 1130 -424 1164 -390
rect 1230 -424 1264 -390
rect 1330 -424 1364 -390
rect 1430 -424 1464 -390
rect 1530 -424 1564 -390
rect 1030 -522 1064 -490
rect 1030 -524 1036 -522
rect 1036 -524 1064 -522
rect 1130 -524 1164 -490
rect 1230 -524 1264 -490
rect 1330 -522 1364 -490
rect 1430 -522 1464 -490
rect 1530 -522 1564 -490
rect 1330 -524 1362 -522
rect 1362 -524 1364 -522
rect 1430 -524 1452 -522
rect 1452 -524 1464 -522
rect 1530 -524 1542 -522
rect 1542 -524 1564 -522
rect 1030 -612 1064 -590
rect 1030 -624 1036 -612
rect 1036 -624 1064 -612
rect 1130 -624 1164 -590
rect 1230 -624 1264 -590
rect 1330 -612 1364 -590
rect 1430 -612 1464 -590
rect 1530 -612 1564 -590
rect 1330 -624 1362 -612
rect 1362 -624 1364 -612
rect 1430 -624 1452 -612
rect 1452 -624 1464 -612
rect 1530 -624 1542 -612
rect 1542 -624 1564 -612
rect 1030 -702 1064 -690
rect 1030 -724 1036 -702
rect 1036 -724 1064 -702
rect 1130 -724 1164 -690
rect 1230 -724 1264 -690
rect 1330 -702 1364 -690
rect 1430 -702 1464 -690
rect 1530 -702 1564 -690
rect 1330 -724 1362 -702
rect 1362 -724 1364 -702
rect 1430 -724 1452 -702
rect 1452 -724 1464 -702
rect 1530 -724 1542 -702
rect 1542 -724 1564 -702
rect 2390 -196 2396 -190
rect 2396 -196 2424 -190
rect 2390 -224 2424 -196
rect 2490 -224 2524 -190
rect 2590 -224 2624 -190
rect 2690 -196 2722 -190
rect 2722 -196 2724 -190
rect 2790 -196 2812 -190
rect 2812 -196 2824 -190
rect 2890 -196 2902 -190
rect 2902 -196 2924 -190
rect 2690 -224 2724 -196
rect 2790 -224 2824 -196
rect 2890 -224 2924 -196
rect 2390 -324 2424 -290
rect 2490 -324 2524 -290
rect 2590 -324 2624 -290
rect 2690 -324 2724 -290
rect 2790 -324 2824 -290
rect 2890 -324 2924 -290
rect 2390 -424 2424 -390
rect 2490 -424 2524 -390
rect 2590 -424 2624 -390
rect 2690 -424 2724 -390
rect 2790 -424 2824 -390
rect 2890 -424 2924 -390
rect 2390 -522 2424 -490
rect 2390 -524 2396 -522
rect 2396 -524 2424 -522
rect 2490 -524 2524 -490
rect 2590 -524 2624 -490
rect 2690 -522 2724 -490
rect 2790 -522 2824 -490
rect 2890 -522 2924 -490
rect 2690 -524 2722 -522
rect 2722 -524 2724 -522
rect 2790 -524 2812 -522
rect 2812 -524 2824 -522
rect 2890 -524 2902 -522
rect 2902 -524 2924 -522
rect 2390 -612 2424 -590
rect 2390 -624 2396 -612
rect 2396 -624 2424 -612
rect 2490 -624 2524 -590
rect 2590 -624 2624 -590
rect 2690 -612 2724 -590
rect 2790 -612 2824 -590
rect 2890 -612 2924 -590
rect 2690 -624 2722 -612
rect 2722 -624 2724 -612
rect 2790 -624 2812 -612
rect 2812 -624 2824 -612
rect 2890 -624 2902 -612
rect 2902 -624 2924 -612
rect 2390 -702 2424 -690
rect 2390 -724 2396 -702
rect 2396 -724 2424 -702
rect 2490 -724 2524 -690
rect 2590 -724 2624 -690
rect 2690 -702 2724 -690
rect 2790 -702 2824 -690
rect 2890 -702 2924 -690
rect 2690 -724 2722 -702
rect 2722 -724 2724 -702
rect 2790 -724 2812 -702
rect 2812 -724 2824 -702
rect 2890 -724 2902 -702
rect 2902 -724 2924 -702
rect -1290 -2267 -1250 -2240
rect -2730 -2280 -2690 -2270
rect -1290 -2280 -1250 -2267
rect -330 -1556 -324 -1550
rect -324 -1556 -296 -1550
rect -330 -1584 -296 -1556
rect -230 -1584 -196 -1550
rect -130 -1584 -96 -1550
rect -30 -1556 2 -1550
rect 2 -1556 4 -1550
rect 70 -1556 92 -1550
rect 92 -1556 104 -1550
rect 170 -1556 182 -1550
rect 182 -1556 204 -1550
rect -30 -1584 4 -1556
rect 70 -1584 104 -1556
rect 170 -1584 204 -1556
rect -330 -1684 -296 -1650
rect -230 -1684 -196 -1650
rect -130 -1684 -96 -1650
rect -30 -1684 4 -1650
rect 70 -1684 104 -1650
rect 170 -1684 204 -1650
rect -330 -1784 -296 -1750
rect -230 -1784 -196 -1750
rect -130 -1784 -96 -1750
rect -30 -1784 4 -1750
rect 70 -1784 104 -1750
rect 170 -1784 204 -1750
rect -330 -1882 -296 -1850
rect -330 -1884 -324 -1882
rect -324 -1884 -296 -1882
rect -230 -1884 -196 -1850
rect -130 -1884 -96 -1850
rect -30 -1882 4 -1850
rect 70 -1882 104 -1850
rect 170 -1882 204 -1850
rect -30 -1884 2 -1882
rect 2 -1884 4 -1882
rect 70 -1884 92 -1882
rect 92 -1884 104 -1882
rect 170 -1884 182 -1882
rect 182 -1884 204 -1882
rect -330 -1972 -296 -1950
rect -330 -1984 -324 -1972
rect -324 -1984 -296 -1972
rect -230 -1984 -196 -1950
rect -130 -1984 -96 -1950
rect -30 -1972 4 -1950
rect 70 -1972 104 -1950
rect 170 -1972 204 -1950
rect -30 -1984 2 -1972
rect 2 -1984 4 -1972
rect 70 -1984 92 -1972
rect 92 -1984 104 -1972
rect 170 -1984 182 -1972
rect 182 -1984 204 -1972
rect -330 -2062 -296 -2050
rect -330 -2084 -324 -2062
rect -324 -2084 -296 -2062
rect -230 -2084 -196 -2050
rect -130 -2084 -96 -2050
rect -30 -2062 4 -2050
rect 70 -2062 104 -2050
rect 170 -2062 204 -2050
rect -30 -2084 2 -2062
rect 2 -2084 4 -2062
rect 70 -2084 92 -2062
rect 92 -2084 104 -2062
rect 170 -2084 182 -2062
rect 182 -2084 204 -2062
rect 1030 -1556 1036 -1550
rect 1036 -1556 1064 -1550
rect 1030 -1584 1064 -1556
rect 1130 -1584 1164 -1550
rect 1230 -1584 1264 -1550
rect 1330 -1556 1362 -1550
rect 1362 -1556 1364 -1550
rect 1430 -1556 1452 -1550
rect 1452 -1556 1464 -1550
rect 1530 -1556 1542 -1550
rect 1542 -1556 1564 -1550
rect 1330 -1584 1364 -1556
rect 1430 -1584 1464 -1556
rect 1530 -1584 1564 -1556
rect 1030 -1684 1064 -1650
rect 1130 -1684 1164 -1650
rect 1230 -1684 1264 -1650
rect 1330 -1684 1364 -1650
rect 1430 -1684 1464 -1650
rect 1530 -1684 1564 -1650
rect 1030 -1784 1064 -1750
rect 1130 -1784 1164 -1750
rect 1230 -1784 1264 -1750
rect 1330 -1784 1364 -1750
rect 1430 -1784 1464 -1750
rect 1530 -1784 1564 -1750
rect 1030 -1882 1064 -1850
rect 1030 -1884 1036 -1882
rect 1036 -1884 1064 -1882
rect 1130 -1884 1164 -1850
rect 1230 -1884 1264 -1850
rect 1330 -1882 1364 -1850
rect 1430 -1882 1464 -1850
rect 1530 -1882 1564 -1850
rect 1330 -1884 1362 -1882
rect 1362 -1884 1364 -1882
rect 1430 -1884 1452 -1882
rect 1452 -1884 1464 -1882
rect 1530 -1884 1542 -1882
rect 1542 -1884 1564 -1882
rect 1030 -1972 1064 -1950
rect 1030 -1984 1036 -1972
rect 1036 -1984 1064 -1972
rect 1130 -1984 1164 -1950
rect 1230 -1984 1264 -1950
rect 1330 -1972 1364 -1950
rect 1430 -1972 1464 -1950
rect 1530 -1972 1564 -1950
rect 1330 -1984 1362 -1972
rect 1362 -1984 1364 -1972
rect 1430 -1984 1452 -1972
rect 1452 -1984 1464 -1972
rect 1530 -1984 1542 -1972
rect 1542 -1984 1564 -1972
rect 1030 -2062 1064 -2050
rect 1030 -2084 1036 -2062
rect 1036 -2084 1064 -2062
rect 1130 -2084 1164 -2050
rect 1230 -2084 1264 -2050
rect 1330 -2062 1364 -2050
rect 1430 -2062 1464 -2050
rect 1530 -2062 1564 -2050
rect 1330 -2084 1362 -2062
rect 1362 -2084 1364 -2062
rect 1430 -2084 1452 -2062
rect 1452 -2084 1464 -2062
rect 1530 -2084 1542 -2062
rect 1542 -2084 1564 -2062
rect 2390 -1556 2396 -1550
rect 2396 -1556 2424 -1550
rect 2390 -1584 2424 -1556
rect 2490 -1584 2524 -1550
rect 2590 -1584 2624 -1550
rect 2690 -1556 2722 -1550
rect 2722 -1556 2724 -1550
rect 2790 -1556 2812 -1550
rect 2812 -1556 2824 -1550
rect 2890 -1556 2902 -1550
rect 2902 -1556 2924 -1550
rect 2690 -1584 2724 -1556
rect 2790 -1584 2824 -1556
rect 2890 -1584 2924 -1556
rect 2390 -1684 2424 -1650
rect 2490 -1684 2524 -1650
rect 2590 -1684 2624 -1650
rect 2690 -1684 2724 -1650
rect 2790 -1684 2824 -1650
rect 2890 -1684 2924 -1650
rect 2390 -1784 2424 -1750
rect 2490 -1784 2524 -1750
rect 2590 -1784 2624 -1750
rect 2690 -1784 2724 -1750
rect 2790 -1784 2824 -1750
rect 2890 -1784 2924 -1750
rect 2390 -1882 2424 -1850
rect 2390 -1884 2396 -1882
rect 2396 -1884 2424 -1882
rect 2490 -1884 2524 -1850
rect 2590 -1884 2624 -1850
rect 2690 -1882 2724 -1850
rect 2790 -1882 2824 -1850
rect 2890 -1882 2924 -1850
rect 2690 -1884 2722 -1882
rect 2722 -1884 2724 -1882
rect 2790 -1884 2812 -1882
rect 2812 -1884 2824 -1882
rect 2890 -1884 2902 -1882
rect 2902 -1884 2924 -1882
rect 2390 -1972 2424 -1950
rect 2390 -1984 2396 -1972
rect 2396 -1984 2424 -1972
rect 2490 -1984 2524 -1950
rect 2590 -1984 2624 -1950
rect 2690 -1972 2724 -1950
rect 2790 -1972 2824 -1950
rect 2890 -1972 2924 -1950
rect 2690 -1984 2722 -1972
rect 2722 -1984 2724 -1972
rect 2790 -1984 2812 -1972
rect 2812 -1984 2824 -1972
rect 2890 -1984 2902 -1972
rect 2902 -1984 2924 -1972
rect 2390 -2062 2424 -2050
rect 2390 -2084 2396 -2062
rect 2396 -2084 2424 -2062
rect 2490 -2084 2524 -2050
rect 2590 -2084 2624 -2050
rect 2690 -2062 2724 -2050
rect 2790 -2062 2824 -2050
rect 2890 -2062 2924 -2050
rect 2690 -2084 2722 -2062
rect 2722 -2084 2724 -2062
rect 2790 -2084 2812 -2062
rect 2812 -2084 2824 -2062
rect 2890 -2084 2902 -2062
rect 2902 -2084 2924 -2062
rect 4030 -370 4070 20
rect 3700 -2110 3740 -1720
rect 3700 -2267 3740 -2240
rect 4813 -1508 4851 -1111
rect 4813 -2107 4851 -1710
rect 4810 -2264 4850 -2240
rect 5600 -1301 5638 -904
rect 5600 -2110 5638 -1713
rect 3700 -2280 3740 -2267
rect 4810 -2280 4850 -2264
rect 5600 -2267 5640 -2240
rect 5600 -2280 5640 -2267
rect 1270 -2580 1310 -2540
rect 1270 -2660 1310 -2620
rect 1270 -2740 1310 -2700
rect 3020 -3160 3417 -3122
rect 4923 -3160 5320 -3122
rect 4150 -3333 4190 -3310
rect 4150 -3350 4190 -3333
<< metal1 >>
rect 11320 14830 11400 14840
rect 11320 14770 11330 14830
rect 11390 14770 11400 14830
rect 10820 14720 11060 14730
rect 10820 14660 10830 14720
rect 10890 14660 10910 14720
rect 10970 14660 10990 14720
rect 11050 14660 11060 14720
rect 10820 14640 11060 14660
rect 10820 14580 10830 14640
rect 10890 14580 10910 14640
rect 10970 14580 10990 14640
rect 11050 14580 11060 14640
rect 10820 14560 11060 14580
rect 10820 14500 10830 14560
rect 10890 14500 10910 14560
rect 10970 14500 10990 14560
rect 11050 14500 11060 14560
rect 550 13430 630 13440
rect 550 13370 560 13430
rect 620 13370 630 13430
rect 550 13360 630 13370
rect 770 13430 850 13440
rect 770 13370 780 13430
rect 840 13370 850 13430
rect 770 13360 850 13370
rect 1240 13430 1320 13440
rect 1240 13370 1250 13430
rect 1310 13370 1320 13430
rect 1240 13360 1320 13370
rect 1580 13430 1660 13440
rect 1580 13370 1590 13430
rect 1650 13370 1660 13430
rect 1580 13360 1660 13370
rect 1800 13430 1880 13440
rect 1800 13370 1810 13430
rect 1870 13370 1880 13430
rect 1800 13360 1880 13370
rect 2240 13430 2320 13440
rect 2240 13370 2250 13430
rect 2310 13370 2320 13430
rect 2240 13360 2320 13370
rect 2920 13430 3000 13440
rect 2920 13370 2930 13430
rect 2990 13370 3000 13430
rect 2920 13360 3000 13370
rect 3140 13430 3220 13440
rect 3140 13370 3150 13430
rect 3210 13370 3220 13430
rect 3140 13360 3220 13370
rect 3610 13430 3690 13440
rect 3610 13370 3620 13430
rect 3680 13370 3690 13430
rect 3610 13360 3690 13370
rect 4070 13430 4150 13440
rect 4070 13370 4080 13430
rect 4140 13370 4150 13430
rect 4070 13360 4150 13370
rect 4420 13430 4500 13440
rect 4420 13370 4430 13430
rect 4490 13370 4500 13430
rect 4420 13360 4500 13370
rect 4670 13430 4750 13440
rect 4670 13370 4680 13430
rect 4740 13370 4750 13430
rect 4670 13360 4750 13370
rect 4890 13430 4970 13440
rect 4890 13370 4900 13430
rect 4960 13370 4970 13430
rect 4890 13360 4970 13370
rect 5220 13430 5300 13440
rect 5220 13370 5230 13430
rect 5290 13370 5300 13430
rect 5220 13360 5300 13370
rect 5880 13430 5960 13440
rect 5880 13370 5890 13430
rect 5950 13370 5960 13430
rect 5880 13360 5960 13370
rect 6100 13430 6180 13440
rect 6100 13370 6110 13430
rect 6170 13370 6180 13430
rect 6100 13360 6180 13370
rect 6670 13430 6750 13440
rect 6670 13370 6680 13430
rect 6740 13370 6750 13430
rect 6670 13360 6750 13370
rect 6930 13430 7010 13440
rect 6930 13370 6940 13430
rect 7000 13370 7010 13430
rect 6930 13360 7010 13370
rect 7180 13430 7260 13440
rect 7180 13370 7190 13430
rect 7250 13370 7260 13430
rect 7180 13360 7260 13370
rect 7400 13430 7480 13440
rect 7400 13370 7410 13430
rect 7470 13370 7480 13430
rect 7400 13360 7480 13370
rect 7950 13430 8030 13440
rect 7950 13370 7960 13430
rect 8020 13370 8030 13430
rect 7950 13360 8030 13370
rect 8230 13430 8310 13440
rect 8230 13370 8240 13430
rect 8300 13370 8310 13430
rect 8230 13360 8310 13370
rect 8480 13430 8560 13440
rect 8480 13370 8490 13430
rect 8550 13370 8560 13430
rect 8480 13360 8560 13370
rect 8700 13430 8780 13440
rect 8700 13370 8710 13430
rect 8770 13370 8780 13430
rect 8700 13360 8780 13370
rect 9250 13430 9330 13440
rect 9250 13370 9260 13430
rect 9320 13370 9330 13430
rect 9250 13360 9330 13370
rect 9530 13430 9610 13440
rect 9530 13370 9540 13430
rect 9600 13370 9610 13430
rect 9530 13360 9610 13370
rect 9780 13430 9860 13440
rect 9780 13370 9790 13430
rect 9850 13370 9860 13430
rect 9780 13360 9860 13370
rect 10000 13430 10080 13440
rect 10000 13370 10010 13430
rect 10070 13370 10080 13430
rect 10000 13360 10080 13370
rect 10550 13430 10630 13440
rect 10550 13370 10560 13430
rect 10620 13370 10630 13430
rect 10550 13360 10630 13370
rect 390 13310 470 13330
rect 390 13270 410 13310
rect 450 13290 1420 13310
rect 450 13270 1360 13290
rect 390 13250 470 13270
rect 1340 13250 1360 13270
rect 1400 13250 1420 13290
rect 1470 13300 4050 13320
rect 1470 13260 1490 13300
rect 1530 13280 2430 13300
rect 1530 13260 1550 13280
rect 1470 13250 1550 13260
rect 2410 13260 2430 13280
rect 2470 13280 3990 13300
rect 2470 13260 2490 13280
rect 2410 13250 2490 13260
rect 3970 13260 3990 13280
rect 4030 13260 4050 13300
rect 6584 13310 6650 13330
rect 6584 13290 6594 13310
rect 3970 13250 4050 13260
rect 4240 13270 6594 13290
rect 6634 13270 6650 13310
rect 4240 13250 6650 13270
rect 1340 13230 1420 13250
rect 2000 13070 2080 13090
rect 120 13050 200 13060
rect 120 12990 130 13050
rect 190 12990 200 13050
rect 120 8580 200 12990
rect 330 13050 410 13060
rect 330 12990 340 13050
rect 400 12990 410 13050
rect 2000 13030 2020 13070
rect 2060 13060 2080 13070
rect 2520 13070 2600 13090
rect 2520 13060 2540 13070
rect 2060 13030 2540 13060
rect 2580 13030 2600 13070
rect 2000 13020 2600 13030
rect 4240 13080 4280 13250
rect 10820 13140 11060 14500
rect 11320 14450 11400 14770
rect 11320 14410 11340 14450
rect 11380 14410 11400 14450
rect 11320 14390 11400 14410
rect 11840 14830 11920 14840
rect 11840 14770 11850 14830
rect 11910 14770 11920 14830
rect 11840 14450 11920 14770
rect 11840 14410 11860 14450
rect 11900 14410 11920 14450
rect 11840 14390 11920 14410
rect 12360 14830 12440 14840
rect 12360 14770 12370 14830
rect 12430 14770 12440 14830
rect 12360 14450 12440 14770
rect 12360 14410 12380 14450
rect 12420 14410 12440 14450
rect 12360 14390 12440 14410
rect 12850 14830 12930 14840
rect 12850 14770 12860 14830
rect 12920 14770 12930 14830
rect 12850 14450 12930 14770
rect 12850 14410 12870 14450
rect 12910 14410 12930 14450
rect 12850 14390 12930 14410
rect 13180 14720 13420 14730
rect 13180 14660 13190 14720
rect 13250 14660 13270 14720
rect 13330 14660 13350 14720
rect 13410 14660 13420 14720
rect 13180 14640 13420 14660
rect 13180 14580 13190 14640
rect 13250 14580 13270 14640
rect 13330 14580 13350 14640
rect 13410 14580 13420 14640
rect 13180 14560 13420 14580
rect 13180 14500 13190 14560
rect 13250 14500 13270 14560
rect 13330 14500 13350 14560
rect 13410 14500 13420 14560
rect 11330 14340 11390 14390
rect 11850 14340 11910 14390
rect 12370 14340 12430 14390
rect 11180 14320 11280 14340
rect 11180 14280 11230 14320
rect 11270 14280 11280 14320
rect 11180 14220 11280 14280
rect 11180 14180 11230 14220
rect 11270 14180 11280 14220
rect 11180 14160 11280 14180
rect 11330 14320 11430 14340
rect 11330 14280 11340 14320
rect 11380 14280 11430 14320
rect 11330 14220 11430 14280
rect 11330 14180 11340 14220
rect 11380 14180 11430 14220
rect 11330 14160 11430 14180
rect 11180 13960 11220 14160
rect 11276 14112 11334 14120
rect 11276 14060 11280 14112
rect 11332 14060 11334 14112
rect 11276 14050 11334 14060
rect 11390 13960 11430 14160
rect 11180 13940 11280 13960
rect 11180 13900 11230 13940
rect 11270 13900 11280 13940
rect 11180 13840 11280 13900
rect 11180 13800 11230 13840
rect 11270 13800 11280 13840
rect 11180 13740 11280 13800
rect 11180 13700 11230 13740
rect 11270 13700 11280 13740
rect 11180 13680 11280 13700
rect 11330 13940 11430 13960
rect 11330 13900 11340 13940
rect 11380 13900 11430 13940
rect 11330 13840 11430 13900
rect 11330 13800 11340 13840
rect 11380 13800 11430 13840
rect 11330 13750 11430 13800
rect 11700 14320 11800 14340
rect 11700 14280 11750 14320
rect 11790 14280 11800 14320
rect 11700 14220 11800 14280
rect 11700 14180 11750 14220
rect 11790 14180 11800 14220
rect 11700 14160 11800 14180
rect 11850 14320 11950 14340
rect 11850 14280 11860 14320
rect 11900 14280 11950 14320
rect 11850 14220 11950 14280
rect 11850 14180 11860 14220
rect 11900 14180 11950 14220
rect 11850 14160 11950 14180
rect 11700 13960 11740 14160
rect 11796 14112 11854 14120
rect 11796 14060 11800 14112
rect 11852 14060 11854 14112
rect 11796 14050 11854 14060
rect 11910 13960 11950 14160
rect 11700 13940 11800 13960
rect 11700 13900 11750 13940
rect 11790 13900 11800 13940
rect 11700 13840 11800 13900
rect 11700 13800 11750 13840
rect 11790 13800 11800 13840
rect 11390 13690 11430 13750
rect 11330 13680 11430 13690
rect 11530 13750 11610 13760
rect 11530 13690 11540 13750
rect 11600 13690 11610 13750
rect 11180 13530 11220 13680
rect 11290 13632 11348 13640
rect 11290 13580 11294 13632
rect 11346 13580 11348 13632
rect 11290 13570 11348 13580
rect 11420 13630 11500 13640
rect 11420 13570 11430 13630
rect 11490 13570 11500 13630
rect 11420 13560 11500 13570
rect 11180 13480 11222 13530
rect 11180 13460 11278 13480
rect 11180 13420 11228 13460
rect 11268 13420 11278 13460
rect 11180 13360 11278 13420
rect 11180 13320 11228 13360
rect 11268 13320 11278 13360
rect 11180 13300 11278 13320
rect 11330 13460 11390 13480
rect 11330 13420 11340 13460
rect 11380 13420 11390 13460
rect 11330 13360 11390 13420
rect 11330 13320 11340 13360
rect 11380 13320 11390 13360
rect 11330 13300 11390 13320
rect 11262 13242 11320 13260
rect 11262 13208 11274 13242
rect 11308 13208 11320 13242
rect 11262 13190 11320 13208
rect 11270 13150 11320 13190
rect 10820 13080 10830 13140
rect 10890 13080 10910 13140
rect 10970 13080 10990 13140
rect 11050 13080 11060 13140
rect 4240 13060 4320 13080
rect 10820 13070 11060 13080
rect 4240 13020 4260 13060
rect 4300 13020 4320 13060
rect 4240 13000 4320 13020
rect 10762 13060 11060 13070
rect 10762 13052 10830 13060
rect 10762 13000 10766 13052
rect 10818 13000 10830 13052
rect 10890 13000 10910 13060
rect 10970 13000 10990 13060
rect 11050 13000 11060 13060
rect 10762 12990 11060 13000
rect 330 12980 410 12990
rect 10820 12980 11060 12990
rect 10820 12920 10830 12980
rect 10890 12920 10910 12980
rect 10970 12920 10990 12980
rect 11050 12920 11060 12980
rect 10820 12910 11060 12920
rect 11260 13140 11320 13150
rect 11260 13060 11320 13080
rect 11260 12980 11320 13000
rect 11260 12910 11320 12920
rect 2740 12870 2820 12890
rect 11270 12870 11320 12910
rect 2740 12830 2760 12870
rect 2800 12830 2820 12870
rect 2740 12810 2820 12830
rect 11262 12852 11320 12870
rect 11262 12818 11274 12852
rect 11308 12818 11320 12852
rect 1340 12770 1420 12790
rect 2740 12770 2780 12810
rect 7160 12770 7200 12810
rect 8460 12770 8500 12810
rect 9760 12770 9800 12810
rect 11262 12800 11320 12818
rect 11350 13150 11390 13300
rect 11350 13140 11410 13150
rect 11350 13060 11410 13080
rect 11350 12980 11410 13000
rect 11350 12910 11410 12920
rect 11350 12770 11390 12910
rect 1030 12750 1300 12770
rect 1030 12710 1050 12750
rect 1090 12730 1240 12750
rect 1090 12710 1110 12730
rect 1030 12690 1110 12710
rect 1230 12710 1240 12730
rect 1280 12710 1300 12750
rect 1340 12730 1360 12770
rect 1400 12750 2230 12770
rect 1400 12730 2170 12750
rect 1340 12710 1420 12730
rect 2150 12710 2170 12730
rect 2210 12710 2230 12750
rect 1230 12690 1300 12710
rect 2150 12690 2230 12710
rect 2290 12750 2780 12770
rect 2290 12710 2300 12750
rect 2340 12730 2780 12750
rect 3410 12750 3710 12770
rect 2340 12710 2350 12730
rect 2290 12690 2350 12710
rect 3410 12710 3430 12750
rect 3470 12730 3650 12750
rect 3470 12710 3490 12730
rect 3410 12690 3490 12710
rect 3630 12710 3650 12730
rect 3690 12710 3710 12750
rect 3630 12690 3710 12710
rect 4760 12740 5250 12760
rect 4760 12700 4780 12740
rect 4820 12720 5190 12740
rect 4820 12700 4840 12720
rect 4760 12690 4840 12700
rect 5170 12700 5190 12720
rect 5230 12700 5250 12740
rect 5170 12690 5250 12700
rect 7120 12750 7780 12770
rect 7120 12710 7140 12750
rect 7180 12730 7720 12750
rect 7180 12710 7200 12730
rect 7120 12690 7200 12710
rect 7700 12710 7720 12730
rect 7760 12710 7780 12750
rect 7700 12690 7780 12710
rect 8420 12750 9080 12770
rect 8420 12710 8440 12750
rect 8480 12730 9020 12750
rect 8480 12710 8500 12730
rect 8420 12690 8500 12710
rect 9000 12710 9020 12730
rect 9060 12710 9080 12750
rect 9000 12690 9080 12710
rect 9720 12750 10380 12770
rect 9720 12710 9740 12750
rect 9780 12730 10320 12750
rect 9780 12710 9800 12730
rect 9720 12690 9800 12710
rect 10300 12710 10320 12730
rect 10360 12710 10380 12750
rect 10300 12690 10380 12710
rect 11218 12740 11278 12760
rect 11218 12700 11228 12740
rect 11268 12700 11278 12740
rect 710 12650 790 12660
rect 710 12590 720 12650
rect 780 12590 790 12650
rect 710 12580 790 12590
rect 1130 12650 1210 12660
rect 1130 12590 1140 12650
rect 1200 12590 1210 12650
rect 1130 12580 1210 12590
rect 1800 12650 1880 12660
rect 1800 12590 1810 12650
rect 1870 12590 1880 12650
rect 1800 12580 1880 12590
rect 2370 12650 2450 12660
rect 2370 12590 2380 12650
rect 2440 12590 2450 12650
rect 2370 12580 2450 12590
rect 3080 12650 3160 12660
rect 3080 12590 3090 12650
rect 3150 12590 3160 12650
rect 3080 12580 3160 12590
rect 3510 12650 3590 12660
rect 3510 12590 3520 12650
rect 3580 12590 3590 12650
rect 3510 12580 3590 12590
rect 3950 12650 4030 12660
rect 3950 12590 3960 12650
rect 4020 12590 4030 12650
rect 3950 12580 4030 12590
rect 4200 12650 4280 12660
rect 4200 12590 4210 12650
rect 4270 12590 4280 12650
rect 4200 12580 4280 12590
rect 4420 12650 4500 12660
rect 4420 12590 4430 12650
rect 4490 12590 4500 12650
rect 4420 12580 4500 12590
rect 4890 12650 4970 12660
rect 4890 12590 4900 12650
rect 4960 12590 4970 12650
rect 4890 12580 4970 12590
rect 5330 12650 5410 12660
rect 5330 12590 5340 12650
rect 5400 12590 5410 12650
rect 5330 12580 5410 12590
rect 5950 12650 6030 12660
rect 5950 12590 5960 12650
rect 6020 12590 6030 12650
rect 5950 12580 6030 12590
rect 6290 12650 6370 12660
rect 6290 12590 6300 12650
rect 6360 12590 6370 12650
rect 6290 12580 6370 12590
rect 6650 12650 6730 12660
rect 6650 12590 6660 12650
rect 6720 12590 6730 12650
rect 6650 12580 6730 12590
rect 7250 12650 7330 12660
rect 7250 12590 7260 12650
rect 7320 12590 7330 12650
rect 7250 12580 7330 12590
rect 7590 12650 7670 12660
rect 7590 12590 7600 12650
rect 7660 12590 7670 12650
rect 7590 12580 7670 12590
rect 7950 12650 8030 12660
rect 7950 12590 7960 12650
rect 8020 12590 8030 12650
rect 7950 12580 8030 12590
rect 8550 12650 8630 12660
rect 8550 12590 8560 12650
rect 8620 12590 8630 12650
rect 8550 12580 8630 12590
rect 8890 12650 8970 12660
rect 8890 12590 8900 12650
rect 8960 12590 8970 12650
rect 8890 12580 8970 12590
rect 9250 12650 9330 12660
rect 9250 12590 9260 12650
rect 9320 12590 9330 12650
rect 9250 12580 9330 12590
rect 9850 12650 9930 12660
rect 9850 12590 9860 12650
rect 9920 12590 9930 12650
rect 9850 12580 9930 12590
rect 10190 12650 10270 12660
rect 10190 12590 10200 12650
rect 10260 12590 10270 12650
rect 10190 12580 10270 12590
rect 10550 12650 10630 12660
rect 10550 12590 10560 12650
rect 10620 12590 10630 12650
rect 10550 12580 10630 12590
rect 11218 12640 11278 12700
rect 11218 12600 11228 12640
rect 11268 12600 11278 12640
rect 11218 12540 11278 12600
rect 11218 12500 11228 12540
rect 11268 12500 11278 12540
rect 11218 12440 11278 12500
rect 11218 12400 11228 12440
rect 11268 12400 11278 12440
rect 11218 12380 11278 12400
rect 11330 12740 11390 12770
rect 11330 12700 11340 12740
rect 11380 12700 11390 12740
rect 11330 12640 11390 12700
rect 11330 12600 11340 12640
rect 11380 12600 11390 12640
rect 11330 12540 11390 12600
rect 11330 12500 11340 12540
rect 11380 12500 11390 12540
rect 11330 12440 11390 12500
rect 11330 12400 11340 12440
rect 11380 12400 11390 12440
rect 11330 12380 11390 12400
rect 11220 12180 11260 12380
rect 11290 12282 11348 12290
rect 11290 12230 11294 12282
rect 11346 12230 11348 12282
rect 11290 12220 11348 12230
rect 11440 12180 11500 13560
rect 11530 12290 11610 13690
rect 11700 13740 11800 13800
rect 11700 13700 11750 13740
rect 11790 13700 11800 13740
rect 11700 13680 11800 13700
rect 11850 13940 11950 13960
rect 11850 13900 11860 13940
rect 11900 13900 11950 13940
rect 11850 13840 11950 13900
rect 11850 13800 11860 13840
rect 11900 13800 11950 13840
rect 11850 13750 11950 13800
rect 12220 14320 12320 14340
rect 12220 14280 12270 14320
rect 12310 14280 12320 14320
rect 12220 14220 12320 14280
rect 12220 14180 12270 14220
rect 12310 14180 12320 14220
rect 12220 14160 12320 14180
rect 12370 14320 12470 14340
rect 12370 14280 12380 14320
rect 12420 14280 12470 14320
rect 12370 14220 12470 14280
rect 12370 14180 12380 14220
rect 12420 14180 12470 14220
rect 12370 14160 12470 14180
rect 12860 14320 12920 14390
rect 12860 14280 12870 14320
rect 12910 14280 12920 14320
rect 12860 14220 12920 14280
rect 12860 14180 12870 14220
rect 12910 14180 12920 14220
rect 12860 14160 12920 14180
rect 12970 14320 13030 14340
rect 12970 14280 12980 14320
rect 13020 14280 13030 14320
rect 12970 14220 13030 14280
rect 12970 14180 12980 14220
rect 13020 14180 13030 14220
rect 12220 13960 12260 14160
rect 12316 14112 12374 14120
rect 12316 14060 12320 14112
rect 12372 14060 12374 14112
rect 12316 14050 12374 14060
rect 12430 13960 12470 14160
rect 12884 14112 12942 14120
rect 12884 14060 12886 14112
rect 12938 14060 12942 14112
rect 12884 14050 12942 14060
rect 12220 13940 12320 13960
rect 12220 13900 12270 13940
rect 12310 13900 12320 13940
rect 12220 13840 12320 13900
rect 12220 13800 12270 13840
rect 12310 13800 12320 13840
rect 11910 13690 11950 13750
rect 11850 13680 11950 13690
rect 12050 13750 12130 13760
rect 12050 13690 12060 13750
rect 12120 13690 12130 13750
rect 11700 13530 11740 13680
rect 11810 13632 11868 13640
rect 11810 13580 11814 13632
rect 11866 13580 11868 13632
rect 11810 13570 11868 13580
rect 11940 13630 12020 13640
rect 11940 13570 11950 13630
rect 12010 13570 12020 13630
rect 11940 13560 12020 13570
rect 11700 13480 11742 13530
rect 11700 13460 11798 13480
rect 11700 13420 11748 13460
rect 11788 13420 11798 13460
rect 11700 13360 11798 13420
rect 11700 13320 11748 13360
rect 11788 13320 11798 13360
rect 11700 13300 11798 13320
rect 11850 13460 11910 13480
rect 11850 13420 11860 13460
rect 11900 13420 11910 13460
rect 11850 13360 11910 13420
rect 11850 13320 11860 13360
rect 11900 13320 11910 13360
rect 11850 13300 11910 13320
rect 11782 13242 11840 13260
rect 11782 13208 11794 13242
rect 11828 13208 11840 13242
rect 11782 13190 11840 13208
rect 11790 13150 11840 13190
rect 11780 13140 11840 13150
rect 11780 13060 11840 13080
rect 11780 12980 11840 13000
rect 11780 12910 11840 12920
rect 11790 12870 11840 12910
rect 11782 12852 11840 12870
rect 11782 12818 11794 12852
rect 11828 12818 11840 12852
rect 11782 12800 11840 12818
rect 11870 13150 11910 13300
rect 11870 13140 11930 13150
rect 11870 13060 11930 13080
rect 11870 12980 11930 13000
rect 11870 12910 11930 12920
rect 11870 12770 11910 12910
rect 11738 12740 11798 12760
rect 11738 12700 11748 12740
rect 11788 12700 11798 12740
rect 11738 12640 11798 12700
rect 11738 12600 11748 12640
rect 11788 12600 11798 12640
rect 11738 12540 11798 12600
rect 11738 12500 11748 12540
rect 11788 12500 11798 12540
rect 11738 12440 11798 12500
rect 11738 12400 11748 12440
rect 11788 12400 11798 12440
rect 11738 12380 11798 12400
rect 11850 12740 11910 12770
rect 11850 12700 11860 12740
rect 11900 12700 11910 12740
rect 11850 12640 11910 12700
rect 11850 12600 11860 12640
rect 11900 12600 11910 12640
rect 11850 12540 11910 12600
rect 11850 12500 11860 12540
rect 11900 12500 11910 12540
rect 11850 12440 11910 12500
rect 11850 12400 11860 12440
rect 11900 12400 11910 12440
rect 11850 12380 11910 12400
rect 11530 12230 11540 12290
rect 11600 12230 11610 12290
rect 11530 12220 11610 12230
rect 11220 12160 11280 12180
rect 11220 12120 11230 12160
rect 11270 12120 11280 12160
rect 11220 12060 11280 12120
rect 11220 12020 11230 12060
rect 11270 12020 11280 12060
rect 11220 11960 11280 12020
rect 11220 11920 11230 11960
rect 11270 11920 11280 11960
rect 11220 11860 11280 11920
rect 11220 11820 11230 11860
rect 11270 11820 11280 11860
rect 11220 11760 11280 11820
rect 11220 11720 11230 11760
rect 11270 11720 11280 11760
rect 11220 11660 11280 11720
rect 11220 11620 11230 11660
rect 11270 11620 11280 11660
rect 11220 11270 11280 11620
rect 11330 12170 11390 12180
rect 11330 12060 11390 12110
rect 11420 12170 11500 12180
rect 11420 12110 11430 12170
rect 11490 12110 11500 12170
rect 11420 12100 11500 12110
rect 11740 12180 11780 12380
rect 11810 12282 11868 12290
rect 11810 12230 11814 12282
rect 11866 12230 11868 12282
rect 11810 12220 11868 12230
rect 11960 12180 12020 13560
rect 12050 12290 12130 13690
rect 12220 13740 12320 13800
rect 12220 13700 12270 13740
rect 12310 13700 12320 13740
rect 12220 13680 12320 13700
rect 12370 13940 12470 13960
rect 12370 13900 12380 13940
rect 12420 13900 12470 13940
rect 12370 13840 12470 13900
rect 12370 13800 12380 13840
rect 12420 13800 12470 13840
rect 12370 13750 12470 13800
rect 12430 13690 12470 13750
rect 12370 13680 12470 13690
rect 12570 13750 12650 13760
rect 12570 13690 12580 13750
rect 12640 13690 12650 13750
rect 12220 13530 12260 13680
rect 12330 13632 12388 13640
rect 12330 13580 12334 13632
rect 12386 13580 12388 13632
rect 12330 13570 12388 13580
rect 12460 13630 12540 13640
rect 12460 13570 12470 13630
rect 12530 13570 12540 13630
rect 12460 13560 12540 13570
rect 12220 13480 12262 13530
rect 12220 13460 12318 13480
rect 12220 13420 12268 13460
rect 12308 13420 12318 13460
rect 12220 13360 12318 13420
rect 12220 13320 12268 13360
rect 12308 13320 12318 13360
rect 12220 13300 12318 13320
rect 12370 13460 12430 13480
rect 12370 13420 12380 13460
rect 12420 13420 12430 13460
rect 12370 13360 12430 13420
rect 12370 13320 12380 13360
rect 12420 13320 12430 13360
rect 12370 13300 12430 13320
rect 12302 13242 12360 13260
rect 12302 13208 12314 13242
rect 12348 13208 12360 13242
rect 12302 13190 12360 13208
rect 12310 13150 12360 13190
rect 12300 13140 12360 13150
rect 12300 13060 12360 13080
rect 12300 12980 12360 13000
rect 12300 12910 12360 12920
rect 12310 12870 12360 12910
rect 12302 12852 12360 12870
rect 12302 12818 12314 12852
rect 12348 12818 12360 12852
rect 12302 12800 12360 12818
rect 12390 13150 12430 13300
rect 12390 13140 12450 13150
rect 12390 13060 12450 13080
rect 12390 12980 12450 13000
rect 12390 12910 12450 12920
rect 12390 12770 12430 12910
rect 12258 12740 12318 12760
rect 12258 12700 12268 12740
rect 12308 12700 12318 12740
rect 12258 12640 12318 12700
rect 12258 12600 12268 12640
rect 12308 12600 12318 12640
rect 12258 12540 12318 12600
rect 12258 12500 12268 12540
rect 12308 12500 12318 12540
rect 12258 12440 12318 12500
rect 12258 12400 12268 12440
rect 12308 12400 12318 12440
rect 12258 12380 12318 12400
rect 12370 12740 12430 12770
rect 12370 12700 12380 12740
rect 12420 12700 12430 12740
rect 12370 12640 12430 12700
rect 12370 12600 12380 12640
rect 12420 12600 12430 12640
rect 12370 12540 12430 12600
rect 12370 12500 12380 12540
rect 12420 12500 12430 12540
rect 12370 12440 12430 12500
rect 12370 12400 12380 12440
rect 12420 12400 12430 12440
rect 12370 12380 12430 12400
rect 12050 12230 12060 12290
rect 12120 12230 12130 12290
rect 12050 12220 12130 12230
rect 11740 12160 11800 12180
rect 11740 12120 11750 12160
rect 11790 12120 11800 12160
rect 11330 12020 11340 12060
rect 11380 12020 11390 12060
rect 11330 11960 11390 12020
rect 11330 11920 11340 11960
rect 11380 11920 11390 11960
rect 11330 11860 11390 11920
rect 11330 11820 11340 11860
rect 11380 11820 11390 11860
rect 11330 11760 11390 11820
rect 11330 11720 11340 11760
rect 11380 11720 11390 11760
rect 11330 11660 11390 11720
rect 11330 11620 11340 11660
rect 11380 11620 11390 11660
rect 11330 11590 11390 11620
rect 11740 12060 11800 12120
rect 11740 12020 11750 12060
rect 11790 12020 11800 12060
rect 11740 11960 11800 12020
rect 11740 11920 11750 11960
rect 11790 11920 11800 11960
rect 11740 11860 11800 11920
rect 11740 11820 11750 11860
rect 11790 11820 11800 11860
rect 11740 11760 11800 11820
rect 11740 11720 11750 11760
rect 11790 11720 11800 11760
rect 11740 11660 11800 11720
rect 11740 11620 11750 11660
rect 11790 11620 11800 11660
rect 11320 11580 11400 11590
rect 11320 11520 11330 11580
rect 11390 11520 11400 11580
rect 11320 11510 11400 11520
rect 11590 11580 11670 11590
rect 11590 11520 11600 11580
rect 11660 11520 11670 11580
rect 11590 11510 11670 11520
rect 11400 11400 11480 11410
rect 11400 11340 11410 11400
rect 11470 11340 11480 11400
rect 11400 11330 11480 11340
rect 11220 11230 11230 11270
rect 11270 11230 11280 11270
rect 11220 11170 11280 11230
rect 11220 11130 11230 11170
rect 11270 11130 11280 11170
rect 11220 11070 11280 11130
rect 11220 11030 11230 11070
rect 11270 11030 11280 11070
rect 11220 10970 11280 11030
rect 11220 10930 11230 10970
rect 11270 10930 11280 10970
rect 11220 10910 11280 10930
rect 11600 11270 11660 11510
rect 11600 11230 11610 11270
rect 11650 11230 11660 11270
rect 11600 11170 11660 11230
rect 11600 11130 11610 11170
rect 11650 11130 11660 11170
rect 11600 11070 11660 11130
rect 11600 11030 11610 11070
rect 11650 11030 11660 11070
rect 11600 10970 11660 11030
rect 11600 10930 11610 10970
rect 11650 10930 11660 10970
rect 11600 10860 11660 10930
rect 11740 11270 11800 11620
rect 11850 12170 11910 12180
rect 11850 12060 11910 12110
rect 11940 12170 12020 12180
rect 11940 12110 11950 12170
rect 12010 12110 12020 12170
rect 11940 12100 12020 12110
rect 12260 12180 12300 12380
rect 12330 12282 12388 12290
rect 12330 12230 12334 12282
rect 12386 12230 12388 12282
rect 12330 12220 12388 12230
rect 12480 12180 12540 13560
rect 12570 12290 12650 13690
rect 12570 12230 12580 12290
rect 12640 12230 12650 12290
rect 12570 12220 12650 12230
rect 12260 12160 12320 12180
rect 12260 12120 12270 12160
rect 12310 12120 12320 12160
rect 11850 12020 11860 12060
rect 11900 12020 11910 12060
rect 11850 11960 11910 12020
rect 11850 11920 11860 11960
rect 11900 11920 11910 11960
rect 11850 11860 11910 11920
rect 11850 11820 11860 11860
rect 11900 11820 11910 11860
rect 11850 11760 11910 11820
rect 11850 11720 11860 11760
rect 11900 11720 11910 11760
rect 11850 11660 11910 11720
rect 11850 11620 11860 11660
rect 11900 11620 11910 11660
rect 11850 11590 11910 11620
rect 12260 12060 12320 12120
rect 12260 12020 12270 12060
rect 12310 12020 12320 12060
rect 12260 11960 12320 12020
rect 12260 11920 12270 11960
rect 12310 11920 12320 11960
rect 12260 11860 12320 11920
rect 12260 11820 12270 11860
rect 12310 11820 12320 11860
rect 12260 11760 12320 11820
rect 12260 11720 12270 11760
rect 12310 11720 12320 11760
rect 12260 11660 12320 11720
rect 12260 11620 12270 11660
rect 12310 11620 12320 11660
rect 11840 11580 11920 11590
rect 11840 11520 11850 11580
rect 11910 11520 11920 11580
rect 11840 11510 11920 11520
rect 12110 11580 12190 11590
rect 12110 11520 12120 11580
rect 12180 11520 12190 11580
rect 12110 11510 12190 11520
rect 11920 11400 12000 11410
rect 11920 11340 11930 11400
rect 11990 11340 12000 11400
rect 11920 11330 12000 11340
rect 11740 11230 11750 11270
rect 11790 11230 11800 11270
rect 11740 11170 11800 11230
rect 11740 11130 11750 11170
rect 11790 11130 11800 11170
rect 11740 11070 11800 11130
rect 11740 11030 11750 11070
rect 11790 11030 11800 11070
rect 11740 10970 11800 11030
rect 11740 10930 11750 10970
rect 11790 10930 11800 10970
rect 11740 10910 11800 10930
rect 12120 11270 12180 11510
rect 12120 11230 12130 11270
rect 12170 11230 12180 11270
rect 12120 11170 12180 11230
rect 12120 11130 12130 11170
rect 12170 11130 12180 11170
rect 12120 11070 12180 11130
rect 12120 11030 12130 11070
rect 12170 11030 12180 11070
rect 12120 10970 12180 11030
rect 12120 10930 12130 10970
rect 12170 10930 12180 10970
rect 12120 10860 12180 10930
rect 12260 11270 12320 11620
rect 12370 12170 12430 12180
rect 12370 12060 12430 12110
rect 12460 12170 12540 12180
rect 12460 12110 12470 12170
rect 12530 12110 12540 12170
rect 12460 12100 12540 12110
rect 12370 12020 12380 12060
rect 12420 12020 12430 12060
rect 12370 11960 12430 12020
rect 12370 11920 12380 11960
rect 12420 11920 12430 11960
rect 12370 11860 12430 11920
rect 12370 11820 12380 11860
rect 12420 11820 12430 11860
rect 12370 11760 12430 11820
rect 12370 11720 12380 11760
rect 12420 11720 12430 11760
rect 12370 11660 12430 11720
rect 12370 11620 12380 11660
rect 12420 11620 12430 11660
rect 12370 11590 12430 11620
rect 12360 11580 12440 11590
rect 12360 11520 12370 11580
rect 12430 11520 12440 11580
rect 12360 11510 12440 11520
rect 12630 11580 12710 11590
rect 12630 11520 12640 11580
rect 12700 11520 12710 11580
rect 12630 11510 12710 11520
rect 12440 11400 12520 11410
rect 12440 11340 12450 11400
rect 12510 11340 12520 11400
rect 12440 11330 12520 11340
rect 12260 11230 12270 11270
rect 12310 11230 12320 11270
rect 12260 11170 12320 11230
rect 12260 11130 12270 11170
rect 12310 11130 12320 11170
rect 12260 11070 12320 11130
rect 12260 11030 12270 11070
rect 12310 11030 12320 11070
rect 12260 10970 12320 11030
rect 12260 10930 12270 10970
rect 12310 10930 12320 10970
rect 12260 10910 12320 10930
rect 12640 11270 12700 11510
rect 12640 11230 12650 11270
rect 12690 11230 12700 11270
rect 12640 11170 12700 11230
rect 12640 11130 12650 11170
rect 12690 11130 12700 11170
rect 12640 11070 12700 11130
rect 12640 11030 12650 11070
rect 12690 11030 12700 11070
rect 12640 10970 12700 11030
rect 12640 10930 12650 10970
rect 12690 10930 12700 10970
rect 12640 10860 12700 10930
rect 12780 11400 12840 11410
rect 12780 11270 12840 11340
rect 12970 11400 13030 14180
rect 13180 13140 13420 14500
rect 13180 13080 13190 13140
rect 13250 13080 13270 13140
rect 13330 13080 13350 13140
rect 13410 13080 13420 13140
rect 13180 13060 13420 13080
rect 13180 13000 13190 13060
rect 13250 13000 13270 13060
rect 13330 13000 13350 13060
rect 13410 13000 13420 13060
rect 13180 12980 13420 13000
rect 13180 12920 13190 12980
rect 13250 12920 13270 12980
rect 13330 12920 13350 12980
rect 13410 12920 13420 12980
rect 13180 12910 13420 12920
rect 14010 14110 14090 14120
rect 14010 14050 14020 14110
rect 14080 14050 14090 14110
rect 12970 11330 13030 11340
rect 12780 11230 12790 11270
rect 12830 11230 12840 11270
rect 12780 11170 12840 11230
rect 12780 11130 12790 11170
rect 12830 11130 12840 11170
rect 12780 11070 12840 11130
rect 12780 11030 12790 11070
rect 12830 11030 12840 11070
rect 12780 10970 12840 11030
rect 12780 10930 12790 10970
rect 12830 10930 12840 10970
rect 12780 10910 12840 10930
rect 13160 11270 13220 11290
rect 13160 11230 13170 11270
rect 13210 11230 13220 11270
rect 13160 11170 13220 11230
rect 13160 11130 13170 11170
rect 13210 11130 13220 11170
rect 13160 11070 13220 11130
rect 13160 11030 13170 11070
rect 13210 11030 13220 11070
rect 13160 10970 13220 11030
rect 13160 10930 13170 10970
rect 13210 10930 13220 10970
rect 13160 10860 13220 10930
rect 11590 10840 11670 10860
rect 11590 10800 11610 10840
rect 11650 10800 11670 10840
rect 11590 10750 11670 10800
rect 11590 10690 11600 10750
rect 11660 10690 11670 10750
rect 11590 10680 11670 10690
rect 12110 10840 12190 10860
rect 12110 10800 12130 10840
rect 12170 10800 12190 10840
rect 12110 10750 12190 10800
rect 12110 10690 12120 10750
rect 12180 10690 12190 10750
rect 12110 10680 12190 10690
rect 12630 10840 12710 10860
rect 12630 10800 12650 10840
rect 12690 10800 12710 10840
rect 12630 10750 12710 10800
rect 12630 10690 12640 10750
rect 12700 10690 12710 10750
rect 12630 10680 12710 10690
rect 13150 10840 13230 10860
rect 13150 10800 13170 10840
rect 13210 10800 13230 10840
rect 13150 10750 13230 10800
rect 13150 10690 13160 10750
rect 13220 10690 13230 10750
rect 13150 10680 13230 10690
rect 10990 10520 11100 10540
rect 5700 10510 5780 10520
rect 1260 10450 1340 10460
rect 1260 10390 1270 10450
rect 1330 10390 1340 10450
rect 1260 10380 1340 10390
rect 1480 10450 1560 10460
rect 1480 10390 1490 10450
rect 1550 10390 1560 10450
rect 1480 10380 1560 10390
rect 1780 10450 1860 10460
rect 1780 10390 1790 10450
rect 1850 10390 1860 10450
rect 1780 10380 1860 10390
rect 2000 10450 2080 10460
rect 2000 10390 2010 10450
rect 2070 10390 2080 10450
rect 2000 10380 2080 10390
rect 2160 10450 2240 10460
rect 2160 10390 2170 10450
rect 2230 10390 2240 10450
rect 2160 10380 2240 10390
rect 2380 10450 2460 10460
rect 2380 10390 2390 10450
rect 2450 10390 2460 10450
rect 2380 10380 2460 10390
rect 2680 10450 2760 10460
rect 2680 10390 2690 10450
rect 2750 10390 2760 10450
rect 2680 10380 2760 10390
rect 2900 10450 2980 10460
rect 2900 10390 2910 10450
rect 2970 10390 2980 10450
rect 2900 10380 2980 10390
rect 3200 10450 3280 10460
rect 3200 10390 3210 10450
rect 3270 10390 3280 10450
rect 3200 10380 3280 10390
rect 3640 10450 3720 10460
rect 3640 10390 3650 10450
rect 3710 10390 3720 10450
rect 3640 10380 3720 10390
rect 3970 10450 4050 10460
rect 3970 10390 3980 10450
rect 4040 10390 4050 10450
rect 3970 10380 4050 10390
rect 4400 10450 4480 10460
rect 4400 10390 4410 10450
rect 4470 10390 4480 10450
rect 4400 10380 4480 10390
rect 4790 10450 4870 10460
rect 4790 10390 4800 10450
rect 4860 10390 4870 10450
rect 4790 10380 4870 10390
rect 5180 10450 5260 10460
rect 5180 10390 5190 10450
rect 5250 10390 5260 10450
rect 5180 10380 5260 10390
rect 5700 10450 5710 10510
rect 5770 10450 5780 10510
rect 1670 10340 1750 10350
rect 1670 10280 1680 10340
rect 1740 10280 1750 10340
rect 1670 10270 1750 10280
rect 3390 10340 3470 10350
rect 3390 10280 3400 10340
rect 3460 10280 3470 10340
rect 5470 10340 5550 10350
rect 3390 10270 3470 10280
rect 4240 10320 4320 10330
rect 4240 10260 4250 10320
rect 4310 10260 4320 10320
rect 5470 10280 5480 10340
rect 5540 10280 5550 10340
rect 5470 10270 5550 10280
rect 4240 10250 4320 10260
rect 3040 9990 3120 10000
rect 1140 9960 1220 9970
rect 1140 9900 1150 9960
rect 1210 9900 1220 9960
rect 3040 9930 3050 9990
rect 3110 9930 3120 9990
rect 4260 9990 4300 10250
rect 4260 9970 4340 9990
rect 3040 9920 3120 9930
rect 1140 9890 1220 9900
rect 1260 9270 1340 9280
rect 1260 9210 1270 9270
rect 1330 9210 1340 9270
rect 1260 9200 1340 9210
rect 2000 9270 2080 9280
rect 2000 9210 2010 9270
rect 2070 9210 2080 9270
rect 2000 9200 2080 9210
rect 2160 9270 2240 9280
rect 2160 9210 2170 9270
rect 2230 9210 2240 9270
rect 2160 9200 2240 9210
rect 2900 9270 2980 9280
rect 2900 9210 2910 9270
rect 2970 9210 2980 9270
rect 2900 9200 2980 9210
rect 1710 9160 1790 9170
rect 1710 9100 1720 9160
rect 1780 9100 1790 9160
rect 1710 9090 1790 9100
rect 3080 8600 3120 9920
rect 4130 9950 4210 9960
rect 4130 9890 4140 9950
rect 4200 9890 4210 9950
rect 4260 9930 4280 9970
rect 4320 9930 4340 9970
rect 4260 9910 4340 9930
rect 5700 9920 5780 10450
rect 10990 10450 11010 10520
rect 11080 10450 11100 10520
rect 10990 10430 11100 10450
rect 6410 10340 6490 10350
rect 6410 10280 6420 10340
rect 6480 10280 6490 10340
rect 6010 10000 6090 10010
rect 6010 9940 6020 10000
rect 6080 9940 6090 10000
rect 6010 9930 6090 9940
rect 6300 10000 6380 10010
rect 6300 9940 6310 10000
rect 6370 9940 6380 10000
rect 4130 9880 4210 9890
rect 3260 9380 3340 9390
rect 3260 9320 3270 9380
rect 3330 9320 3340 9380
rect 3150 9270 3230 9280
rect 3150 9210 3160 9270
rect 3220 9210 3230 9270
rect 3150 9200 3230 9210
rect 3260 9170 3300 9320
rect 3340 9270 3500 9280
rect 3340 9210 3350 9270
rect 3410 9210 3430 9270
rect 3490 9210 3500 9270
rect 3340 9200 3500 9210
rect 3630 9270 3710 9280
rect 3630 9210 3640 9270
rect 3700 9210 3710 9270
rect 3630 9200 3710 9210
rect 3960 9270 4040 9280
rect 3960 9210 3970 9270
rect 4030 9210 4040 9270
rect 3960 9200 4040 9210
rect 3240 9160 3320 9170
rect 3240 9100 3250 9160
rect 3310 9100 3320 9160
rect 3240 9090 3320 9100
rect 4170 8600 4210 9880
rect 5700 9860 5710 9920
rect 5770 9860 5780 9920
rect 5700 9850 5780 9860
rect 4400 9270 4480 9280
rect 4400 9210 4410 9270
rect 4470 9210 4480 9270
rect 4400 9200 4480 9210
rect 4790 9270 4870 9280
rect 4790 9210 4800 9270
rect 4860 9210 4870 9270
rect 4790 9200 4870 9210
rect 5000 9270 5080 9280
rect 5000 9210 5010 9270
rect 5070 9210 5080 9270
rect 5000 9200 5080 9210
rect 5180 9270 5260 9280
rect 5180 9210 5190 9270
rect 5250 9210 5260 9270
rect 5180 9200 5260 9210
rect 5860 9270 5940 9280
rect 5860 9210 5870 9270
rect 5930 9210 5940 9270
rect 5860 9200 5940 9210
rect 3060 8590 3140 8600
rect 120 8520 130 8580
rect 190 8520 200 8580
rect 120 8510 200 8520
rect 1140 8580 1220 8590
rect 1140 8520 1150 8580
rect 1210 8520 1220 8580
rect 3060 8530 3070 8590
rect 3130 8530 3140 8590
rect 3060 8520 3140 8530
rect 4090 8590 4210 8600
rect 4090 8530 4100 8590
rect 4160 8530 4210 8590
rect 4090 8520 4210 8530
rect 4240 9150 4320 9160
rect 4240 9090 4250 9150
rect 4310 9090 4320 9150
rect 4660 9100 4670 9160
rect 4730 9100 4740 9160
rect 4830 9100 4840 9160
rect 4900 9100 4910 9160
rect 4240 9080 4320 9090
rect 4240 8590 4280 9080
rect 4240 8570 4320 8590
rect 4240 8530 4260 8570
rect 4300 8530 4320 8570
rect 1140 8510 1220 8520
rect 4240 8510 4320 8530
rect 4680 8100 4720 9100
rect 4830 9090 4910 9100
rect 5020 8210 5060 9200
rect 5470 9160 5550 9170
rect 5470 9100 5480 9160
rect 5540 9100 5550 9160
rect 5470 9090 5550 9100
rect 6190 9160 6270 9170
rect 6190 9100 6200 9160
rect 6260 9100 6270 9160
rect 6190 9010 6270 9100
rect 6300 9120 6380 9940
rect 6410 9230 6490 10280
rect 7550 10000 7630 10010
rect 7550 9940 7560 10000
rect 7620 9940 7630 10000
rect 7550 9880 7630 9940
rect 7550 9840 7570 9880
rect 7610 9840 7630 9880
rect 7550 9760 7630 9840
rect 7550 9720 7570 9760
rect 7610 9720 7630 9760
rect 7550 9660 7630 9720
rect 7550 9620 7570 9660
rect 7610 9620 7630 9660
rect 7550 9560 7630 9620
rect 7550 9520 7570 9560
rect 7610 9520 7630 9560
rect 7550 9460 7630 9520
rect 7550 9420 7570 9460
rect 7610 9420 7630 9460
rect 7550 9400 7630 9420
rect 7770 10000 7850 10010
rect 7770 9940 7780 10000
rect 7840 9940 7850 10000
rect 7770 9760 7850 9940
rect 8210 10000 8290 10010
rect 8210 9940 8220 10000
rect 8280 9940 8290 10000
rect 7770 9720 7790 9760
rect 7830 9720 7850 9760
rect 7770 9660 7850 9720
rect 7770 9620 7790 9660
rect 7830 9620 7850 9660
rect 7770 9560 7850 9620
rect 7770 9520 7790 9560
rect 7830 9520 7850 9560
rect 7770 9460 7850 9520
rect 7770 9420 7790 9460
rect 7830 9420 7850 9460
rect 7770 9400 7850 9420
rect 7990 9760 8070 9780
rect 7990 9720 8010 9760
rect 8050 9720 8070 9760
rect 7990 9660 8070 9720
rect 7990 9620 8010 9660
rect 8050 9620 8070 9660
rect 7990 9560 8070 9620
rect 7990 9520 8010 9560
rect 8050 9520 8070 9560
rect 7990 9460 8070 9520
rect 7990 9420 8010 9460
rect 8050 9420 8070 9460
rect 6410 9170 6420 9230
rect 6480 9170 6490 9230
rect 6410 9160 6490 9170
rect 6930 9350 7010 9360
rect 6930 9290 6940 9350
rect 7000 9290 7010 9350
rect 6300 9060 6310 9120
rect 6370 9060 6380 9120
rect 6300 9050 6380 9060
rect 6190 8950 6200 9010
rect 6260 8950 6270 9010
rect 6190 8940 6270 8950
rect 6660 9010 6900 9020
rect 6660 8950 6670 9010
rect 6730 8950 6750 9010
rect 6810 8950 6830 9010
rect 6890 8950 6900 9010
rect 6190 8900 6270 8910
rect 6190 8840 6200 8900
rect 6260 8840 6270 8900
rect 6010 8540 6090 8550
rect 6010 8480 6020 8540
rect 6080 8480 6090 8540
rect 6010 8470 6090 8480
rect 6190 8540 6270 8840
rect 6190 8480 6200 8540
rect 6260 8480 6270 8540
rect 6190 8470 6270 8480
rect 4910 8200 5060 8210
rect 4910 8140 4920 8200
rect 4980 8140 5060 8200
rect 4910 8130 5060 8140
rect 5540 8200 5620 8210
rect 5540 8140 5550 8200
rect 5610 8140 5620 8200
rect 5540 8130 5620 8140
rect 6110 8200 6190 8210
rect 6110 8140 6120 8200
rect 6180 8140 6190 8200
rect 1260 8090 1340 8100
rect 1260 8030 1270 8090
rect 1330 8030 1340 8090
rect 1260 8020 1340 8030
rect 1480 8090 1560 8100
rect 1480 8030 1490 8090
rect 1550 8030 1560 8090
rect 1480 8020 1560 8030
rect 1780 8090 1860 8100
rect 1780 8030 1790 8090
rect 1850 8030 1860 8090
rect 1780 8020 1860 8030
rect 2010 8090 2090 8100
rect 2010 8030 2020 8090
rect 2080 8030 2090 8090
rect 2010 8020 2090 8030
rect 2160 8090 2240 8100
rect 2160 8030 2170 8090
rect 2230 8030 2240 8090
rect 2160 8020 2240 8030
rect 2380 8090 2460 8100
rect 2380 8030 2390 8090
rect 2450 8030 2460 8090
rect 2380 8020 2460 8030
rect 2680 8090 2760 8100
rect 2680 8030 2690 8090
rect 2750 8030 2760 8090
rect 2680 8020 2760 8030
rect 2900 8090 2980 8100
rect 2900 8030 2910 8090
rect 2970 8030 2980 8090
rect 2900 8020 2980 8030
rect 3300 8090 3380 8100
rect 3300 8030 3310 8090
rect 3370 8030 3380 8090
rect 3300 8020 3380 8030
rect 3630 8090 3710 8100
rect 3630 8030 3640 8090
rect 3700 8030 3710 8090
rect 3630 8020 3710 8030
rect 3960 8090 4040 8100
rect 3960 8030 3970 8090
rect 4030 8030 4040 8090
rect 3960 8020 4040 8030
rect 4400 8090 4480 8100
rect 4400 8030 4410 8090
rect 4470 8030 4480 8090
rect 4400 8020 4480 8030
rect 4660 8090 4740 8100
rect 4660 8030 4670 8090
rect 4730 8030 4740 8090
rect 4660 8020 4740 8030
rect 5180 8090 5260 8100
rect 5180 8030 5190 8090
rect 5250 8030 5260 8090
rect 5180 8020 5260 8030
rect 5860 8090 5940 8100
rect 5860 8030 5870 8090
rect 5930 8030 5940 8090
rect 5860 8020 5940 8030
rect 6110 8020 6190 8140
rect 6110 7960 6120 8020
rect 6180 7960 6190 8020
rect 6110 7950 6190 7960
rect 1650 7250 1730 7260
rect 1650 7190 1660 7250
rect 1720 7190 1730 7250
rect 1650 7170 1730 7190
rect 1650 7110 1660 7170
rect 1720 7110 1730 7170
rect 1650 7090 1730 7110
rect -2310 7080 -2230 7090
rect -2310 7020 -2300 7080
rect -2240 7020 -2230 7080
rect -3540 6630 -3460 6640
rect -3540 6570 -3530 6630
rect -3470 6570 -3460 6630
rect -3540 4810 -3460 6570
rect -3540 4750 -3530 4810
rect -3470 4750 -3460 4810
rect -3540 -900 -3460 4750
rect -2530 5300 -2450 5310
rect -2530 5240 -2520 5300
rect -2460 5240 -2450 5300
rect -2530 2180 -2450 5240
rect -2530 2120 -2520 2180
rect -2460 2120 -2450 2180
rect -2530 2110 -2450 2120
rect -2420 5190 -2340 5200
rect -2420 5130 -2410 5190
rect -2350 5130 -2340 5190
rect -2420 3870 -2340 5130
rect -2420 3810 -2410 3870
rect -2350 3810 -2340 3870
rect -2420 -506 -2340 3810
rect -2310 3640 -2230 7020
rect -250 7080 -170 7090
rect -250 7020 -240 7080
rect -180 7020 -170 7080
rect -250 7010 -170 7020
rect -30 7080 50 7090
rect -30 7020 -20 7080
rect 40 7020 50 7080
rect -30 7010 50 7020
rect 190 7080 270 7090
rect 190 7020 200 7080
rect 260 7020 270 7080
rect 190 7010 270 7020
rect 410 7080 490 7090
rect 410 7020 420 7080
rect 480 7020 490 7080
rect 410 7010 490 7020
rect 630 7080 710 7090
rect 630 7020 640 7080
rect 700 7020 710 7080
rect 630 7010 710 7020
rect 850 7080 930 7090
rect 850 7020 860 7080
rect 920 7020 930 7080
rect 1650 7030 1660 7090
rect 1720 7030 1730 7090
rect 1650 7020 1730 7030
rect 1870 7250 1950 7260
rect 1870 7190 1880 7250
rect 1940 7190 1950 7250
rect 1870 7170 1950 7190
rect 1870 7110 1880 7170
rect 1940 7110 1950 7170
rect 1870 7090 1950 7110
rect 1870 7030 1880 7090
rect 1940 7030 1950 7090
rect 1870 7020 1950 7030
rect 2090 7250 2170 7260
rect 2090 7190 2100 7250
rect 2160 7190 2170 7250
rect 2090 7170 2170 7190
rect 2090 7110 2100 7170
rect 2160 7110 2170 7170
rect 2090 7090 2170 7110
rect 2090 7030 2100 7090
rect 2160 7030 2170 7090
rect 2090 7020 2170 7030
rect 2310 7250 2390 7260
rect 2310 7190 2320 7250
rect 2380 7190 2390 7250
rect 2310 7170 2390 7190
rect 2310 7110 2320 7170
rect 2380 7110 2390 7170
rect 2310 7090 2390 7110
rect 2310 7030 2320 7090
rect 2380 7030 2390 7090
rect 2310 7020 2390 7030
rect 2530 7250 2610 7260
rect 2530 7190 2540 7250
rect 2600 7190 2610 7250
rect 2530 7170 2610 7190
rect 2530 7110 2540 7170
rect 2600 7110 2610 7170
rect 2530 7090 2610 7110
rect 2530 7030 2540 7090
rect 2600 7030 2610 7090
rect 2530 7020 2610 7030
rect 2750 7250 2830 7260
rect 2750 7190 2760 7250
rect 2820 7190 2830 7250
rect 2750 7170 2830 7190
rect 2750 7110 2760 7170
rect 2820 7110 2830 7170
rect 2750 7090 2830 7110
rect 2750 7030 2760 7090
rect 2820 7030 2830 7090
rect 2750 7020 2830 7030
rect 6660 7250 6900 8950
rect 6660 7190 6670 7250
rect 6730 7190 6750 7250
rect 6810 7190 6830 7250
rect 6890 7190 6900 7250
rect 6660 7170 6900 7190
rect 6660 7110 6670 7170
rect 6730 7110 6750 7170
rect 6810 7110 6830 7170
rect 6890 7110 6900 7170
rect 6660 7090 6900 7110
rect 6660 7030 6670 7090
rect 6730 7030 6750 7090
rect 6810 7030 6830 7090
rect 6890 7030 6900 7090
rect 6660 7020 6900 7030
rect 850 7010 930 7020
rect -360 6970 -280 6980
rect -360 6910 -350 6970
rect -290 6910 -280 6970
rect -360 6900 -280 6910
rect -350 6860 -290 6900
rect -430 6840 -290 6860
rect -430 6800 -420 6840
rect -380 6800 -340 6840
rect -300 6800 -290 6840
rect -430 6740 -290 6800
rect -430 6700 -420 6740
rect -380 6700 -340 6740
rect -300 6700 -290 6740
rect -430 6680 -290 6700
rect -240 6840 -180 7010
rect -140 6970 -60 6980
rect -140 6910 -130 6970
rect -70 6910 -60 6970
rect -140 6900 -60 6910
rect -240 6800 -230 6840
rect -190 6800 -180 6840
rect -240 6740 -180 6800
rect -240 6700 -230 6740
rect -190 6700 -180 6740
rect -240 6680 -180 6700
rect -130 6840 -70 6900
rect -130 6800 -120 6840
rect -80 6800 -70 6840
rect -130 6740 -70 6800
rect -130 6700 -120 6740
rect -80 6700 -70 6740
rect -130 6680 -70 6700
rect -20 6840 40 7010
rect 80 6970 160 6980
rect 80 6910 90 6970
rect 150 6910 160 6970
rect 80 6900 160 6910
rect -20 6800 -10 6840
rect 30 6800 40 6840
rect -20 6740 40 6800
rect -20 6700 -10 6740
rect 30 6700 40 6740
rect -20 6680 40 6700
rect 90 6840 150 6900
rect 90 6800 100 6840
rect 140 6800 150 6840
rect 90 6740 150 6800
rect 90 6700 100 6740
rect 140 6700 150 6740
rect 90 6680 150 6700
rect 200 6840 260 7010
rect 300 6970 380 6980
rect 300 6910 310 6970
rect 370 6910 380 6970
rect 300 6900 380 6910
rect 200 6800 210 6840
rect 250 6800 260 6840
rect 200 6740 260 6800
rect 200 6700 210 6740
rect 250 6700 260 6740
rect 200 6680 260 6700
rect 310 6840 370 6900
rect 310 6800 320 6840
rect 360 6800 370 6840
rect 310 6740 370 6800
rect 310 6700 320 6740
rect 360 6700 370 6740
rect 310 6680 370 6700
rect 420 6840 480 7010
rect 520 6970 600 6980
rect 520 6910 530 6970
rect 590 6910 600 6970
rect 520 6900 600 6910
rect 420 6800 430 6840
rect 470 6800 480 6840
rect 420 6740 480 6800
rect 420 6700 430 6740
rect 470 6700 480 6740
rect 420 6680 480 6700
rect 530 6840 590 6900
rect 530 6800 540 6840
rect 580 6800 590 6840
rect 530 6740 590 6800
rect 530 6700 540 6740
rect 580 6700 590 6740
rect 530 6680 590 6700
rect 640 6840 700 7010
rect 740 6970 820 6980
rect 740 6910 750 6970
rect 810 6910 820 6970
rect 740 6900 820 6910
rect 640 6800 650 6840
rect 690 6800 700 6840
rect 640 6740 700 6800
rect 640 6700 650 6740
rect 690 6700 700 6740
rect 640 6680 700 6700
rect 750 6840 810 6900
rect 750 6800 760 6840
rect 800 6800 810 6840
rect 750 6740 810 6800
rect 750 6700 760 6740
rect 800 6700 810 6740
rect 750 6680 810 6700
rect 860 6840 920 7010
rect 960 6970 1040 6980
rect 960 6910 970 6970
rect 1030 6910 1040 6970
rect 960 6900 1040 6910
rect 1540 6970 1620 6980
rect 1540 6910 1550 6970
rect 1610 6910 1620 6970
rect 1540 6900 1620 6910
rect 860 6800 870 6840
rect 910 6800 920 6840
rect 860 6740 920 6800
rect 860 6700 870 6740
rect 910 6700 920 6740
rect 860 6680 920 6700
rect 970 6860 1030 6900
rect 1550 6860 1610 6900
rect 970 6840 1110 6860
rect 970 6800 980 6840
rect 1020 6800 1060 6840
rect 1100 6800 1110 6840
rect 970 6740 1110 6800
rect 970 6700 980 6740
rect 1020 6700 1060 6740
rect 1100 6700 1110 6740
rect 970 6680 1110 6700
rect 1470 6840 1610 6860
rect 1470 6800 1480 6840
rect 1520 6800 1560 6840
rect 1600 6800 1610 6840
rect 1470 6740 1610 6800
rect 1470 6700 1480 6740
rect 1520 6700 1560 6740
rect 1600 6700 1610 6740
rect 1470 6680 1610 6700
rect 1660 6840 1720 7020
rect 1760 6970 1840 6980
rect 1760 6910 1770 6970
rect 1830 6910 1840 6970
rect 1760 6900 1840 6910
rect 1660 6800 1670 6840
rect 1710 6800 1720 6840
rect 1660 6740 1720 6800
rect 1660 6700 1670 6740
rect 1710 6700 1720 6740
rect 1660 6680 1720 6700
rect 1770 6840 1830 6900
rect 1770 6800 1780 6840
rect 1820 6800 1830 6840
rect 1770 6740 1830 6800
rect 1770 6700 1780 6740
rect 1820 6700 1830 6740
rect 1770 6680 1830 6700
rect 1880 6840 1940 7020
rect 1980 6970 2060 6980
rect 1980 6910 1990 6970
rect 2050 6910 2060 6970
rect 1980 6900 2060 6910
rect 1880 6800 1890 6840
rect 1930 6800 1940 6840
rect 1880 6740 1940 6800
rect 1880 6700 1890 6740
rect 1930 6700 1940 6740
rect 1880 6680 1940 6700
rect 1990 6840 2050 6900
rect 1990 6800 2000 6840
rect 2040 6800 2050 6840
rect 1990 6740 2050 6800
rect 1990 6700 2000 6740
rect 2040 6700 2050 6740
rect 1990 6680 2050 6700
rect 2100 6840 2160 7020
rect 2200 6970 2280 6980
rect 2200 6910 2210 6970
rect 2270 6910 2280 6970
rect 2200 6900 2280 6910
rect 2100 6800 2110 6840
rect 2150 6800 2160 6840
rect 2100 6740 2160 6800
rect 2100 6700 2110 6740
rect 2150 6700 2160 6740
rect 2100 6680 2160 6700
rect 2210 6840 2270 6900
rect 2210 6800 2220 6840
rect 2260 6800 2270 6840
rect 2210 6740 2270 6800
rect 2210 6700 2220 6740
rect 2260 6700 2270 6740
rect 2210 6680 2270 6700
rect 2320 6840 2380 7020
rect 2420 6970 2500 6980
rect 2420 6910 2430 6970
rect 2490 6910 2500 6970
rect 2420 6900 2500 6910
rect 2320 6800 2330 6840
rect 2370 6800 2380 6840
rect 2320 6740 2380 6800
rect 2320 6700 2330 6740
rect 2370 6700 2380 6740
rect 2320 6680 2380 6700
rect 2430 6840 2490 6900
rect 2430 6800 2440 6840
rect 2480 6800 2490 6840
rect 2430 6740 2490 6800
rect 2430 6700 2440 6740
rect 2480 6700 2490 6740
rect 2430 6680 2490 6700
rect 2540 6840 2600 7020
rect 2640 6970 2720 6980
rect 2640 6910 2650 6970
rect 2710 6910 2720 6970
rect 2640 6900 2720 6910
rect 2540 6800 2550 6840
rect 2590 6800 2600 6840
rect 2540 6740 2600 6800
rect 2540 6700 2550 6740
rect 2590 6700 2600 6740
rect 2540 6680 2600 6700
rect 2650 6840 2710 6900
rect 2650 6800 2660 6840
rect 2700 6800 2710 6840
rect 2650 6740 2710 6800
rect 2650 6700 2660 6740
rect 2700 6700 2710 6740
rect 2650 6680 2710 6700
rect 2760 6840 2820 7020
rect 2860 6970 2940 6980
rect 2860 6910 2870 6970
rect 2930 6910 2940 6970
rect 2860 6900 2940 6910
rect 2760 6800 2770 6840
rect 2810 6800 2820 6840
rect 2760 6740 2820 6800
rect 2760 6700 2770 6740
rect 2810 6700 2820 6740
rect 2760 6680 2820 6700
rect 2870 6860 2930 6900
rect 2870 6840 3010 6860
rect 2870 6800 2880 6840
rect 2920 6800 2960 6840
rect 3000 6800 3010 6840
rect 2870 6740 3010 6800
rect 2870 6700 2880 6740
rect 2920 6700 2960 6740
rect 3000 6700 3010 6740
rect 2870 6680 3010 6700
rect -184 6632 -126 6640
rect -184 6580 -182 6632
rect -130 6580 -126 6632
rect -184 6570 -126 6580
rect -74 6632 -16 6640
rect -74 6580 -72 6632
rect -20 6580 -16 6632
rect -74 6570 -16 6580
rect 36 6632 94 6640
rect 36 6580 38 6632
rect 90 6580 94 6632
rect 36 6570 94 6580
rect 146 6632 204 6640
rect 146 6580 148 6632
rect 200 6580 204 6632
rect 146 6570 204 6580
rect 256 6632 314 6640
rect 256 6580 258 6632
rect 310 6580 314 6632
rect 256 6570 314 6580
rect 366 6632 424 6640
rect 366 6580 368 6632
rect 420 6580 424 6632
rect 366 6570 424 6580
rect 476 6632 534 6640
rect 476 6580 478 6632
rect 530 6580 534 6632
rect 476 6570 534 6580
rect 586 6632 644 6640
rect 586 6580 588 6632
rect 640 6580 644 6632
rect 586 6570 644 6580
rect 696 6632 754 6640
rect 696 6580 698 6632
rect 750 6580 754 6632
rect 696 6570 754 6580
rect 806 6632 864 6640
rect 806 6580 808 6632
rect 860 6580 864 6632
rect 806 6570 864 6580
rect 1716 6632 1774 6640
rect 1716 6580 1718 6632
rect 1770 6580 1774 6632
rect 1716 6570 1774 6580
rect 1826 6632 1884 6640
rect 1826 6580 1828 6632
rect 1880 6580 1884 6632
rect 1826 6570 1884 6580
rect 1936 6632 1994 6640
rect 1936 6580 1938 6632
rect 1990 6580 1994 6632
rect 1936 6570 1994 6580
rect 2046 6632 2104 6640
rect 2046 6580 2048 6632
rect 2100 6580 2104 6632
rect 2046 6570 2104 6580
rect 2156 6632 2214 6640
rect 2156 6580 2158 6632
rect 2210 6580 2214 6632
rect 2156 6570 2214 6580
rect 2266 6632 2324 6640
rect 2266 6580 2268 6632
rect 2320 6580 2324 6632
rect 2266 6570 2324 6580
rect 2376 6632 2434 6640
rect 2376 6580 2378 6632
rect 2430 6580 2434 6632
rect 2376 6570 2434 6580
rect 2486 6632 2544 6640
rect 2486 6580 2488 6632
rect 2540 6580 2544 6632
rect 2486 6570 2544 6580
rect 2596 6632 2654 6640
rect 2596 6580 2598 6632
rect 2650 6580 2654 6632
rect 2596 6570 2654 6580
rect 2706 6632 2764 6640
rect 2706 6580 2708 6632
rect 2760 6580 2764 6632
rect 2706 6570 2764 6580
rect -370 6530 -290 6540
rect -370 6470 -360 6530
rect -300 6470 -290 6530
rect -370 6450 -290 6470
rect -370 6390 -360 6450
rect -300 6390 -290 6450
rect -370 6370 -290 6390
rect -370 6310 -360 6370
rect -300 6310 -290 6370
rect -370 6300 -290 6310
rect -10 6530 70 6540
rect -10 6470 0 6530
rect 60 6470 70 6530
rect -10 6450 70 6470
rect -10 6390 0 6450
rect 60 6390 70 6450
rect -10 6370 70 6390
rect -10 6310 0 6370
rect 60 6310 70 6370
rect -10 6300 70 6310
rect 350 6530 430 6540
rect 350 6470 360 6530
rect 420 6470 430 6530
rect 350 6450 430 6470
rect 350 6390 360 6450
rect 420 6390 430 6450
rect 350 6370 430 6390
rect 350 6310 360 6370
rect 420 6310 430 6370
rect 350 6300 430 6310
rect 710 6530 790 6540
rect 710 6470 720 6530
rect 780 6470 790 6530
rect 710 6450 790 6470
rect 710 6390 720 6450
rect 780 6390 790 6450
rect 710 6370 790 6390
rect 710 6310 720 6370
rect 780 6310 790 6370
rect 710 6300 790 6310
rect 1070 6530 1150 6540
rect 1070 6470 1080 6530
rect 1140 6470 1150 6530
rect 1070 6450 1150 6470
rect 1070 6390 1080 6450
rect 1140 6390 1150 6450
rect 1070 6370 1150 6390
rect 1070 6310 1080 6370
rect 1140 6310 1150 6370
rect 1070 6300 1150 6310
rect 1430 6530 1510 6540
rect 1430 6470 1440 6530
rect 1500 6470 1510 6530
rect 1430 6450 1510 6470
rect 1430 6390 1440 6450
rect 1500 6390 1510 6450
rect 1430 6370 1510 6390
rect 1430 6310 1440 6370
rect 1500 6310 1510 6370
rect 1430 6300 1510 6310
rect 1790 6530 1870 6540
rect 1790 6470 1800 6530
rect 1860 6470 1870 6530
rect 1790 6450 1870 6470
rect 1790 6390 1800 6450
rect 1860 6390 1870 6450
rect 1790 6370 1870 6390
rect 1790 6310 1800 6370
rect 1860 6310 1870 6370
rect 1790 6300 1870 6310
rect 2150 6530 2230 6540
rect 2150 6470 2160 6530
rect 2220 6470 2230 6530
rect 2150 6450 2230 6470
rect 2150 6390 2160 6450
rect 2220 6390 2230 6450
rect 2150 6370 2230 6390
rect 2150 6310 2160 6370
rect 2220 6310 2230 6370
rect 2150 6300 2230 6310
rect 2510 6530 2590 6540
rect 2510 6470 2520 6530
rect 2580 6470 2590 6530
rect 2510 6450 2590 6470
rect 2510 6390 2520 6450
rect 2580 6390 2590 6450
rect 2510 6370 2590 6390
rect 2510 6310 2520 6370
rect 2580 6310 2590 6370
rect 2510 6300 2590 6310
rect 2870 6530 2950 6540
rect 2870 6470 2880 6530
rect 2940 6470 2950 6530
rect 2870 6450 2950 6470
rect 2870 6390 2880 6450
rect 2940 6390 2950 6450
rect 2870 6370 2950 6390
rect 2870 6310 2880 6370
rect 2940 6310 2950 6370
rect 2870 6300 2950 6310
rect 3500 6530 3580 6540
rect 3500 6470 3510 6530
rect 3570 6470 3580 6530
rect 3500 6450 3580 6470
rect 3500 6390 3510 6450
rect 3570 6390 3580 6450
rect 3500 6370 3580 6390
rect 3500 6310 3510 6370
rect 3570 6310 3580 6370
rect 3500 6300 3580 6310
rect 3940 6530 4020 6540
rect 3940 6470 3950 6530
rect 4010 6470 4020 6530
rect 3940 6450 4020 6470
rect 3940 6390 3950 6450
rect 4010 6390 4020 6450
rect 3940 6370 4020 6390
rect 3940 6310 3950 6370
rect 4010 6310 4020 6370
rect 3940 6300 4020 6310
rect -360 6240 -300 6260
rect -360 6200 -350 6240
rect -310 6200 -300 6240
rect -360 6140 -300 6200
rect -360 6100 -350 6140
rect -310 6100 -300 6140
rect -360 6040 -300 6100
rect -360 6000 -350 6040
rect -310 6000 -300 6040
rect -360 5940 -300 6000
rect -360 5900 -350 5940
rect -310 5900 -300 5940
rect -360 5840 -300 5900
rect -360 5800 -350 5840
rect -310 5800 -300 5840
rect -360 5740 -300 5800
rect -360 5700 -350 5740
rect -310 5700 -300 5740
rect -360 5680 -300 5700
rect -180 6240 -120 6260
rect -180 6200 -170 6240
rect -130 6200 -120 6240
rect -180 6140 -120 6200
rect -180 6100 -170 6140
rect -130 6100 -120 6140
rect -180 6040 -120 6100
rect -180 6000 -170 6040
rect -130 6000 -120 6040
rect -180 5940 -120 6000
rect -180 5900 -170 5940
rect -130 5900 -120 5940
rect -180 5840 -120 5900
rect -180 5800 -170 5840
rect -130 5800 -120 5840
rect -180 5740 -120 5800
rect -180 5700 -170 5740
rect -130 5700 -120 5740
rect -180 5200 -120 5700
rect 0 6240 60 6260
rect 0 6200 10 6240
rect 50 6200 60 6240
rect 0 6140 60 6200
rect 0 6100 10 6140
rect 50 6100 60 6140
rect 0 6040 60 6100
rect 0 6000 10 6040
rect 50 6000 60 6040
rect 0 5940 60 6000
rect 0 5900 10 5940
rect 50 5900 60 5940
rect 0 5840 60 5900
rect 0 5800 10 5840
rect 50 5800 60 5840
rect 0 5740 60 5800
rect 0 5700 10 5740
rect 50 5700 60 5740
rect 0 5680 60 5700
rect 180 6240 240 6260
rect 180 6200 190 6240
rect 230 6200 240 6240
rect 180 6140 240 6200
rect 180 6100 190 6140
rect 230 6100 240 6140
rect 180 6040 240 6100
rect 180 6000 190 6040
rect 230 6000 240 6040
rect 180 5940 240 6000
rect 180 5900 190 5940
rect 230 5900 240 5940
rect 180 5840 240 5900
rect 180 5800 190 5840
rect 230 5800 240 5840
rect 180 5740 240 5800
rect 180 5700 190 5740
rect 230 5700 240 5740
rect 180 5680 240 5700
rect 360 6240 420 6260
rect 360 6200 370 6240
rect 410 6200 420 6240
rect 360 6140 420 6200
rect 360 6100 370 6140
rect 410 6100 420 6140
rect 360 6040 420 6100
rect 360 6000 370 6040
rect 410 6000 420 6040
rect 360 5940 420 6000
rect 360 5900 370 5940
rect 410 5900 420 5940
rect 360 5840 420 5900
rect 360 5800 370 5840
rect 410 5800 420 5840
rect 360 5740 420 5800
rect 360 5700 370 5740
rect 410 5700 420 5740
rect 360 5680 420 5700
rect 540 6240 600 6260
rect 540 6200 550 6240
rect 590 6200 600 6240
rect 540 6140 600 6200
rect 540 6100 550 6140
rect 590 6100 600 6140
rect 540 6040 600 6100
rect 540 6000 550 6040
rect 590 6000 600 6040
rect 540 5940 600 6000
rect 540 5900 550 5940
rect 590 5900 600 5940
rect 540 5840 600 5900
rect 540 5800 550 5840
rect 590 5800 600 5840
rect 540 5740 600 5800
rect 540 5700 550 5740
rect 590 5700 600 5740
rect 540 5680 600 5700
rect 720 6240 780 6260
rect 720 6200 730 6240
rect 770 6200 780 6240
rect 720 6140 780 6200
rect 720 6100 730 6140
rect 770 6100 780 6140
rect 720 6040 780 6100
rect 720 6000 730 6040
rect 770 6000 780 6040
rect 720 5940 780 6000
rect 720 5900 730 5940
rect 770 5900 780 5940
rect 720 5840 780 5900
rect 720 5800 730 5840
rect 770 5800 780 5840
rect 720 5740 780 5800
rect 720 5700 730 5740
rect 770 5700 780 5740
rect 720 5680 780 5700
rect 900 6240 960 6260
rect 900 6200 910 6240
rect 950 6200 960 6240
rect 900 6140 960 6200
rect 900 6100 910 6140
rect 950 6100 960 6140
rect 900 6040 960 6100
rect 900 6000 910 6040
rect 950 6000 960 6040
rect 900 5940 960 6000
rect 900 5900 910 5940
rect 950 5900 960 5940
rect 900 5840 960 5900
rect 900 5800 910 5840
rect 950 5800 960 5840
rect 900 5740 960 5800
rect 900 5700 910 5740
rect 950 5700 960 5740
rect 900 5680 960 5700
rect 1080 6240 1140 6260
rect 1080 6200 1090 6240
rect 1130 6200 1140 6240
rect 1080 6140 1140 6200
rect 1080 6100 1090 6140
rect 1130 6100 1140 6140
rect 1080 6040 1140 6100
rect 1080 6000 1090 6040
rect 1130 6000 1140 6040
rect 1080 5940 1140 6000
rect 1080 5900 1090 5940
rect 1130 5900 1140 5940
rect 1080 5840 1140 5900
rect 1080 5800 1090 5840
rect 1130 5800 1140 5840
rect 1080 5740 1140 5800
rect 1080 5700 1090 5740
rect 1130 5700 1140 5740
rect 1080 5680 1140 5700
rect 1260 6240 1320 6260
rect 1260 6200 1270 6240
rect 1310 6200 1320 6240
rect 1260 6140 1320 6200
rect 1260 6100 1270 6140
rect 1310 6100 1320 6140
rect 1260 6040 1320 6100
rect 1260 6000 1270 6040
rect 1310 6000 1320 6040
rect 1260 5940 1320 6000
rect 1260 5900 1270 5940
rect 1310 5900 1320 5940
rect 1260 5840 1320 5900
rect 1260 5800 1270 5840
rect 1310 5800 1320 5840
rect 1260 5740 1320 5800
rect 1260 5700 1270 5740
rect 1310 5700 1320 5740
rect -90 5630 -20 5640
rect -30 5570 -20 5630
rect -90 5560 -20 5570
rect 80 5630 160 5640
rect 80 5570 90 5630
rect 150 5570 160 5630
rect 80 5560 160 5570
rect 190 5310 230 5680
rect 260 5630 340 5640
rect 260 5570 270 5630
rect 330 5570 340 5630
rect 260 5560 340 5570
rect 440 5630 520 5640
rect 440 5570 450 5630
rect 510 5570 520 5630
rect 440 5560 520 5570
rect 550 5420 590 5680
rect 620 5630 700 5640
rect 620 5570 630 5630
rect 690 5570 700 5630
rect 620 5560 700 5570
rect 800 5630 880 5640
rect 800 5570 810 5630
rect 870 5570 880 5630
rect 800 5560 880 5570
rect 910 5530 950 5680
rect 980 5630 1060 5640
rect 980 5570 990 5630
rect 1050 5570 1060 5630
rect 980 5560 1060 5570
rect 1160 5630 1230 5640
rect 1160 5570 1170 5630
rect 1160 5560 1230 5570
rect 890 5520 970 5530
rect 890 5460 900 5520
rect 960 5460 970 5520
rect 890 5450 970 5460
rect 530 5410 610 5420
rect 530 5350 540 5410
rect 600 5350 610 5410
rect 530 5340 610 5350
rect 170 5300 250 5310
rect 170 5240 180 5300
rect 240 5240 250 5300
rect 170 5230 250 5240
rect 1260 5200 1320 5700
rect 1440 6240 1500 6260
rect 1440 6200 1450 6240
rect 1490 6200 1500 6240
rect 1440 6140 1500 6200
rect 1440 6100 1450 6140
rect 1490 6100 1500 6140
rect 1440 6040 1500 6100
rect 1440 6000 1450 6040
rect 1490 6000 1500 6040
rect 1440 5940 1500 6000
rect 1440 5900 1450 5940
rect 1490 5900 1500 5940
rect 1440 5840 1500 5900
rect 1440 5800 1450 5840
rect 1490 5800 1500 5840
rect 1440 5740 1500 5800
rect 1440 5700 1450 5740
rect 1490 5700 1500 5740
rect 1440 5680 1500 5700
rect 1620 6240 1680 6260
rect 1620 6200 1630 6240
rect 1670 6200 1680 6240
rect 1620 6140 1680 6200
rect 1620 6100 1630 6140
rect 1670 6100 1680 6140
rect 1620 6040 1680 6100
rect 1620 6000 1630 6040
rect 1670 6000 1680 6040
rect 1620 5940 1680 6000
rect 1620 5900 1630 5940
rect 1670 5900 1680 5940
rect 1620 5840 1680 5900
rect 1620 5800 1630 5840
rect 1670 5800 1680 5840
rect 1620 5740 1680 5800
rect 1620 5700 1630 5740
rect 1670 5700 1680 5740
rect 1620 5680 1680 5700
rect 1800 6240 1860 6260
rect 1800 6200 1810 6240
rect 1850 6200 1860 6240
rect 1800 6140 1860 6200
rect 1800 6100 1810 6140
rect 1850 6100 1860 6140
rect 1800 6040 1860 6100
rect 1800 6000 1810 6040
rect 1850 6000 1860 6040
rect 1800 5940 1860 6000
rect 1800 5900 1810 5940
rect 1850 5900 1860 5940
rect 1800 5840 1860 5900
rect 1800 5800 1810 5840
rect 1850 5800 1860 5840
rect 1800 5740 1860 5800
rect 1800 5700 1810 5740
rect 1850 5700 1860 5740
rect 1800 5680 1860 5700
rect 1980 6240 2040 6260
rect 1980 6200 1990 6240
rect 2030 6200 2040 6240
rect 1980 6140 2040 6200
rect 1980 6100 1990 6140
rect 2030 6100 2040 6140
rect 1980 6040 2040 6100
rect 1980 6000 1990 6040
rect 2030 6000 2040 6040
rect 1980 5940 2040 6000
rect 1980 5900 1990 5940
rect 2030 5900 2040 5940
rect 1980 5840 2040 5900
rect 1980 5800 1990 5840
rect 2030 5800 2040 5840
rect 1980 5740 2040 5800
rect 1980 5700 1990 5740
rect 2030 5700 2040 5740
rect 1980 5680 2040 5700
rect 2160 6240 2220 6260
rect 2160 6200 2170 6240
rect 2210 6200 2220 6240
rect 2160 6140 2220 6200
rect 2160 6100 2170 6140
rect 2210 6100 2220 6140
rect 2160 6040 2220 6100
rect 2160 6000 2170 6040
rect 2210 6000 2220 6040
rect 2160 5940 2220 6000
rect 2160 5900 2170 5940
rect 2210 5900 2220 5940
rect 2160 5840 2220 5900
rect 2160 5800 2170 5840
rect 2210 5800 2220 5840
rect 2160 5740 2220 5800
rect 2160 5700 2170 5740
rect 2210 5700 2220 5740
rect 2160 5680 2220 5700
rect 2340 6240 2400 6260
rect 2340 6200 2350 6240
rect 2390 6200 2400 6240
rect 2340 6140 2400 6200
rect 2340 6100 2350 6140
rect 2390 6100 2400 6140
rect 2340 6040 2400 6100
rect 2340 6000 2350 6040
rect 2390 6000 2400 6040
rect 2340 5940 2400 6000
rect 2340 5900 2350 5940
rect 2390 5900 2400 5940
rect 2340 5840 2400 5900
rect 2340 5800 2350 5840
rect 2390 5800 2400 5840
rect 2340 5740 2400 5800
rect 2340 5700 2350 5740
rect 2390 5700 2400 5740
rect 2340 5680 2400 5700
rect 2520 6240 2580 6260
rect 2520 6200 2530 6240
rect 2570 6200 2580 6240
rect 2520 6140 2580 6200
rect 2520 6100 2530 6140
rect 2570 6100 2580 6140
rect 2520 6040 2580 6100
rect 2520 6000 2530 6040
rect 2570 6000 2580 6040
rect 2520 5940 2580 6000
rect 2520 5900 2530 5940
rect 2570 5900 2580 5940
rect 2520 5840 2580 5900
rect 2520 5800 2530 5840
rect 2570 5800 2580 5840
rect 2520 5740 2580 5800
rect 2520 5700 2530 5740
rect 2570 5700 2580 5740
rect 2520 5680 2580 5700
rect 2700 6240 2760 6260
rect 2700 6200 2710 6240
rect 2750 6200 2760 6240
rect 2700 6140 2760 6200
rect 2700 6100 2710 6140
rect 2750 6100 2760 6140
rect 2700 6040 2760 6100
rect 2700 6000 2710 6040
rect 2750 6000 2760 6040
rect 2700 5940 2760 6000
rect 2700 5900 2710 5940
rect 2750 5900 2760 5940
rect 2700 5840 2760 5900
rect 2700 5800 2710 5840
rect 2750 5800 2760 5840
rect 2700 5740 2760 5800
rect 2700 5700 2710 5740
rect 2750 5700 2760 5740
rect 1350 5630 1600 5640
rect 1410 5570 1440 5630
rect 1500 5570 1530 5630
rect 1590 5570 1600 5630
rect 1350 5560 1600 5570
rect -190 5190 -110 5200
rect -190 5130 -180 5190
rect -120 5130 -110 5190
rect -190 5120 -110 5130
rect 1250 5190 1330 5200
rect 1250 5130 1260 5190
rect 1320 5130 1330 5190
rect 1250 5120 1330 5130
rect -1470 5080 -1390 5090
rect -1470 5020 -1460 5080
rect -1400 5020 -1390 5080
rect -1470 5000 -1390 5020
rect -1470 4940 -1460 5000
rect -1400 4940 -1390 5000
rect -1470 4920 -1390 4940
rect -1470 4860 -1460 4920
rect -1400 4860 -1390 4920
rect -1470 4850 -1390 4860
rect -1230 5080 -1150 5090
rect -1230 5020 -1220 5080
rect -1160 5020 -1150 5080
rect -1230 5000 -1150 5020
rect -1230 4940 -1220 5000
rect -1160 4940 -1150 5000
rect -1230 4920 -1150 4940
rect -1230 4860 -1220 4920
rect -1160 4860 -1150 4920
rect -1230 4850 -1150 4860
rect -990 5080 -910 5090
rect -990 5020 -980 5080
rect -920 5020 -910 5080
rect -990 5000 -910 5020
rect -990 4940 -980 5000
rect -920 4940 -910 5000
rect -990 4920 -910 4940
rect -990 4860 -980 4920
rect -920 4860 -910 4920
rect -990 4850 -910 4860
rect -750 5080 -670 5090
rect -750 5020 -740 5080
rect -680 5020 -670 5080
rect -750 5000 -670 5020
rect -750 4940 -740 5000
rect -680 4940 -670 5000
rect -750 4920 -670 4940
rect -750 4860 -740 4920
rect -680 4860 -670 4920
rect -750 4850 -670 4860
rect -510 5080 -430 5090
rect -510 5020 -500 5080
rect -440 5020 -430 5080
rect -510 5000 -430 5020
rect -510 4940 -500 5000
rect -440 4940 -430 5000
rect -510 4920 -430 4940
rect -510 4860 -500 4920
rect -440 4860 -430 4920
rect -510 4850 -430 4860
rect -270 5080 -190 5090
rect -270 5020 -260 5080
rect -200 5020 -190 5080
rect -270 5000 -190 5020
rect -270 4940 -260 5000
rect -200 4940 -190 5000
rect -270 4920 -190 4940
rect -270 4860 -260 4920
rect -200 4860 -190 4920
rect -270 4850 -190 4860
rect -30 5080 50 5090
rect -30 5020 -20 5080
rect 40 5020 50 5080
rect -30 5000 50 5020
rect -30 4940 -20 5000
rect 40 4940 50 5000
rect -30 4920 50 4940
rect -30 4860 -20 4920
rect 40 4860 50 4920
rect -30 4850 50 4860
rect 210 5080 290 5090
rect 210 5020 220 5080
rect 280 5020 290 5080
rect 210 5000 290 5020
rect 210 4940 220 5000
rect 280 4940 290 5000
rect 210 4920 290 4940
rect 210 4860 220 4920
rect 280 4860 290 4920
rect 210 4850 290 4860
rect 450 5080 530 5090
rect 450 5020 460 5080
rect 520 5020 530 5080
rect 450 5000 530 5020
rect 450 4940 460 5000
rect 520 4940 530 5000
rect 450 4920 530 4940
rect 450 4860 460 4920
rect 520 4860 530 4920
rect 450 4850 530 4860
rect 690 5080 770 5090
rect 690 5020 700 5080
rect 760 5020 770 5080
rect 690 5000 770 5020
rect 690 4940 700 5000
rect 760 4940 770 5000
rect 690 4920 770 4940
rect 690 4860 700 4920
rect 760 4860 770 4920
rect 690 4850 770 4860
rect 930 5080 1010 5090
rect 930 5020 940 5080
rect 1000 5020 1010 5080
rect 930 5000 1010 5020
rect 930 4940 940 5000
rect 1000 4940 1010 5000
rect 930 4920 1010 4940
rect 930 4860 940 4920
rect 1000 4860 1010 4920
rect 930 4850 1010 4860
rect -1460 4800 -1400 4850
rect -1460 4760 -1450 4800
rect -1410 4760 -1400 4800
rect -1460 4680 -1400 4760
rect -1350 4810 -1270 4820
rect -1350 4750 -1340 4810
rect -1280 4750 -1270 4810
rect -1350 4740 -1270 4750
rect -1460 4640 -1450 4680
rect -1410 4640 -1400 4680
rect -1460 4580 -1400 4640
rect -1460 4540 -1450 4580
rect -1410 4540 -1400 4580
rect -1460 4520 -1400 4540
rect -1340 4680 -1280 4740
rect -1340 4640 -1330 4680
rect -1290 4640 -1280 4680
rect -1340 4580 -1280 4640
rect -1340 4540 -1330 4580
rect -1290 4540 -1280 4580
rect -1340 4520 -1280 4540
rect -1220 4680 -1160 4850
rect -1220 4640 -1210 4680
rect -1170 4640 -1160 4680
rect -1220 4580 -1160 4640
rect -1220 4540 -1210 4580
rect -1170 4540 -1160 4580
rect -1220 4520 -1160 4540
rect -1100 4680 -1040 4700
rect -1100 4640 -1090 4680
rect -1050 4640 -1040 4680
rect -1100 4580 -1040 4640
rect -1100 4540 -1090 4580
rect -1050 4540 -1040 4580
rect -1100 4480 -1040 4540
rect -980 4680 -920 4850
rect -980 4640 -970 4680
rect -930 4640 -920 4680
rect -980 4580 -920 4640
rect -980 4540 -970 4580
rect -930 4540 -920 4580
rect -980 4520 -920 4540
rect -860 4680 -800 4700
rect -860 4640 -850 4680
rect -810 4640 -800 4680
rect -860 4580 -800 4640
rect -860 4540 -850 4580
rect -810 4540 -800 4580
rect -1110 4470 -1030 4480
rect -1280 4450 -1220 4470
rect -1280 4410 -1270 4450
rect -1230 4410 -1220 4450
rect -1280 4360 -1220 4410
rect -1110 4410 -1100 4470
rect -1040 4410 -1030 4470
rect -1110 4400 -1030 4410
rect -860 4360 -800 4540
rect -740 4680 -680 4850
rect -630 4810 -550 4820
rect -630 4750 -620 4810
rect -560 4750 -550 4810
rect -630 4740 -550 4750
rect -740 4640 -730 4680
rect -690 4640 -680 4680
rect -740 4580 -680 4640
rect -740 4540 -730 4580
rect -690 4540 -680 4580
rect -740 4520 -680 4540
rect -620 4680 -560 4740
rect -620 4640 -610 4680
rect -570 4640 -560 4680
rect -620 4580 -560 4640
rect -620 4540 -610 4580
rect -570 4540 -560 4580
rect -620 4520 -560 4540
rect -500 4680 -440 4850
rect -500 4640 -490 4680
rect -450 4640 -440 4680
rect -500 4580 -440 4640
rect -500 4540 -490 4580
rect -450 4540 -440 4580
rect -500 4520 -440 4540
rect -380 4680 -320 4700
rect -380 4640 -370 4680
rect -330 4640 -320 4680
rect -380 4580 -320 4640
rect -380 4540 -370 4580
rect -330 4540 -320 4580
rect -380 4480 -320 4540
rect -260 4680 -200 4850
rect -260 4640 -250 4680
rect -210 4640 -200 4680
rect -260 4580 -200 4640
rect -260 4540 -250 4580
rect -210 4540 -200 4580
rect -260 4520 -200 4540
rect -140 4680 -80 4700
rect -140 4640 -130 4680
rect -90 4640 -80 4680
rect -140 4580 -80 4640
rect -140 4540 -130 4580
rect -90 4540 -80 4580
rect -620 4460 -560 4480
rect -620 4420 -610 4460
rect -570 4420 -560 4460
rect -620 4360 -560 4420
rect -390 4470 -310 4480
rect -390 4410 -380 4470
rect -320 4410 -310 4470
rect -2310 3580 -2300 3640
rect -2240 3580 -2230 3640
rect -2310 1900 -2230 3580
rect -1370 4350 -1210 4360
rect -1370 4290 -1360 4350
rect -1300 4290 -1280 4350
rect -1220 4290 -1210 4350
rect -1370 4280 -1210 4290
rect -870 4350 -790 4360
rect -870 4290 -860 4350
rect -800 4290 -790 4350
rect -870 4280 -790 4290
rect -630 4350 -550 4360
rect -630 4290 -620 4350
rect -560 4290 -550 4350
rect -1370 2010 -1290 4280
rect -630 4080 -550 4290
rect -630 4020 -620 4080
rect -560 4020 -550 4080
rect -630 4010 -550 4020
rect -620 3740 -560 4010
rect -390 3970 -310 4410
rect -140 4360 -80 4540
rect -20 4680 40 4850
rect 90 4810 170 4820
rect 90 4750 100 4810
rect 160 4750 170 4810
rect 90 4740 170 4750
rect -20 4640 -10 4680
rect 30 4640 40 4680
rect -20 4580 40 4640
rect -20 4540 -10 4580
rect 30 4540 40 4580
rect -20 4520 40 4540
rect 100 4680 160 4740
rect 100 4640 110 4680
rect 150 4640 160 4680
rect 100 4580 160 4640
rect 100 4540 110 4580
rect 150 4540 160 4580
rect 100 4520 160 4540
rect 220 4680 280 4850
rect 220 4640 230 4680
rect 270 4640 280 4680
rect 220 4580 280 4640
rect 220 4540 230 4580
rect 270 4540 280 4580
rect 220 4520 280 4540
rect 340 4680 400 4700
rect 340 4640 350 4680
rect 390 4640 400 4680
rect 340 4580 400 4640
rect 340 4540 350 4580
rect 390 4540 400 4580
rect 340 4480 400 4540
rect 460 4680 520 4850
rect 460 4640 470 4680
rect 510 4640 520 4680
rect 460 4580 520 4640
rect 460 4540 470 4580
rect 510 4540 520 4580
rect 460 4520 520 4540
rect 580 4680 640 4700
rect 580 4640 590 4680
rect 630 4640 640 4680
rect 580 4580 640 4640
rect 580 4540 590 4580
rect 630 4540 640 4580
rect 100 4460 160 4480
rect 100 4420 110 4460
rect 150 4420 160 4460
rect 100 4360 160 4420
rect 330 4470 410 4480
rect 330 4410 340 4470
rect 400 4410 410 4470
rect 330 4400 410 4410
rect 580 4360 640 4540
rect 700 4680 760 4850
rect 810 4810 890 4820
rect 810 4750 820 4810
rect 880 4750 890 4810
rect 810 4740 890 4750
rect 940 4800 1000 4850
rect 940 4760 950 4800
rect 990 4760 1000 4800
rect 700 4640 710 4680
rect 750 4640 760 4680
rect 700 4580 760 4640
rect 700 4540 710 4580
rect 750 4540 760 4580
rect 700 4520 760 4540
rect 820 4680 880 4740
rect 820 4640 830 4680
rect 870 4640 880 4680
rect 820 4580 880 4640
rect 820 4540 830 4580
rect 870 4540 880 4580
rect 820 4520 880 4540
rect 940 4680 1000 4760
rect 1070 4810 1150 4820
rect 1070 4750 1080 4810
rect 1140 4750 1150 4810
rect 1070 4740 1150 4750
rect 1430 4810 1510 5560
rect 1630 5530 1670 5680
rect 1700 5630 1780 5640
rect 1700 5570 1710 5630
rect 1770 5570 1780 5630
rect 1700 5560 1780 5570
rect 1880 5630 1960 5640
rect 1880 5570 1890 5630
rect 1950 5570 1960 5630
rect 1880 5560 1960 5570
rect 1610 5520 1690 5530
rect 1610 5460 1620 5520
rect 1680 5460 1690 5520
rect 1610 5450 1690 5460
rect 1990 5420 2030 5680
rect 2060 5630 2140 5640
rect 2060 5570 2070 5630
rect 2130 5570 2140 5630
rect 2060 5560 2140 5570
rect 2240 5630 2320 5640
rect 2240 5570 2250 5630
rect 2310 5570 2320 5630
rect 2240 5560 2320 5570
rect 1970 5410 2050 5420
rect 1970 5350 1980 5410
rect 2040 5350 2050 5410
rect 1970 5340 2050 5350
rect 2350 5310 2390 5680
rect 2420 5630 2500 5640
rect 2420 5570 2430 5630
rect 2490 5570 2500 5630
rect 2420 5560 2500 5570
rect 2600 5630 2670 5640
rect 2600 5570 2610 5630
rect 2600 5560 2670 5570
rect 2330 5300 2410 5310
rect 2330 5240 2340 5300
rect 2400 5240 2410 5300
rect 2330 5230 2410 5240
rect 2700 5200 2760 5700
rect 2880 6240 2940 6260
rect 2880 6200 2890 6240
rect 2930 6200 2940 6240
rect 2880 6140 2940 6200
rect 3510 6180 3570 6300
rect 3950 6180 4010 6300
rect 2880 6100 2890 6140
rect 2930 6100 2940 6140
rect 3250 6170 3330 6180
rect 3250 6110 3260 6170
rect 3320 6110 3330 6170
rect 3250 6100 3330 6110
rect 3500 6160 3580 6180
rect 3500 6120 3520 6160
rect 3560 6120 3580 6160
rect 3500 6100 3580 6120
rect 3720 6170 3800 6180
rect 3720 6110 3730 6170
rect 3790 6110 3800 6170
rect 3720 6100 3800 6110
rect 3940 6160 4020 6180
rect 3940 6120 3960 6160
rect 4000 6120 4020 6160
rect 3940 6100 4020 6120
rect 2880 6040 2940 6100
rect 2880 6000 2890 6040
rect 2930 6000 2940 6040
rect 2880 5940 2940 6000
rect 2880 5900 2890 5940
rect 2930 5900 2940 5940
rect 2880 5840 2940 5900
rect 2880 5800 2890 5840
rect 2930 5800 2940 5840
rect 2880 5740 2940 5800
rect 2880 5700 2890 5740
rect 2930 5700 2940 5740
rect 2880 5680 2940 5700
rect 3270 5420 3310 6100
rect 3510 6040 3570 6100
rect 3510 6000 3520 6040
rect 3560 6000 3570 6040
rect 3510 5940 3570 6000
rect 3510 5900 3520 5940
rect 3560 5900 3570 5940
rect 3510 5880 3570 5900
rect 3620 6040 3680 6060
rect 3620 6000 3630 6040
rect 3670 6000 3680 6040
rect 3620 5940 3680 6000
rect 3620 5900 3630 5940
rect 3670 5900 3680 5940
rect 3620 5840 3680 5900
rect 3730 6040 3790 6100
rect 3730 6000 3740 6040
rect 3780 6000 3790 6040
rect 3730 5940 3790 6000
rect 3730 5900 3740 5940
rect 3780 5900 3790 5940
rect 3730 5880 3790 5900
rect 3840 6040 3900 6060
rect 3840 6000 3850 6040
rect 3890 6000 3900 6040
rect 3840 5940 3900 6000
rect 3840 5900 3850 5940
rect 3890 5900 3900 5940
rect 3840 5840 3900 5900
rect 3950 6040 4010 6100
rect 3950 6000 3960 6040
rect 4000 6000 4010 6040
rect 3950 5940 4010 6000
rect 3950 5900 3960 5940
rect 4000 5900 4010 5940
rect 3950 5880 4010 5900
rect 3600 5830 3680 5840
rect 3600 5770 3610 5830
rect 3670 5770 3680 5830
rect 3600 5760 3680 5770
rect 3720 5820 3800 5840
rect 3720 5780 3740 5820
rect 3780 5780 3800 5820
rect 3250 5410 3330 5420
rect 3250 5350 3260 5410
rect 3320 5350 3330 5410
rect 3250 5340 3330 5350
rect 3720 5300 3800 5780
rect 3840 5830 3920 5840
rect 3840 5770 3850 5830
rect 3910 5770 3920 5830
rect 3840 5760 3920 5770
rect 3720 5240 3730 5300
rect 3790 5240 3800 5300
rect 3720 5230 3800 5240
rect 2690 5190 2770 5200
rect 2690 5130 2700 5190
rect 2760 5130 2770 5190
rect 2690 5120 2770 5130
rect 1570 5080 1650 5090
rect 1570 5020 1580 5080
rect 1640 5020 1650 5080
rect 1570 5000 1650 5020
rect 1570 4940 1580 5000
rect 1640 4940 1650 5000
rect 1570 4920 1650 4940
rect 1570 4860 1580 4920
rect 1640 4860 1650 4920
rect 1570 4850 1650 4860
rect 1810 5080 1890 5090
rect 1810 5020 1820 5080
rect 1880 5020 1890 5080
rect 1810 5000 1890 5020
rect 1810 4940 1820 5000
rect 1880 4940 1890 5000
rect 1810 4920 1890 4940
rect 1810 4860 1820 4920
rect 1880 4860 1890 4920
rect 1810 4850 1890 4860
rect 2050 5080 2130 5090
rect 2050 5020 2060 5080
rect 2120 5020 2130 5080
rect 2050 5000 2130 5020
rect 2050 4940 2060 5000
rect 2120 4940 2130 5000
rect 2050 4920 2130 4940
rect 2050 4860 2060 4920
rect 2120 4860 2130 4920
rect 2050 4850 2130 4860
rect 2290 5080 2370 5090
rect 2290 5020 2300 5080
rect 2360 5020 2370 5080
rect 2290 5000 2370 5020
rect 2290 4940 2300 5000
rect 2360 4940 2370 5000
rect 2290 4920 2370 4940
rect 2290 4860 2300 4920
rect 2360 4860 2370 4920
rect 2290 4850 2370 4860
rect 2530 5080 2610 5090
rect 2530 5020 2540 5080
rect 2600 5020 2610 5080
rect 2530 5000 2610 5020
rect 2530 4940 2540 5000
rect 2600 4940 2610 5000
rect 2530 4920 2610 4940
rect 2530 4860 2540 4920
rect 2600 4860 2610 4920
rect 2530 4850 2610 4860
rect 2770 5080 2850 5090
rect 2770 5020 2780 5080
rect 2840 5020 2850 5080
rect 2770 5000 2850 5020
rect 2770 4940 2780 5000
rect 2840 4940 2850 5000
rect 2770 4920 2850 4940
rect 2770 4860 2780 4920
rect 2840 4860 2850 4920
rect 2770 4850 2850 4860
rect 3010 5080 3090 5090
rect 3010 5020 3020 5080
rect 3080 5020 3090 5080
rect 3010 5000 3090 5020
rect 3010 4940 3020 5000
rect 3080 4940 3090 5000
rect 3010 4920 3090 4940
rect 3010 4860 3020 4920
rect 3080 4860 3090 4920
rect 3010 4850 3090 4860
rect 3250 5080 3330 5090
rect 3250 5020 3260 5080
rect 3320 5020 3330 5080
rect 3250 5000 3330 5020
rect 3250 4940 3260 5000
rect 3320 4940 3330 5000
rect 3250 4920 3330 4940
rect 3250 4860 3260 4920
rect 3320 4860 3330 4920
rect 3250 4850 3330 4860
rect 3490 5080 3570 5090
rect 3490 5020 3500 5080
rect 3560 5020 3570 5080
rect 3490 5000 3570 5020
rect 3490 4940 3500 5000
rect 3560 4940 3570 5000
rect 3490 4920 3570 4940
rect 3490 4860 3500 4920
rect 3560 4860 3570 4920
rect 3490 4850 3570 4860
rect 3730 5080 3810 5090
rect 3730 5020 3740 5080
rect 3800 5020 3810 5080
rect 3730 5000 3810 5020
rect 3730 4940 3740 5000
rect 3800 4940 3810 5000
rect 3730 4920 3810 4940
rect 3730 4860 3740 4920
rect 3800 4860 3810 4920
rect 3730 4850 3810 4860
rect 1430 4750 1440 4810
rect 1500 4750 1510 4810
rect 1430 4740 1510 4750
rect 1580 4800 1640 4850
rect 1580 4760 1590 4800
rect 1630 4760 1640 4800
rect 940 4640 950 4680
rect 990 4640 1000 4680
rect 940 4580 1000 4640
rect 940 4540 950 4580
rect 990 4540 1000 4580
rect 940 4520 1000 4540
rect 760 4460 820 4480
rect 760 4420 770 4460
rect 810 4420 820 4460
rect 760 4360 820 4420
rect -150 4350 -70 4360
rect -150 4290 -140 4350
rect -80 4290 -70 4350
rect -150 4280 -70 4290
rect 90 4350 170 4360
rect 90 4290 100 4350
rect 160 4290 170 4350
rect 90 4280 170 4290
rect 570 4350 650 4360
rect 570 4290 580 4350
rect 640 4290 650 4350
rect 570 4280 650 4290
rect 750 4350 830 4360
rect 750 4290 760 4350
rect 820 4290 830 4350
rect 750 4280 830 4290
rect -150 4080 -70 4090
rect -150 4020 -140 4080
rect -80 4020 -70 4080
rect -150 4010 -70 4020
rect 330 4080 410 4090
rect 330 4020 340 4080
rect 400 4020 410 4080
rect 330 4010 410 4020
rect -390 3910 -380 3970
rect -320 3910 -310 3970
rect -390 3900 -310 3910
rect -458 3860 -400 3870
rect -458 3808 -454 3860
rect -402 3808 -400 3860
rect -458 3800 -400 3808
rect -370 3760 -330 3900
rect -300 3860 -242 3870
rect -300 3808 -296 3860
rect -244 3808 -242 3860
rect -300 3800 -242 3808
rect -130 3760 -90 4010
rect 90 3970 170 3980
rect 90 3910 100 3970
rect 160 3910 170 3970
rect 90 3900 170 3910
rect 24 3860 82 3870
rect 24 3808 28 3860
rect 80 3808 82 3860
rect 24 3800 82 3808
rect 110 3760 150 3900
rect 178 3860 236 3870
rect 178 3808 182 3860
rect 234 3808 236 3860
rect 178 3800 236 3808
rect 350 3760 390 4010
rect 570 3970 650 3980
rect 570 3910 580 3970
rect 640 3910 650 3970
rect 570 3900 650 3910
rect 502 3860 560 3870
rect 502 3808 506 3860
rect 558 3808 560 3860
rect 502 3800 560 3808
rect 590 3760 630 3900
rect 810 3820 890 3830
rect 810 3760 820 3820
rect 880 3760 890 3820
rect -620 3700 -610 3740
rect -570 3700 -560 3740
rect -620 3680 -560 3700
rect -500 3740 -440 3760
rect -500 3700 -490 3740
rect -450 3700 -440 3740
rect -500 3680 -440 3700
rect -380 3740 -320 3760
rect -380 3700 -370 3740
rect -330 3700 -320 3740
rect -380 3680 -320 3700
rect -260 3740 -200 3760
rect -260 3700 -250 3740
rect -210 3700 -200 3740
rect -260 3680 -200 3700
rect -140 3740 -80 3760
rect -140 3700 -130 3740
rect -90 3700 -80 3740
rect -140 3680 -80 3700
rect -20 3740 40 3760
rect -20 3700 -10 3740
rect 30 3700 40 3740
rect -20 3680 40 3700
rect 100 3740 160 3760
rect 100 3700 110 3740
rect 150 3700 160 3740
rect 100 3680 160 3700
rect 220 3740 280 3760
rect 220 3700 230 3740
rect 270 3700 280 3740
rect 220 3680 280 3700
rect 340 3740 400 3760
rect 340 3700 350 3740
rect 390 3700 400 3740
rect 340 3680 400 3700
rect 460 3740 520 3760
rect 460 3700 470 3740
rect 510 3700 520 3740
rect 460 3680 520 3700
rect 580 3740 640 3760
rect 580 3700 590 3740
rect 630 3700 640 3740
rect 580 3680 640 3700
rect 810 3740 890 3760
rect 810 3680 820 3740
rect 880 3680 890 3740
rect -559 3632 -501 3640
rect -559 3580 -557 3632
rect -505 3580 -501 3632
rect -559 3570 -501 3580
rect -470 3540 -440 3680
rect -260 3540 -230 3680
rect -199 3632 -141 3640
rect -199 3580 -197 3632
rect -145 3580 -141 3632
rect -199 3570 -141 3580
rect -79 3632 -21 3640
rect -79 3580 -77 3632
rect -25 3580 -21 3632
rect -79 3570 -21 3580
rect 10 3540 40 3680
rect 220 3540 250 3680
rect 281 3632 339 3640
rect 281 3580 283 3632
rect 335 3580 339 3632
rect 281 3570 339 3580
rect 401 3632 459 3640
rect 401 3580 403 3632
rect 455 3580 459 3632
rect 401 3570 459 3580
rect 490 3540 520 3680
rect 810 3660 890 3680
rect 810 3600 820 3660
rect 880 3600 890 3660
rect 810 3590 890 3600
rect -1250 3530 -1170 3540
rect -1250 3470 -1240 3530
rect -1180 3470 -1170 3530
rect -1250 3210 -1170 3470
rect -500 3530 -420 3540
rect -500 3470 -490 3530
rect -430 3470 -420 3530
rect -500 3460 -420 3470
rect -280 3530 -200 3540
rect -280 3470 -270 3530
rect -210 3470 -200 3530
rect -280 3460 -200 3470
rect -20 3530 60 3540
rect -20 3470 -10 3530
rect 50 3470 60 3530
rect -20 3460 60 3470
rect 200 3530 280 3540
rect 200 3470 210 3530
rect 270 3470 280 3530
rect 200 3460 280 3470
rect 460 3530 540 3540
rect 460 3470 470 3530
rect 530 3470 540 3530
rect 460 3460 540 3470
rect -1250 3170 -1230 3210
rect -1190 3170 -1170 3210
rect -1070 3420 -990 3430
rect -1070 3360 -1060 3420
rect -1000 3360 -990 3420
rect -1070 3340 -990 3360
rect -1070 3280 -1060 3340
rect -1000 3280 -990 3340
rect -1070 3260 -990 3280
rect -1070 3200 -1060 3260
rect -1000 3200 -990 3260
rect -1070 3190 -990 3200
rect -830 3420 -750 3430
rect -830 3360 -820 3420
rect -760 3360 -750 3420
rect -830 3340 -750 3360
rect -830 3280 -820 3340
rect -760 3280 -750 3340
rect -830 3260 -750 3280
rect -830 3200 -820 3260
rect -760 3200 -750 3260
rect -830 3190 -750 3200
rect -590 3420 -510 3430
rect -590 3360 -580 3420
rect -520 3360 -510 3420
rect -590 3340 -510 3360
rect -590 3280 -580 3340
rect -520 3280 -510 3340
rect -590 3260 -510 3280
rect -590 3200 -580 3260
rect -520 3200 -510 3260
rect -590 3190 -510 3200
rect -350 3420 -270 3430
rect -350 3360 -340 3420
rect -280 3360 -270 3420
rect -350 3340 -270 3360
rect -350 3280 -340 3340
rect -280 3280 -270 3340
rect -350 3260 -270 3280
rect -350 3200 -340 3260
rect -280 3200 -270 3260
rect -350 3190 -270 3200
rect 290 3420 370 3430
rect 290 3360 300 3420
rect 360 3360 370 3420
rect 290 3340 370 3360
rect 290 3280 300 3340
rect 360 3280 370 3340
rect 290 3260 370 3280
rect 290 3200 300 3260
rect 360 3200 370 3260
rect 290 3190 370 3200
rect 530 3420 610 3430
rect 530 3360 540 3420
rect 600 3360 610 3420
rect 530 3340 610 3360
rect 530 3280 540 3340
rect 600 3280 610 3340
rect 530 3260 610 3280
rect 530 3200 540 3260
rect 600 3200 610 3260
rect 530 3190 610 3200
rect 770 3420 850 3430
rect 770 3360 780 3420
rect 840 3360 850 3420
rect 770 3340 850 3360
rect 770 3280 780 3340
rect 840 3280 850 3340
rect 770 3260 850 3280
rect 770 3200 780 3260
rect 840 3200 850 3260
rect 770 3190 850 3200
rect 1080 3220 1140 4740
rect -1250 3150 -1170 3170
rect 1080 3180 1090 3220
rect 1130 3180 1140 3220
rect 1080 3160 1140 3180
rect 1170 3820 1410 3830
rect 1170 3760 1180 3820
rect 1240 3760 1260 3820
rect 1320 3760 1340 3820
rect 1400 3760 1410 3820
rect 1170 3740 1410 3760
rect 1170 3680 1180 3740
rect 1240 3680 1260 3740
rect 1320 3680 1340 3740
rect 1400 3680 1410 3740
rect 1170 3660 1410 3680
rect 1170 3600 1180 3660
rect 1240 3600 1260 3660
rect 1320 3600 1340 3660
rect 1400 3600 1410 3660
rect -90 2620 -10 2630
rect -90 2560 -80 2620
rect -20 2560 -10 2620
rect -90 2540 -10 2560
rect -90 2480 -80 2540
rect -20 2480 -10 2540
rect -90 2460 -10 2480
rect -90 2400 -80 2460
rect -20 2400 -10 2460
rect -90 2390 -10 2400
rect 1170 2620 1410 3600
rect 1440 3220 1500 4740
rect 1580 4680 1640 4760
rect 1690 4810 1770 4820
rect 1690 4750 1700 4810
rect 1760 4750 1770 4810
rect 1690 4740 1770 4750
rect 1580 4640 1590 4680
rect 1630 4640 1640 4680
rect 1580 4580 1640 4640
rect 1580 4540 1590 4580
rect 1630 4540 1640 4580
rect 1580 4520 1640 4540
rect 1700 4680 1760 4740
rect 1700 4640 1710 4680
rect 1750 4640 1760 4680
rect 1700 4580 1760 4640
rect 1700 4540 1710 4580
rect 1750 4540 1760 4580
rect 1700 4520 1760 4540
rect 1820 4680 1880 4850
rect 1820 4640 1830 4680
rect 1870 4640 1880 4680
rect 1820 4580 1880 4640
rect 1820 4540 1830 4580
rect 1870 4540 1880 4580
rect 1820 4520 1880 4540
rect 1940 4680 2000 4700
rect 1940 4640 1950 4680
rect 1990 4640 2000 4680
rect 1940 4580 2000 4640
rect 1940 4540 1950 4580
rect 1990 4540 2000 4580
rect 1760 4460 1820 4480
rect 1760 4420 1770 4460
rect 1810 4420 1820 4460
rect 1760 4360 1820 4420
rect 1940 4360 2000 4540
rect 2060 4680 2120 4850
rect 2060 4640 2070 4680
rect 2110 4640 2120 4680
rect 2060 4580 2120 4640
rect 2060 4540 2070 4580
rect 2110 4540 2120 4580
rect 2060 4520 2120 4540
rect 2180 4680 2240 4700
rect 2180 4640 2190 4680
rect 2230 4640 2240 4680
rect 2180 4580 2240 4640
rect 2180 4540 2190 4580
rect 2230 4540 2240 4580
rect 2180 4480 2240 4540
rect 2300 4680 2360 4850
rect 2410 4810 2490 4820
rect 2410 4750 2420 4810
rect 2480 4750 2490 4810
rect 2410 4740 2490 4750
rect 2300 4640 2310 4680
rect 2350 4640 2360 4680
rect 2300 4580 2360 4640
rect 2300 4540 2310 4580
rect 2350 4540 2360 4580
rect 2300 4520 2360 4540
rect 2420 4680 2480 4740
rect 2420 4640 2430 4680
rect 2470 4640 2480 4680
rect 2420 4580 2480 4640
rect 2420 4540 2430 4580
rect 2470 4540 2480 4580
rect 2420 4520 2480 4540
rect 2540 4680 2600 4850
rect 2540 4640 2550 4680
rect 2590 4640 2600 4680
rect 2540 4580 2600 4640
rect 2540 4540 2550 4580
rect 2590 4540 2600 4580
rect 2540 4520 2600 4540
rect 2660 4680 2720 4700
rect 2660 4640 2670 4680
rect 2710 4640 2720 4680
rect 2660 4580 2720 4640
rect 2660 4540 2670 4580
rect 2710 4540 2720 4580
rect 2170 4470 2250 4480
rect 2170 4410 2180 4470
rect 2240 4410 2250 4470
rect 2170 4400 2250 4410
rect 2420 4460 2480 4480
rect 2420 4420 2430 4460
rect 2470 4420 2480 4460
rect 2420 4360 2480 4420
rect 2660 4360 2720 4540
rect 2780 4680 2840 4850
rect 2780 4640 2790 4680
rect 2830 4640 2840 4680
rect 2780 4580 2840 4640
rect 2780 4540 2790 4580
rect 2830 4540 2840 4580
rect 2780 4520 2840 4540
rect 2900 4680 2960 4700
rect 2900 4640 2910 4680
rect 2950 4640 2960 4680
rect 2900 4580 2960 4640
rect 2900 4540 2910 4580
rect 2950 4540 2960 4580
rect 2900 4480 2960 4540
rect 3020 4680 3080 4850
rect 3130 4810 3210 4820
rect 3130 4750 3140 4810
rect 3200 4750 3210 4810
rect 3130 4740 3210 4750
rect 3020 4640 3030 4680
rect 3070 4640 3080 4680
rect 3020 4580 3080 4640
rect 3020 4540 3030 4580
rect 3070 4540 3080 4580
rect 3020 4520 3080 4540
rect 3140 4680 3200 4740
rect 3140 4640 3150 4680
rect 3190 4640 3200 4680
rect 3140 4580 3200 4640
rect 3140 4540 3150 4580
rect 3190 4540 3200 4580
rect 3140 4520 3200 4540
rect 3260 4680 3320 4850
rect 3260 4640 3270 4680
rect 3310 4640 3320 4680
rect 3260 4580 3320 4640
rect 3260 4540 3270 4580
rect 3310 4540 3320 4580
rect 3260 4520 3320 4540
rect 3380 4680 3440 4700
rect 3380 4640 3390 4680
rect 3430 4640 3440 4680
rect 3380 4580 3440 4640
rect 3380 4540 3390 4580
rect 3430 4540 3440 4580
rect 2890 4470 2970 4480
rect 2890 4410 2900 4470
rect 2960 4410 2970 4470
rect 1750 4350 1830 4360
rect 1750 4290 1760 4350
rect 1820 4290 1830 4350
rect 1750 4270 1830 4290
rect 1750 4210 1760 4270
rect 1820 4210 1830 4270
rect 1750 4190 1830 4210
rect 1750 4130 1760 4190
rect 1820 4130 1830 4190
rect 1750 4120 1830 4130
rect 1930 4350 2010 4360
rect 1930 4290 1940 4350
rect 2000 4290 2010 4350
rect 1930 4270 2010 4290
rect 1930 4210 1940 4270
rect 2000 4210 2010 4270
rect 1930 4190 2010 4210
rect 1930 4130 1940 4190
rect 2000 4130 2010 4190
rect 1930 4120 2010 4130
rect 2170 4350 2250 4360
rect 2170 4290 2180 4350
rect 2240 4290 2250 4350
rect 2170 4270 2250 4290
rect 2170 4210 2180 4270
rect 2240 4210 2250 4270
rect 2170 4190 2250 4210
rect 2170 4130 2180 4190
rect 2240 4130 2250 4190
rect 2170 4120 2250 4130
rect 2410 4350 2490 4360
rect 2410 4290 2420 4350
rect 2480 4290 2490 4350
rect 2410 4270 2490 4290
rect 2410 4210 2420 4270
rect 2480 4210 2490 4270
rect 2410 4190 2490 4210
rect 2410 4130 2420 4190
rect 2480 4130 2490 4190
rect 2410 4120 2490 4130
rect 2650 4350 2730 4360
rect 2650 4290 2660 4350
rect 2720 4290 2730 4350
rect 2650 4270 2730 4290
rect 2650 4210 2660 4270
rect 2720 4210 2730 4270
rect 2650 4190 2730 4210
rect 2650 4130 2660 4190
rect 2720 4130 2730 4190
rect 2650 4120 2730 4130
rect 2170 4080 2250 4090
rect 2170 4020 2180 4080
rect 2240 4020 2250 4080
rect 2170 4010 2250 4020
rect 2650 4080 2730 4090
rect 2650 4020 2660 4080
rect 2720 4020 2730 4080
rect 2650 4010 2730 4020
rect 1930 3970 2010 3980
rect 1930 3910 1940 3970
rect 2000 3910 2010 3970
rect 1930 3900 2010 3910
rect 1690 3820 1770 3830
rect 1690 3760 1700 3820
rect 1760 3760 1770 3820
rect 1950 3760 1990 3900
rect 2020 3860 2078 3870
rect 2020 3808 2022 3860
rect 2074 3808 2078 3860
rect 2020 3800 2078 3808
rect 2190 3760 2230 4010
rect 2410 3970 2490 3980
rect 2410 3910 2420 3970
rect 2480 3910 2490 3970
rect 2410 3900 2490 3910
rect 2344 3860 2402 3870
rect 2344 3808 2346 3860
rect 2398 3808 2402 3860
rect 2344 3800 2402 3808
rect 2430 3760 2470 3900
rect 2498 3860 2556 3870
rect 2498 3808 2500 3860
rect 2552 3808 2556 3860
rect 2498 3800 2556 3808
rect 2670 3760 2710 4010
rect 2890 3970 2970 4410
rect 3140 4460 3200 4480
rect 3140 4420 3150 4460
rect 3190 4420 3200 4460
rect 3140 4360 3200 4420
rect 3380 4360 3440 4540
rect 3500 4680 3560 4850
rect 3500 4640 3510 4680
rect 3550 4640 3560 4680
rect 3500 4580 3560 4640
rect 3500 4540 3510 4580
rect 3550 4540 3560 4580
rect 3500 4520 3560 4540
rect 3620 4680 3680 4700
rect 3620 4640 3630 4680
rect 3670 4640 3680 4680
rect 3620 4580 3680 4640
rect 3620 4540 3630 4580
rect 3670 4540 3680 4580
rect 3620 4480 3680 4540
rect 3740 4680 3800 4850
rect 3850 4810 3930 5760
rect 4160 5520 4240 5530
rect 4160 5460 4170 5520
rect 4230 5460 4240 5520
rect 4160 5450 4240 5460
rect 3970 5080 4050 5090
rect 3970 5020 3980 5080
rect 4040 5020 4050 5080
rect 3970 5000 4050 5020
rect 3970 4940 3980 5000
rect 4040 4940 4050 5000
rect 3970 4920 4050 4940
rect 3970 4860 3980 4920
rect 4040 4860 4050 4920
rect 3970 4850 4050 4860
rect 3850 4750 3860 4810
rect 3920 4750 3930 4810
rect 3850 4740 3930 4750
rect 3980 4800 4040 4850
rect 3980 4760 3990 4800
rect 4030 4760 4040 4800
rect 3740 4640 3750 4680
rect 3790 4640 3800 4680
rect 3740 4580 3800 4640
rect 3740 4540 3750 4580
rect 3790 4540 3800 4580
rect 3740 4520 3800 4540
rect 3860 4680 3920 4740
rect 3860 4640 3870 4680
rect 3910 4640 3920 4680
rect 3860 4580 3920 4640
rect 3860 4540 3870 4580
rect 3910 4540 3920 4580
rect 3860 4520 3920 4540
rect 3980 4680 4040 4760
rect 3980 4640 3990 4680
rect 4030 4640 4040 4680
rect 3980 4580 4040 4640
rect 3980 4540 3990 4580
rect 4030 4540 4040 4580
rect 3980 4520 4040 4540
rect 3610 4470 3690 4480
rect 3610 4410 3620 4470
rect 3680 4410 3690 4470
rect 3610 4400 3690 4410
rect 3800 4450 3860 4470
rect 3800 4410 3810 4450
rect 3850 4410 3860 4450
rect 3800 4360 3860 4410
rect 3130 4350 3210 4360
rect 3130 4290 3140 4350
rect 3200 4290 3210 4350
rect 3130 4270 3210 4290
rect 3130 4210 3140 4270
rect 3200 4210 3210 4270
rect 3130 4190 3210 4210
rect 3130 4130 3140 4190
rect 3200 4130 3210 4190
rect 3130 4080 3210 4130
rect 3370 4350 3450 4360
rect 3370 4290 3380 4350
rect 3440 4290 3450 4350
rect 3370 4270 3450 4290
rect 3370 4210 3380 4270
rect 3440 4210 3450 4270
rect 3370 4190 3450 4210
rect 3370 4130 3380 4190
rect 3440 4130 3450 4190
rect 3370 4120 3450 4130
rect 3790 4350 3870 4360
rect 3790 4290 3800 4350
rect 3860 4290 3870 4350
rect 3790 4270 3870 4290
rect 3790 4210 3800 4270
rect 3860 4210 3870 4270
rect 3790 4190 3870 4210
rect 3790 4130 3800 4190
rect 3860 4130 3870 4190
rect 3790 4120 3870 4130
rect 3130 4020 3140 4080
rect 3200 4020 3210 4080
rect 3130 4010 3210 4020
rect 2890 3910 2900 3970
rect 2960 3910 2970 3970
rect 2890 3900 2970 3910
rect 2822 3860 2880 3870
rect 2822 3808 2824 3860
rect 2876 3808 2880 3860
rect 2822 3800 2880 3808
rect 2910 3760 2950 3900
rect 2980 3860 3038 3870
rect 2980 3808 2982 3860
rect 3034 3808 3038 3860
rect 2980 3800 3038 3808
rect 1690 3740 1770 3760
rect 1690 3680 1700 3740
rect 1760 3680 1770 3740
rect 1940 3740 2000 3760
rect 1940 3700 1950 3740
rect 1990 3700 2000 3740
rect 1940 3680 2000 3700
rect 2060 3740 2120 3760
rect 2060 3700 2070 3740
rect 2110 3700 2120 3740
rect 2060 3680 2120 3700
rect 2180 3740 2240 3760
rect 2180 3700 2190 3740
rect 2230 3700 2240 3740
rect 2180 3680 2240 3700
rect 2300 3740 2360 3760
rect 2300 3700 2310 3740
rect 2350 3700 2360 3740
rect 2300 3680 2360 3700
rect 2420 3740 2480 3760
rect 2420 3700 2430 3740
rect 2470 3700 2480 3740
rect 2420 3680 2480 3700
rect 2540 3740 2600 3760
rect 2540 3700 2550 3740
rect 2590 3700 2600 3740
rect 2540 3680 2600 3700
rect 2660 3740 2720 3760
rect 2660 3700 2670 3740
rect 2710 3700 2720 3740
rect 2660 3680 2720 3700
rect 2780 3740 2840 3760
rect 2780 3700 2790 3740
rect 2830 3700 2840 3740
rect 2780 3680 2840 3700
rect 2900 3740 2960 3760
rect 2900 3700 2910 3740
rect 2950 3700 2960 3740
rect 2900 3680 2960 3700
rect 3020 3740 3080 3760
rect 3020 3700 3030 3740
rect 3070 3700 3080 3740
rect 3020 3680 3080 3700
rect 3140 3740 3200 4010
rect 3140 3700 3150 3740
rect 3190 3700 3200 3740
rect 3140 3680 3200 3700
rect 1690 3660 1770 3680
rect 1690 3600 1700 3660
rect 1760 3600 1770 3660
rect 1690 3590 1770 3600
rect 2060 3540 2090 3680
rect 2121 3632 2179 3640
rect 2121 3580 2125 3632
rect 2177 3580 2179 3632
rect 2121 3570 2179 3580
rect 2241 3632 2299 3640
rect 2241 3580 2245 3632
rect 2297 3580 2299 3632
rect 2241 3570 2299 3580
rect 2330 3540 2360 3680
rect 2540 3540 2570 3680
rect 2601 3632 2659 3640
rect 2601 3580 2605 3632
rect 2657 3580 2659 3632
rect 2601 3570 2659 3580
rect 2721 3632 2779 3640
rect 2721 3580 2725 3632
rect 2777 3580 2779 3632
rect 2721 3570 2779 3580
rect 2810 3540 2840 3680
rect 3020 3540 3050 3680
rect 4180 3650 4220 5450
rect 4250 5410 4330 5420
rect 4250 5350 4260 5410
rect 4320 5350 4330 5410
rect 4250 5340 4330 5350
rect 4270 3880 4310 5340
rect 6930 5140 7010 9290
rect 7990 9350 8070 9420
rect 8210 9760 8290 9940
rect 8650 10000 8730 10010
rect 8650 9940 8660 10000
rect 8720 9940 8730 10000
rect 8210 9720 8230 9760
rect 8270 9720 8290 9760
rect 8210 9660 8290 9720
rect 8210 9620 8230 9660
rect 8270 9620 8290 9660
rect 8210 9560 8290 9620
rect 8210 9520 8230 9560
rect 8270 9520 8290 9560
rect 8210 9460 8290 9520
rect 8210 9420 8230 9460
rect 8270 9420 8290 9460
rect 8210 9400 8290 9420
rect 8430 9760 8510 9780
rect 8430 9720 8450 9760
rect 8490 9720 8510 9760
rect 8430 9660 8510 9720
rect 8430 9620 8450 9660
rect 8490 9620 8510 9660
rect 8430 9560 8510 9620
rect 8430 9520 8450 9560
rect 8490 9520 8510 9560
rect 8430 9460 8510 9520
rect 8430 9420 8450 9460
rect 8490 9420 8510 9460
rect 7990 9290 8000 9350
rect 8060 9290 8070 9350
rect 7990 9280 8070 9290
rect 8210 9340 8290 9360
rect 8210 9300 8230 9340
rect 8270 9300 8290 9340
rect 7150 9230 7230 9240
rect 7150 9170 7160 9230
rect 7220 9170 7230 9230
rect 7150 7890 7230 9170
rect 8210 9230 8290 9300
rect 8430 9350 8510 9420
rect 8650 9760 8730 9940
rect 8970 10000 9050 10010
rect 8970 9940 8980 10000
rect 9040 9940 9050 10000
rect 8970 9780 9050 9940
rect 9290 10000 9370 10010
rect 9290 9940 9300 10000
rect 9360 9940 9370 10000
rect 8650 9720 8670 9760
rect 8710 9720 8730 9760
rect 8650 9660 8730 9720
rect 8650 9620 8670 9660
rect 8710 9620 8730 9660
rect 8650 9560 8730 9620
rect 8650 9520 8670 9560
rect 8710 9520 8730 9560
rect 8650 9460 8730 9520
rect 8650 9420 8670 9460
rect 8710 9420 8730 9460
rect 8650 9400 8730 9420
rect 8870 9760 9150 9780
rect 8870 9720 8890 9760
rect 8930 9720 8990 9760
rect 9030 9720 9090 9760
rect 9130 9720 9150 9760
rect 8870 9660 9150 9720
rect 8870 9620 8890 9660
rect 8930 9620 8990 9660
rect 9030 9620 9090 9660
rect 9130 9620 9150 9660
rect 8870 9560 9150 9620
rect 8870 9520 8890 9560
rect 8930 9520 8990 9560
rect 9030 9520 9090 9560
rect 9130 9520 9150 9560
rect 8870 9460 9150 9520
rect 8870 9420 8890 9460
rect 8930 9420 8990 9460
rect 9030 9420 9090 9460
rect 9130 9420 9150 9460
rect 8870 9400 9150 9420
rect 9290 9760 9370 9940
rect 9730 10000 9810 10010
rect 9730 9940 9740 10000
rect 9800 9940 9810 10000
rect 9290 9720 9310 9760
rect 9350 9720 9370 9760
rect 9290 9660 9370 9720
rect 9290 9620 9310 9660
rect 9350 9620 9370 9660
rect 9290 9560 9370 9620
rect 9290 9520 9310 9560
rect 9350 9520 9370 9560
rect 9290 9460 9370 9520
rect 9290 9420 9310 9460
rect 9350 9420 9370 9460
rect 9290 9400 9370 9420
rect 9510 9760 9590 9780
rect 9510 9720 9530 9760
rect 9570 9720 9590 9760
rect 9510 9660 9590 9720
rect 9510 9620 9530 9660
rect 9570 9620 9590 9660
rect 9510 9560 9590 9620
rect 9510 9520 9530 9560
rect 9570 9520 9590 9560
rect 9510 9460 9590 9520
rect 9510 9420 9530 9460
rect 9570 9420 9590 9460
rect 8430 9290 8440 9350
rect 8500 9290 8510 9350
rect 8430 9280 8510 9290
rect 8870 9350 8950 9360
rect 8870 9290 8880 9350
rect 8940 9290 8950 9350
rect 9510 9350 9590 9420
rect 9730 9760 9810 9940
rect 10170 10000 10250 10010
rect 10170 9940 10180 10000
rect 10240 9940 10250 10000
rect 9730 9720 9750 9760
rect 9790 9720 9810 9760
rect 9730 9660 9810 9720
rect 9730 9620 9750 9660
rect 9790 9620 9810 9660
rect 9730 9560 9810 9620
rect 9730 9520 9750 9560
rect 9790 9520 9810 9560
rect 9730 9460 9810 9520
rect 9730 9420 9750 9460
rect 9790 9420 9810 9460
rect 9730 9400 9810 9420
rect 9950 9760 10030 9780
rect 9950 9720 9970 9760
rect 10010 9720 10030 9760
rect 9950 9660 10030 9720
rect 9950 9620 9970 9660
rect 10010 9620 10030 9660
rect 9950 9560 10030 9620
rect 9950 9520 9970 9560
rect 10010 9520 10030 9560
rect 9950 9460 10030 9520
rect 9950 9420 9970 9460
rect 10010 9420 10030 9460
rect 8210 9170 8220 9230
rect 8280 9170 8290 9230
rect 8210 9160 8290 9170
rect 7790 9010 7870 9020
rect 7790 8950 7800 9010
rect 7860 8950 7870 9010
rect 7790 8770 7870 8950
rect 7790 8730 7810 8770
rect 7850 8730 7870 8770
rect 7790 8710 7870 8730
rect 7350 8660 7430 8680
rect 7350 8620 7370 8660
rect 7410 8620 7430 8660
rect 7350 8560 7430 8620
rect 7350 8520 7370 8560
rect 7410 8520 7430 8560
rect 7350 8460 7430 8520
rect 7350 8420 7370 8460
rect 7410 8420 7430 8460
rect 7350 8360 7430 8420
rect 7350 8320 7370 8360
rect 7410 8320 7430 8360
rect 7350 8240 7430 8320
rect 7350 8200 7370 8240
rect 7410 8200 7430 8240
rect 7350 8160 7430 8200
rect 7350 8100 7360 8160
rect 7420 8100 7430 8160
rect 7350 8090 7430 8100
rect 7570 8660 7650 8680
rect 7570 8620 7590 8660
rect 7630 8620 7650 8660
rect 7570 8560 7650 8620
rect 7570 8520 7590 8560
rect 7630 8520 7650 8560
rect 7570 8460 7650 8520
rect 7570 8420 7590 8460
rect 7630 8420 7650 8460
rect 7570 8360 7650 8420
rect 7570 8320 7590 8360
rect 7630 8320 7650 8360
rect 7570 8160 7650 8320
rect 7790 8660 7870 8680
rect 7790 8620 7810 8660
rect 7850 8620 7870 8660
rect 7790 8560 7870 8620
rect 7790 8520 7810 8560
rect 7850 8520 7870 8560
rect 7790 8460 7870 8520
rect 7790 8420 7810 8460
rect 7850 8420 7870 8460
rect 7790 8360 7870 8420
rect 7790 8320 7810 8360
rect 7850 8320 7870 8360
rect 7790 8300 7870 8320
rect 8010 8660 8090 8680
rect 8010 8620 8030 8660
rect 8070 8620 8090 8660
rect 8010 8560 8090 8620
rect 8010 8520 8030 8560
rect 8070 8520 8090 8560
rect 8010 8460 8090 8520
rect 8010 8420 8030 8460
rect 8070 8420 8090 8460
rect 8010 8360 8090 8420
rect 8010 8320 8030 8360
rect 8070 8320 8090 8360
rect 7570 8100 7580 8160
rect 7640 8100 7650 8160
rect 7570 8090 7650 8100
rect 8010 8160 8090 8320
rect 8230 8660 8510 8680
rect 8230 8620 8250 8660
rect 8290 8620 8350 8660
rect 8390 8620 8450 8660
rect 8490 8620 8510 8660
rect 8230 8560 8510 8620
rect 8230 8520 8250 8560
rect 8290 8520 8350 8560
rect 8390 8520 8450 8560
rect 8490 8520 8510 8560
rect 8230 8460 8510 8520
rect 8230 8420 8250 8460
rect 8290 8420 8350 8460
rect 8390 8420 8450 8460
rect 8490 8420 8510 8460
rect 8230 8360 8510 8420
rect 8230 8320 8250 8360
rect 8290 8320 8350 8360
rect 8390 8320 8450 8360
rect 8490 8320 8510 8360
rect 8230 8300 8510 8320
rect 8650 8660 8730 8680
rect 8650 8620 8670 8660
rect 8710 8620 8730 8660
rect 8650 8560 8730 8620
rect 8650 8520 8670 8560
rect 8710 8520 8730 8560
rect 8650 8460 8730 8520
rect 8650 8420 8670 8460
rect 8710 8420 8730 8460
rect 8650 8360 8730 8420
rect 8650 8320 8670 8360
rect 8710 8320 8730 8360
rect 8010 8100 8020 8160
rect 8080 8100 8090 8160
rect 8010 8090 8090 8100
rect 8330 8160 8410 8300
rect 8330 8100 8340 8160
rect 8400 8100 8410 8160
rect 8330 8090 8410 8100
rect 8650 8160 8730 8320
rect 8870 8660 8950 9290
rect 9380 9320 9460 9330
rect 9380 9260 9390 9320
rect 9450 9260 9460 9320
rect 9510 9290 9520 9350
rect 9580 9290 9590 9350
rect 9510 9280 9590 9290
rect 9950 9350 10030 9420
rect 10170 9760 10250 9940
rect 10170 9720 10190 9760
rect 10230 9720 10250 9760
rect 10170 9660 10250 9720
rect 10170 9620 10190 9660
rect 10230 9620 10250 9660
rect 10170 9560 10250 9620
rect 10170 9520 10190 9560
rect 10230 9520 10250 9560
rect 10170 9460 10250 9520
rect 10170 9420 10190 9460
rect 10230 9420 10250 9460
rect 10170 9400 10250 9420
rect 10390 10000 10470 10010
rect 10390 9940 10400 10000
rect 10460 9940 10470 10000
rect 10390 9880 10470 9940
rect 10390 9840 10410 9880
rect 10450 9840 10470 9880
rect 10390 9760 10470 9840
rect 10390 9720 10410 9760
rect 10450 9720 10470 9760
rect 10390 9660 10470 9720
rect 10390 9620 10410 9660
rect 10450 9620 10470 9660
rect 10390 9560 10470 9620
rect 10390 9520 10410 9560
rect 10450 9520 10470 9560
rect 10390 9460 10470 9520
rect 10390 9420 10410 9460
rect 10450 9420 10470 9460
rect 10390 9400 10470 9420
rect 9950 9290 9960 9350
rect 10020 9290 10030 9350
rect 10750 9340 10860 9360
rect 9380 9120 9460 9260
rect 9380 9060 9390 9120
rect 9450 9060 9460 9120
rect 9380 9050 9460 9060
rect 9950 9070 10030 9290
rect 10080 9320 10160 9330
rect 10080 9260 10090 9320
rect 10150 9260 10160 9320
rect 10080 9250 10160 9260
rect 10750 9270 10770 9340
rect 10840 9270 10860 9340
rect 10750 9250 10860 9270
rect 9950 9010 9960 9070
rect 10020 9010 10030 9070
rect 9820 8820 9900 8830
rect 9820 8760 9830 8820
rect 9890 8760 9900 8820
rect 9820 8750 9900 8760
rect 8870 8620 8890 8660
rect 8930 8620 8950 8660
rect 8870 8560 8950 8620
rect 8870 8520 8890 8560
rect 8930 8520 8950 8560
rect 8870 8460 8950 8520
rect 8870 8420 8890 8460
rect 8930 8420 8950 8460
rect 8870 8360 8950 8420
rect 8870 8320 8890 8360
rect 8930 8320 8950 8360
rect 8870 8300 8950 8320
rect 9090 8660 9170 8680
rect 9090 8620 9110 8660
rect 9150 8620 9170 8660
rect 9090 8560 9170 8620
rect 9090 8520 9110 8560
rect 9150 8520 9170 8560
rect 9090 8460 9170 8520
rect 9090 8420 9110 8460
rect 9150 8420 9170 8460
rect 9090 8360 9170 8420
rect 9090 8320 9110 8360
rect 9150 8320 9170 8360
rect 8650 8100 8660 8160
rect 8720 8100 8730 8160
rect 8650 8090 8730 8100
rect 9090 8160 9170 8320
rect 9310 8660 9590 8680
rect 9310 8620 9330 8660
rect 9370 8620 9430 8660
rect 9470 8620 9530 8660
rect 9570 8620 9590 8660
rect 9310 8560 9590 8620
rect 9310 8520 9330 8560
rect 9370 8520 9430 8560
rect 9470 8520 9530 8560
rect 9570 8520 9590 8560
rect 9310 8460 9590 8520
rect 9310 8420 9330 8460
rect 9370 8420 9430 8460
rect 9470 8420 9530 8460
rect 9570 8420 9590 8460
rect 9310 8360 9590 8420
rect 9310 8320 9330 8360
rect 9370 8320 9430 8360
rect 9470 8320 9530 8360
rect 9570 8320 9590 8360
rect 9310 8300 9590 8320
rect 9730 8660 9810 8680
rect 9730 8620 9750 8660
rect 9790 8620 9810 8660
rect 9730 8560 9810 8620
rect 9730 8520 9750 8560
rect 9790 8520 9810 8560
rect 9730 8460 9810 8520
rect 9730 8420 9750 8460
rect 9790 8420 9810 8460
rect 9730 8360 9810 8420
rect 9730 8320 9750 8360
rect 9790 8320 9810 8360
rect 9090 8100 9100 8160
rect 9160 8100 9170 8160
rect 9090 8090 9170 8100
rect 9410 8160 9490 8300
rect 9410 8100 9420 8160
rect 9480 8100 9490 8160
rect 9410 8090 9490 8100
rect 9730 8160 9810 8320
rect 9950 8660 10030 9010
rect 14010 9070 14090 14050
rect 14010 9010 14020 9070
rect 14080 9010 14090 9070
rect 10080 8820 10160 8830
rect 10080 8760 10090 8820
rect 10150 8760 10160 8820
rect 10080 8750 10160 8760
rect 10750 8810 10860 8830
rect 10750 8740 10770 8810
rect 10840 8740 10860 8810
rect 10750 8720 10860 8740
rect 9950 8620 9970 8660
rect 10010 8620 10030 8660
rect 9950 8560 10030 8620
rect 9950 8520 9970 8560
rect 10010 8520 10030 8560
rect 9950 8460 10030 8520
rect 9950 8420 9970 8460
rect 10010 8420 10030 8460
rect 9950 8360 10030 8420
rect 9950 8320 9970 8360
rect 10010 8320 10030 8360
rect 9950 8300 10030 8320
rect 10170 8660 10250 8680
rect 10170 8620 10190 8660
rect 10230 8620 10250 8660
rect 10170 8560 10250 8620
rect 10170 8520 10190 8560
rect 10230 8520 10250 8560
rect 10170 8460 10250 8520
rect 10170 8420 10190 8460
rect 10230 8420 10250 8460
rect 10170 8360 10250 8420
rect 10170 8320 10190 8360
rect 10230 8320 10250 8360
rect 9730 8100 9740 8160
rect 9800 8100 9810 8160
rect 9730 8090 9810 8100
rect 10170 8160 10250 8320
rect 10170 8100 10180 8160
rect 10240 8100 10250 8160
rect 10170 8090 10250 8100
rect 10390 8660 10470 8680
rect 10390 8620 10410 8660
rect 10450 8620 10470 8660
rect 10390 8560 10470 8620
rect 10390 8520 10410 8560
rect 10450 8520 10470 8560
rect 10390 8460 10470 8520
rect 10390 8420 10410 8460
rect 10450 8420 10470 8460
rect 10390 8360 10470 8420
rect 10390 8320 10410 8360
rect 10450 8320 10470 8360
rect 10390 8240 10470 8320
rect 10390 8200 10410 8240
rect 10450 8200 10470 8240
rect 10390 8160 10470 8200
rect 10390 8100 10400 8160
rect 10460 8100 10470 8160
rect 10390 8090 10470 8100
rect 11100 8020 11210 8040
rect 11100 7950 11120 8020
rect 11190 7950 11210 8020
rect 11100 7930 11210 7950
rect 7150 7830 7160 7890
rect 7220 7830 7230 7890
rect 7150 7820 7230 7830
rect 13900 7890 13980 7900
rect 13900 7830 13910 7890
rect 13970 7830 13980 7890
rect 6930 5080 6940 5140
rect 7000 5080 7010 5140
rect 6930 5070 7010 5080
rect 7040 7780 7120 7790
rect 7040 7720 7050 7780
rect 7110 7720 7120 7780
rect 7040 7700 7120 7720
rect 7040 7640 7050 7700
rect 7110 7640 7120 7700
rect 7040 7620 7120 7640
rect 7040 7560 7050 7620
rect 7110 7560 7120 7620
rect 7040 4980 7120 7560
rect 11220 7260 11320 7280
rect 11220 7200 11240 7260
rect 11300 7200 11320 7260
rect 11220 7180 11320 7200
rect 11020 6740 11100 6750
rect 11020 6680 11030 6740
rect 11090 6680 11100 6740
rect 11020 6670 11100 6680
rect 11230 6688 11310 7180
rect 7040 4920 7050 4980
rect 7110 4920 7120 4980
rect 7040 4910 7120 4920
rect 7150 6340 7230 6360
rect 7150 6300 7170 6340
rect 7210 6300 7230 6340
rect 5580 4810 5660 4820
rect 5580 4750 5590 4810
rect 5650 4750 5660 4810
rect 4360 4350 4600 4360
rect 4360 4290 4370 4350
rect 4430 4290 4450 4350
rect 4510 4290 4530 4350
rect 4590 4290 4600 4350
rect 4360 4270 4600 4290
rect 4360 4210 4370 4270
rect 4430 4210 4450 4270
rect 4510 4210 4530 4270
rect 4590 4210 4600 4270
rect 4360 4190 4600 4210
rect 4360 4130 4370 4190
rect 4430 4130 4450 4190
rect 4510 4130 4530 4190
rect 4590 4130 4600 4190
rect 4250 3870 4330 3880
rect 4250 3810 4260 3870
rect 4320 3810 4330 3870
rect 4250 3800 4330 3810
rect 4160 3640 4240 3650
rect 3081 3632 3139 3640
rect 3081 3580 3085 3632
rect 3137 3580 3139 3632
rect 3081 3570 3139 3580
rect 4160 3580 4170 3640
rect 4230 3580 4240 3640
rect 4160 3570 4240 3580
rect 2040 3530 2120 3540
rect 2040 3470 2050 3530
rect 2110 3470 2120 3530
rect 2040 3460 2120 3470
rect 2300 3530 2380 3540
rect 2300 3470 2310 3530
rect 2370 3470 2380 3530
rect 2300 3460 2380 3470
rect 2520 3530 2600 3540
rect 2520 3470 2530 3530
rect 2590 3470 2600 3530
rect 2520 3460 2600 3470
rect 2780 3530 2860 3540
rect 2780 3470 2790 3530
rect 2850 3470 2860 3530
rect 2780 3460 2860 3470
rect 3000 3530 3080 3540
rect 3000 3470 3010 3530
rect 3070 3470 3080 3530
rect 3000 3460 3080 3470
rect 3750 3530 3830 3540
rect 3750 3470 3760 3530
rect 3820 3470 3830 3530
rect 3750 3460 3830 3470
rect 1440 3180 1450 3220
rect 1490 3180 1500 3220
rect 1730 3420 1810 3430
rect 1730 3360 1740 3420
rect 1800 3360 1810 3420
rect 1730 3340 1810 3360
rect 1730 3280 1740 3340
rect 1800 3280 1810 3340
rect 1730 3260 1810 3280
rect 1730 3200 1740 3260
rect 1800 3200 1810 3260
rect 1730 3190 1810 3200
rect 1970 3420 2050 3430
rect 1970 3360 1980 3420
rect 2040 3360 2050 3420
rect 1970 3340 2050 3360
rect 1970 3280 1980 3340
rect 2040 3280 2050 3340
rect 1970 3260 2050 3280
rect 1970 3200 1980 3260
rect 2040 3200 2050 3260
rect 1970 3190 2050 3200
rect 2210 3420 2290 3430
rect 2210 3360 2220 3420
rect 2280 3360 2290 3420
rect 2210 3340 2290 3360
rect 2210 3280 2220 3340
rect 2280 3280 2290 3340
rect 2210 3260 2290 3280
rect 2210 3200 2220 3260
rect 2280 3200 2290 3260
rect 2210 3190 2290 3200
rect 2850 3420 2930 3430
rect 2850 3360 2860 3420
rect 2920 3360 2930 3420
rect 2850 3340 2930 3360
rect 2850 3280 2860 3340
rect 2920 3280 2930 3340
rect 2850 3260 2930 3280
rect 2850 3200 2860 3260
rect 2920 3200 2930 3260
rect 2850 3190 2930 3200
rect 3090 3420 3170 3430
rect 3090 3360 3100 3420
rect 3160 3360 3170 3420
rect 3090 3340 3170 3360
rect 3090 3280 3100 3340
rect 3160 3280 3170 3340
rect 3090 3260 3170 3280
rect 3090 3200 3100 3260
rect 3160 3200 3170 3260
rect 3090 3190 3170 3200
rect 3330 3420 3410 3430
rect 3330 3360 3340 3420
rect 3400 3360 3410 3420
rect 3330 3340 3410 3360
rect 3330 3280 3340 3340
rect 3400 3280 3410 3340
rect 3330 3260 3410 3280
rect 3330 3200 3340 3260
rect 3400 3200 3410 3260
rect 3330 3190 3410 3200
rect 3570 3420 3650 3430
rect 3570 3360 3580 3420
rect 3640 3360 3650 3420
rect 3570 3340 3650 3360
rect 3570 3280 3580 3340
rect 3640 3280 3650 3340
rect 3570 3260 3650 3280
rect 3570 3200 3580 3260
rect 3640 3200 3650 3260
rect 3570 3190 3650 3200
rect 1440 3160 1500 3180
rect 3760 3130 3820 3460
rect 3760 3090 3770 3130
rect 3810 3090 3820 3130
rect 3760 3030 3820 3090
rect 3760 2990 3770 3030
rect 3810 2990 3820 3030
rect 3760 2930 3820 2990
rect 3760 2890 3770 2930
rect 3810 2890 3820 2930
rect 3760 2830 3820 2890
rect 3760 2790 3770 2830
rect 3810 2790 3820 2830
rect 3760 2730 3820 2790
rect 3760 2690 3770 2730
rect 3810 2690 3820 2730
rect 3760 2670 3820 2690
rect 1170 2560 1180 2620
rect 1240 2560 1260 2620
rect 1320 2560 1340 2620
rect 1400 2560 1410 2620
rect 1170 2540 1410 2560
rect 1170 2480 1180 2540
rect 1240 2480 1260 2540
rect 1320 2480 1340 2540
rect 1400 2480 1410 2540
rect 1170 2460 1410 2480
rect 1170 2400 1180 2460
rect 1240 2400 1260 2460
rect 1320 2400 1340 2460
rect 1400 2400 1410 2460
rect 1170 2390 1410 2400
rect 2590 2620 2670 2630
rect 2590 2560 2600 2620
rect 2660 2560 2670 2620
rect 2590 2540 2670 2560
rect 2590 2480 2600 2540
rect 2660 2480 2670 2540
rect 2590 2460 2670 2480
rect 2590 2400 2600 2460
rect 2660 2400 2670 2460
rect 2590 2390 2670 2400
rect -830 2350 -750 2360
rect -830 2290 -820 2350
rect -760 2290 -750 2350
rect -830 2280 -750 2290
rect -670 2350 -590 2360
rect -670 2290 -660 2350
rect -600 2290 -590 2350
rect -670 2280 -590 2290
rect -510 2350 -430 2360
rect -510 2290 -500 2350
rect -440 2290 -430 2350
rect -510 2280 -430 2290
rect -350 2350 -270 2360
rect -350 2290 -340 2350
rect -280 2290 -270 2350
rect -350 2280 -270 2290
rect -190 2350 -110 2360
rect -190 2290 -180 2350
rect -120 2290 -110 2350
rect -190 2280 -110 2290
rect -30 2350 50 2360
rect -30 2290 -20 2350
rect 40 2290 50 2350
rect -30 2280 50 2290
rect 130 2350 210 2360
rect 130 2290 140 2350
rect 200 2290 210 2350
rect 130 2280 210 2290
rect 290 2350 370 2360
rect 290 2290 300 2350
rect 360 2290 370 2350
rect 290 2280 370 2290
rect 450 2350 530 2360
rect 450 2290 460 2350
rect 520 2290 530 2350
rect 450 2280 530 2290
rect 610 2350 690 2360
rect 610 2290 620 2350
rect 680 2290 690 2350
rect 610 2280 690 2290
rect 770 2350 850 2360
rect 770 2290 780 2350
rect 840 2290 850 2350
rect 770 2280 850 2290
rect 930 2350 1010 2360
rect 930 2290 940 2350
rect 1000 2290 1010 2350
rect 930 2280 1010 2290
rect 1090 2350 1170 2360
rect 1090 2290 1100 2350
rect 1160 2290 1170 2350
rect 1090 2280 1170 2290
rect 1250 2350 1330 2360
rect 1250 2290 1260 2350
rect 1320 2290 1330 2350
rect 1250 2280 1330 2290
rect 1410 2350 1490 2360
rect 1410 2290 1420 2350
rect 1480 2290 1490 2350
rect 1410 2280 1490 2290
rect 1570 2350 1650 2360
rect 1570 2290 1580 2350
rect 1640 2290 1650 2350
rect 1570 2280 1650 2290
rect 1730 2350 1810 2360
rect 1730 2290 1740 2350
rect 1800 2290 1810 2350
rect 1730 2280 1810 2290
rect 1890 2350 1970 2360
rect 1890 2290 1900 2350
rect 1960 2290 1970 2350
rect 1890 2280 1970 2290
rect 2050 2350 2130 2360
rect 2050 2290 2060 2350
rect 2120 2290 2130 2350
rect 2050 2280 2130 2290
rect 2210 2350 2290 2360
rect 2210 2290 2220 2350
rect 2280 2290 2290 2350
rect 2210 2280 2290 2290
rect 2370 2350 2450 2360
rect 2370 2290 2380 2350
rect 2440 2290 2450 2350
rect 2370 2280 2450 2290
rect 2530 2350 2610 2360
rect 2530 2290 2540 2350
rect 2600 2290 2610 2350
rect 2530 2280 2610 2290
rect 2690 2350 2770 2360
rect 2690 2290 2700 2350
rect 2760 2290 2770 2350
rect 2690 2280 2770 2290
rect 2850 2350 2930 2360
rect 2850 2290 2860 2350
rect 2920 2290 2930 2350
rect 2850 2280 2930 2290
rect 3010 2350 3090 2360
rect 3010 2290 3020 2350
rect 3080 2290 3090 2350
rect 3010 2280 3090 2290
rect 3170 2350 3250 2360
rect 3170 2290 3180 2350
rect 3240 2290 3250 2350
rect 3170 2280 3250 2290
rect 3480 2220 3560 2230
rect -910 2180 -830 2190
rect -910 2120 -900 2180
rect -840 2120 -830 2180
rect -910 2110 -830 2120
rect 3480 2160 3490 2220
rect 3550 2160 3560 2220
rect 3480 2140 3560 2160
rect 3480 2080 3490 2140
rect 3550 2080 3560 2140
rect 3480 2070 3560 2080
rect -1370 1950 -1360 2010
rect -1300 1950 -1290 2010
rect -1370 1940 -1290 1950
rect -960 2010 -880 2020
rect -960 1950 -950 2010
rect -890 1950 -880 2010
rect -2310 1840 -2300 1900
rect -2240 1840 -2230 1900
rect -2310 1830 -2230 1840
rect -1640 1670 -1560 1680
rect -1640 1610 -1630 1670
rect -1570 1610 -1560 1670
rect -1640 20 -1560 1610
rect -1640 -370 -1620 20
rect -1580 -370 -1560 20
rect -1640 -390 -1560 -370
rect -2420 -896 -2400 -506
rect -2360 -896 -2340 -506
rect -3526 -904 -3476 -900
rect -3526 -1301 -3520 -904
rect -3482 -1301 -3476 -904
rect -2420 -916 -2340 -896
rect -3526 -1313 -3476 -1301
rect -3540 -1710 -3460 -1700
rect -3540 -2110 -3530 -1710
rect -3470 -2110 -3460 -1710
rect -3540 -2130 -3460 -2110
rect -3120 -1720 -3040 -1700
rect -3120 -1780 -3110 -1720
rect -3050 -1780 -3040 -1720
rect -3120 -1800 -3040 -1780
rect -3120 -1860 -3110 -1800
rect -3050 -1860 -3040 -1800
rect -3120 -1890 -3040 -1860
rect -3120 -1950 -3110 -1890
rect -3050 -1950 -3040 -1890
rect -3120 -1980 -3040 -1950
rect -3120 -2040 -3110 -1980
rect -3050 -2040 -3040 -1980
rect -3120 -2060 -3040 -2040
rect -3120 -2120 -3110 -2060
rect -3050 -2120 -3040 -2060
rect -3540 -2240 -3460 -2220
rect -3540 -2280 -3520 -2240
rect -3480 -2280 -3460 -2240
rect -3540 -2530 -3460 -2280
rect -3540 -2590 -3530 -2530
rect -3470 -2590 -3460 -2530
rect -3540 -2610 -3460 -2590
rect -3540 -2670 -3530 -2610
rect -3470 -2670 -3460 -2610
rect -3540 -2690 -3460 -2670
rect -3540 -2750 -3530 -2690
rect -3470 -2750 -3460 -2690
rect -3540 -2760 -3460 -2750
rect -3120 -2800 -3040 -2120
rect -2750 -1730 -2670 -1700
rect -2750 -2120 -2740 -1730
rect -2700 -2120 -2670 -1730
rect -2750 -2240 -2670 -2120
rect -2750 -2280 -2730 -2240
rect -2690 -2280 -2670 -2240
rect -2750 -2530 -2670 -2280
rect -2750 -2590 -2740 -2530
rect -2680 -2590 -2670 -2530
rect -2750 -2610 -2670 -2590
rect -2750 -2670 -2740 -2610
rect -2680 -2670 -2670 -2610
rect -2750 -2690 -2670 -2670
rect -2750 -2750 -2740 -2690
rect -2680 -2750 -2670 -2690
rect -2750 -2760 -2670 -2750
rect -1310 -1720 -1230 -1700
rect -1310 -2110 -1290 -1720
rect -1250 -2110 -1230 -1720
rect -1310 -2240 -1230 -2110
rect -1310 -2280 -1290 -2240
rect -1250 -2280 -1230 -2240
rect -1310 -2530 -1230 -2280
rect -1310 -2590 -1300 -2530
rect -1240 -2590 -1230 -2530
rect -1310 -2610 -1230 -2590
rect -1310 -2670 -1300 -2610
rect -1240 -2670 -1230 -2610
rect -1310 -2690 -1230 -2670
rect -1310 -2750 -1300 -2690
rect -1240 -2750 -1230 -2690
rect -1310 -2760 -1230 -2750
rect -3120 -2860 -3110 -2800
rect -3050 -2860 -3040 -2800
rect -3120 -2870 -3040 -2860
rect -960 -2870 -880 1950
rect 4180 1800 4220 3570
rect 4160 1790 4240 1800
rect -850 1780 -770 1790
rect -850 1720 -840 1780
rect -780 1720 -770 1780
rect 552 1720 562 1790
rect 632 1720 642 1790
rect 1950 1720 1960 1790
rect 2030 1720 2040 1790
rect 4160 1730 4170 1790
rect 4230 1730 4240 1790
rect 4160 1720 4240 1730
rect -850 -420 -770 1720
rect 1960 1670 2040 1720
rect 1960 1610 1970 1670
rect 2030 1610 2040 1670
rect 1960 1600 2040 1610
rect 4270 1600 4310 3800
rect 3350 1590 3430 1600
rect 3350 1530 3360 1590
rect 3420 1530 3430 1590
rect -850 -480 -840 -420
rect -780 -480 -770 -420
rect -850 -490 -770 -480
rect -420 1170 3000 1260
rect -420 1136 -330 1170
rect -296 1136 -230 1170
rect -196 1136 -130 1170
rect -96 1136 -30 1170
rect 4 1136 70 1170
rect 104 1136 170 1170
rect 204 1136 1030 1170
rect 1064 1136 1130 1170
rect 1164 1136 1230 1170
rect 1264 1136 1330 1170
rect 1364 1136 1430 1170
rect 1464 1136 1530 1170
rect 1564 1136 2390 1170
rect 2424 1136 2490 1170
rect 2524 1136 2590 1170
rect 2624 1136 2690 1170
rect 2724 1136 2790 1170
rect 2824 1136 2890 1170
rect 2924 1136 3000 1170
rect -420 1070 3000 1136
rect -420 1036 -330 1070
rect -296 1036 -230 1070
rect -196 1036 -130 1070
rect -96 1036 -30 1070
rect 4 1036 70 1070
rect 104 1036 170 1070
rect 204 1036 1030 1070
rect 1064 1036 1130 1070
rect 1164 1036 1230 1070
rect 1264 1036 1330 1070
rect 1364 1036 1430 1070
rect 1464 1036 1530 1070
rect 1564 1036 2390 1070
rect 2424 1036 2490 1070
rect 2524 1036 2590 1070
rect 2624 1036 2690 1070
rect 2724 1036 2790 1070
rect 2824 1036 2890 1070
rect 2924 1036 3000 1070
rect -420 970 3000 1036
rect -420 936 -330 970
rect -296 936 -230 970
rect -196 936 -130 970
rect -96 936 -30 970
rect 4 936 70 970
rect 104 936 170 970
rect 204 936 1030 970
rect 1064 936 1130 970
rect 1164 936 1230 970
rect 1264 936 1330 970
rect 1364 936 1430 970
rect 1464 936 1530 970
rect 1564 936 2390 970
rect 2424 936 2490 970
rect 2524 936 2590 970
rect 2624 936 2690 970
rect 2724 936 2790 970
rect 2824 936 2890 970
rect 2924 936 3000 970
rect -420 870 3000 936
rect -420 836 -330 870
rect -296 836 -230 870
rect -196 836 -130 870
rect -96 836 -30 870
rect 4 836 70 870
rect 104 836 170 870
rect 204 836 1030 870
rect 1064 836 1130 870
rect 1164 836 1230 870
rect 1264 836 1330 870
rect 1364 836 1430 870
rect 1464 836 1530 870
rect 1564 836 2390 870
rect 2424 836 2490 870
rect 2524 836 2590 870
rect 2624 836 2690 870
rect 2724 836 2790 870
rect 2824 836 2890 870
rect 2924 836 3000 870
rect -420 770 3000 836
rect -420 736 -330 770
rect -296 736 -230 770
rect -196 736 -130 770
rect -96 736 -30 770
rect 4 736 70 770
rect 104 736 170 770
rect 204 736 1030 770
rect 1064 736 1130 770
rect 1164 736 1230 770
rect 1264 736 1330 770
rect 1364 736 1430 770
rect 1464 736 1530 770
rect 1564 736 2390 770
rect 2424 736 2490 770
rect 2524 736 2590 770
rect 2624 736 2690 770
rect 2724 736 2790 770
rect 2824 736 2890 770
rect 2924 736 3000 770
rect -420 670 3000 736
rect -420 636 -330 670
rect -296 636 -230 670
rect -196 636 -130 670
rect -96 636 -30 670
rect 4 636 70 670
rect 104 636 170 670
rect 204 636 1030 670
rect 1064 636 1130 670
rect 1164 636 1230 670
rect 1264 636 1330 670
rect 1364 636 1430 670
rect 1464 636 1530 670
rect 1564 636 2390 670
rect 2424 636 2490 670
rect 2524 636 2590 670
rect 2624 636 2690 670
rect 2724 636 2790 670
rect 2824 636 2890 670
rect 2924 636 3000 670
rect -420 560 3000 636
rect -420 -190 280 560
rect -420 -224 -330 -190
rect -296 -224 -230 -190
rect -196 -224 -130 -190
rect -96 -224 -30 -190
rect 4 -224 70 -190
rect 104 -224 170 -190
rect 204 -224 280 -190
rect -420 -290 280 -224
rect -420 -324 -330 -290
rect -296 -324 -230 -290
rect -196 -324 -130 -290
rect -96 -324 -30 -290
rect 4 -324 70 -290
rect 104 -324 170 -290
rect 204 -324 280 -290
rect -420 -390 280 -324
rect -420 -420 -330 -390
rect -420 -480 -410 -420
rect -350 -424 -330 -420
rect -296 -424 -230 -390
rect -196 -424 -130 -390
rect -96 -424 -30 -390
rect 4 -424 70 -390
rect 104 -424 170 -390
rect 204 -424 280 -390
rect -350 -480 280 -424
rect -420 -490 280 -480
rect -420 -524 -330 -490
rect -296 -524 -230 -490
rect -196 -524 -130 -490
rect -96 -524 -30 -490
rect 4 -524 70 -490
rect 104 -524 170 -490
rect 204 -524 280 -490
rect -420 -590 280 -524
rect -420 -624 -330 -590
rect -296 -624 -230 -590
rect -196 -624 -130 -590
rect -96 -624 -30 -590
rect 4 -624 70 -590
rect 104 -624 170 -590
rect 204 -624 280 -590
rect -420 -690 280 -624
rect -420 -724 -330 -690
rect -296 -724 -230 -690
rect -196 -724 -130 -690
rect -96 -724 -30 -690
rect 4 -724 70 -690
rect 104 -724 170 -690
rect 204 -724 280 -690
rect -420 -1460 280 -724
rect 940 -190 1640 -100
rect 940 -224 1030 -190
rect 1064 -224 1130 -190
rect 1164 -224 1230 -190
rect 1264 -224 1330 -190
rect 1364 -224 1430 -190
rect 1464 -224 1530 -190
rect 1564 -224 1640 -190
rect 940 -290 1640 -224
rect 940 -324 1030 -290
rect 1064 -324 1130 -290
rect 1164 -324 1230 -290
rect 1264 -324 1330 -290
rect 1364 -324 1430 -290
rect 1464 -324 1530 -290
rect 1564 -324 1640 -290
rect 940 -390 1640 -324
rect 940 -424 1030 -390
rect 1064 -424 1130 -390
rect 1164 -424 1230 -390
rect 1264 -420 1330 -390
rect 1320 -424 1330 -420
rect 1364 -424 1430 -390
rect 1464 -424 1530 -390
rect 1564 -424 1640 -390
rect 940 -480 1260 -424
rect 1320 -480 1640 -424
rect 940 -490 1640 -480
rect 940 -524 1030 -490
rect 1064 -524 1130 -490
rect 1164 -524 1230 -490
rect 1264 -524 1330 -490
rect 1364 -524 1430 -490
rect 1464 -524 1530 -490
rect 1564 -524 1640 -490
rect 940 -590 1640 -524
rect 940 -624 1030 -590
rect 1064 -624 1130 -590
rect 1164 -624 1230 -590
rect 1264 -624 1330 -590
rect 1364 -624 1430 -590
rect 1464 -624 1530 -590
rect 1564 -624 1640 -590
rect 940 -690 1640 -624
rect 940 -724 1030 -690
rect 1064 -724 1130 -690
rect 1164 -724 1230 -690
rect 1264 -724 1330 -690
rect 1364 -724 1430 -690
rect 1464 -724 1530 -690
rect 1564 -724 1640 -690
rect 940 -800 1640 -724
rect 2300 -190 3000 560
rect 2300 -224 2390 -190
rect 2424 -224 2490 -190
rect 2524 -224 2590 -190
rect 2624 -224 2690 -190
rect 2724 -224 2790 -190
rect 2824 -224 2890 -190
rect 2924 -224 3000 -190
rect 2300 -290 3000 -224
rect 2300 -324 2390 -290
rect 2424 -324 2490 -290
rect 2524 -324 2590 -290
rect 2624 -324 2690 -290
rect 2724 -324 2790 -290
rect 2824 -324 2890 -290
rect 2924 -324 3000 -290
rect 2300 -390 3000 -324
rect 2300 -424 2390 -390
rect 2424 -424 2490 -390
rect 2524 -424 2590 -390
rect 2624 -424 2690 -390
rect 2724 -424 2790 -390
rect 2824 -424 2890 -390
rect 2924 -424 3000 -390
rect 2300 -490 3000 -424
rect 3350 -420 3430 1530
rect 4010 1590 4090 1600
rect 4010 1530 4020 1590
rect 4080 1530 4090 1590
rect 4010 20 4090 1530
rect 4250 1590 4330 1600
rect 4250 1530 4260 1590
rect 4320 1530 4330 1590
rect 4250 1520 4330 1530
rect 4360 1040 4600 4130
rect 4360 980 4370 1040
rect 4430 980 4450 1040
rect 4510 980 4530 1040
rect 4590 980 4600 1040
rect 4360 960 4600 980
rect 4790 1900 4870 1910
rect 4790 1840 4800 1900
rect 4860 1840 4870 1900
rect 4010 -370 4030 20
rect 4070 -370 4090 20
rect 4010 -390 4090 -370
rect 3350 -480 3360 -420
rect 3420 -480 3430 -420
rect 3350 -490 3430 -480
rect 2300 -524 2390 -490
rect 2424 -524 2490 -490
rect 2524 -524 2590 -490
rect 2624 -524 2690 -490
rect 2724 -524 2790 -490
rect 2824 -524 2890 -490
rect 2924 -524 3000 -490
rect 2300 -590 3000 -524
rect 2300 -624 2390 -590
rect 2424 -624 2490 -590
rect 2524 -624 2590 -590
rect 2624 -624 2690 -590
rect 2724 -624 2790 -590
rect 2824 -624 2890 -590
rect 2924 -624 3000 -590
rect 2300 -690 3000 -624
rect 2300 -724 2390 -690
rect 2424 -724 2490 -690
rect 2524 -724 2590 -690
rect 2624 -724 2690 -690
rect 2724 -724 2790 -690
rect 2824 -724 2890 -690
rect 2924 -724 3000 -690
rect 2300 -1460 3000 -724
rect -420 -1550 3000 -1460
rect 4790 -1111 4870 1840
rect 4790 -1508 4813 -1111
rect 4851 -1508 4870 -1111
rect 5580 -360 5660 4750
rect 7150 3600 7230 6300
rect 11230 6291 11250 6688
rect 11288 6291 11310 6688
rect 11230 6280 11310 6291
rect 11244 6279 11294 6280
rect 11230 6117 11310 6130
rect 7610 6030 7690 6050
rect 7610 5980 7630 6030
rect 7670 5980 7690 6030
rect 7610 5890 7690 5980
rect 7610 5840 7630 5890
rect 7670 5840 7690 5890
rect 7410 5760 7490 5780
rect 7410 5720 7430 5760
rect 7470 5720 7490 5760
rect 7410 5620 7490 5720
rect 7410 5560 7420 5620
rect 7480 5560 7490 5620
rect 7410 5550 7490 5560
rect 7610 5620 7690 5840
rect 8010 6030 8090 6050
rect 8010 5980 8030 6030
rect 8070 5980 8090 6030
rect 8010 5890 8090 5980
rect 8010 5840 8030 5890
rect 8070 5840 8090 5890
rect 7610 5560 7620 5620
rect 7680 5560 7690 5620
rect 7610 5550 7690 5560
rect 7850 5620 7930 5630
rect 7850 5560 7860 5620
rect 7920 5560 7930 5620
rect 7850 5550 7930 5560
rect 8010 5620 8090 5840
rect 8010 5560 8020 5620
rect 8080 5560 8090 5620
rect 8010 5550 8090 5560
rect 8410 6030 8490 6050
rect 8410 5980 8430 6030
rect 8470 5980 8490 6030
rect 8410 5890 8490 5980
rect 8410 5840 8430 5890
rect 8470 5840 8490 5890
rect 8410 5620 8490 5840
rect 8410 5560 8420 5620
rect 8480 5560 8490 5620
rect 8410 5550 8490 5560
rect 8810 6030 8890 6050
rect 8810 5980 8830 6030
rect 8870 5980 8890 6030
rect 8810 5890 8890 5980
rect 8810 5840 8830 5890
rect 8870 5840 8890 5890
rect 8810 5620 8890 5840
rect 9210 6030 9290 6050
rect 9210 5980 9230 6030
rect 9270 5980 9290 6030
rect 9210 5890 9290 5980
rect 9210 5840 9230 5890
rect 9270 5840 9290 5890
rect 8810 5560 8820 5620
rect 8880 5560 8890 5620
rect 8810 5550 8890 5560
rect 8990 5730 9070 5740
rect 8990 5670 9000 5730
rect 9060 5670 9070 5730
rect 8990 5510 9070 5670
rect 9210 5620 9290 5840
rect 9210 5560 9220 5620
rect 9280 5560 9290 5620
rect 9210 5550 9290 5560
rect 9410 5760 9490 5780
rect 9410 5720 9430 5760
rect 9470 5720 9490 5760
rect 9410 5620 9490 5720
rect 11230 5720 11250 6117
rect 11288 5720 11310 6117
rect 9410 5560 9420 5620
rect 9480 5560 9490 5620
rect 9410 5550 9490 5560
rect 10130 5620 10210 5630
rect 10130 5560 10140 5620
rect 10200 5560 10210 5620
rect 10130 5550 10210 5560
rect 8990 5450 9000 5510
rect 9060 5450 9070 5510
rect 8990 5440 9070 5450
rect 7460 5340 7540 5360
rect 7460 5300 7480 5340
rect 7520 5300 7540 5340
rect 7460 5280 7540 5300
rect 7590 5340 7670 5360
rect 7590 5300 7610 5340
rect 7650 5300 7670 5340
rect 7590 5280 7670 5300
rect 7720 5340 7800 5360
rect 7720 5300 7740 5340
rect 7780 5300 7800 5340
rect 7720 5220 7800 5300
rect 7850 5340 7930 5360
rect 7850 5300 7870 5340
rect 7910 5300 7930 5340
rect 7850 5280 7930 5300
rect 7980 5340 8060 5360
rect 7980 5300 8000 5340
rect 8040 5300 8060 5340
rect 7980 5240 8060 5300
rect 8110 5340 8190 5360
rect 8110 5300 8130 5340
rect 8170 5300 8190 5340
rect 8110 5280 8190 5300
rect 8240 5340 8320 5360
rect 8240 5300 8260 5340
rect 8300 5300 8320 5340
rect 8240 5280 8320 5300
rect 8600 5340 8680 5360
rect 8600 5300 8620 5340
rect 8660 5300 8680 5340
rect 8600 5280 8680 5300
rect 8730 5340 8810 5360
rect 8730 5300 8750 5340
rect 8790 5300 8810 5340
rect 8730 5280 8810 5300
rect 8860 5340 8940 5360
rect 8860 5300 8880 5340
rect 8920 5300 8940 5340
rect 8860 5280 8940 5300
rect 8990 5340 9070 5360
rect 8990 5300 9010 5340
rect 9050 5300 9070 5340
rect 8990 5280 9070 5300
rect 9120 5340 9200 5360
rect 9120 5300 9140 5340
rect 9180 5300 9200 5340
rect 9120 5280 9200 5300
rect 9250 5340 9330 5360
rect 9250 5300 9270 5340
rect 9310 5300 9330 5340
rect 9250 5280 9330 5300
rect 9380 5340 9460 5360
rect 9380 5300 9400 5340
rect 9440 5300 9460 5340
rect 9380 5280 9460 5300
rect 7720 5180 7740 5220
rect 7780 5180 7800 5220
rect 7720 5160 7800 5180
rect 7630 4890 7710 4900
rect 7630 4830 7640 4890
rect 7700 4830 7710 4890
rect 7630 4820 7710 4830
rect 7740 4780 7780 5160
rect 8000 5060 8040 5240
rect 8770 5230 8850 5240
rect 8770 5170 8780 5230
rect 8840 5170 8850 5230
rect 8070 5160 8150 5170
rect 8070 5100 8080 5160
rect 8140 5100 8150 5160
rect 8070 5090 8150 5100
rect 8770 5160 8850 5170
rect 7980 5000 7990 5060
rect 8050 5000 8060 5060
rect 8000 4780 8040 5000
rect 8090 4900 8130 5090
rect 8770 4980 8810 5160
rect 8730 4920 8740 4980
rect 8800 4920 8810 4980
rect 8880 4910 8920 5280
rect 9140 4920 9180 5280
rect 9210 5230 9290 5240
rect 9210 5170 9220 5230
rect 9280 5170 9290 5230
rect 9210 5160 9290 5170
rect 10750 5230 10830 5240
rect 10750 5170 10760 5230
rect 10820 5170 10830 5230
rect 10750 5160 10830 5170
rect 11230 5230 11310 5720
rect 11450 5330 11560 5350
rect 11450 5260 11470 5330
rect 11540 5260 11560 5330
rect 11450 5240 11560 5260
rect 11230 5170 11240 5230
rect 11300 5170 11310 5230
rect 11230 5160 11310 5170
rect 9910 5110 9990 5120
rect 9910 5050 9920 5110
rect 9980 5050 9990 5110
rect 9910 5040 9990 5050
rect 11620 5060 11700 5070
rect 11620 5000 11630 5060
rect 11690 5000 11700 5060
rect 11620 4990 11700 5000
rect 13900 5060 13980 7830
rect 13900 5000 13910 5060
rect 13970 5000 13980 5060
rect 13900 4990 13980 5000
rect 14010 7780 14090 9010
rect 14010 7720 14020 7780
rect 14080 7720 14090 7780
rect 14010 7700 14090 7720
rect 14010 7640 14020 7700
rect 14080 7640 14090 7700
rect 14010 7620 14090 7640
rect 14010 7560 14020 7620
rect 14080 7560 14090 7620
rect 9140 4910 9220 4920
rect 8070 4890 8150 4900
rect 8070 4830 8080 4890
rect 8140 4830 8150 4890
rect 8070 4820 8150 4830
rect 8860 4890 8940 4910
rect 8860 4850 8880 4890
rect 8920 4850 8940 4890
rect 7460 4760 7540 4780
rect 7460 4720 7480 4760
rect 7520 4720 7540 4760
rect 7460 4660 7540 4720
rect 7460 4620 7480 4660
rect 7520 4620 7540 4660
rect 7460 4600 7540 4620
rect 7590 4760 7670 4780
rect 7590 4720 7610 4760
rect 7650 4720 7670 4760
rect 7590 4660 7670 4720
rect 7590 4620 7610 4660
rect 7650 4620 7670 4660
rect 7590 4600 7670 4620
rect 7720 4760 7800 4780
rect 7720 4720 7740 4760
rect 7780 4720 7800 4760
rect 7720 4660 7800 4720
rect 7720 4620 7740 4660
rect 7780 4620 7800 4660
rect 7720 4600 7800 4620
rect 7850 4760 7930 4780
rect 7850 4720 7870 4760
rect 7910 4720 7930 4760
rect 7850 4660 7930 4720
rect 7850 4620 7870 4660
rect 7910 4620 7930 4660
rect 7850 4600 7930 4620
rect 7980 4760 8060 4780
rect 7980 4720 8000 4760
rect 8040 4720 8060 4760
rect 7980 4660 8060 4720
rect 7980 4620 8000 4660
rect 8040 4620 8060 4660
rect 7980 4600 8060 4620
rect 8110 4760 8190 4780
rect 8110 4720 8130 4760
rect 8170 4720 8190 4760
rect 8110 4660 8190 4720
rect 8110 4620 8130 4660
rect 8170 4620 8190 4660
rect 8110 4600 8190 4620
rect 8240 4760 8320 4780
rect 8240 4720 8260 4760
rect 8300 4720 8320 4760
rect 8240 4660 8320 4720
rect 8240 4620 8260 4660
rect 8300 4620 8320 4660
rect 8240 4600 8320 4620
rect 8600 4760 8680 4780
rect 8600 4720 8620 4760
rect 8660 4720 8680 4760
rect 8600 4660 8680 4720
rect 8600 4620 8620 4660
rect 8660 4620 8680 4660
rect 8600 4600 8680 4620
rect 8730 4760 8810 4780
rect 8730 4720 8750 4760
rect 8790 4720 8810 4760
rect 8730 4660 8810 4720
rect 8730 4620 8750 4660
rect 8790 4620 8810 4660
rect 8730 4600 8810 4620
rect 8860 4760 8940 4850
rect 9140 4850 9150 4910
rect 9210 4850 9220 4910
rect 9140 4840 9220 4850
rect 9910 4890 9990 4900
rect 9140 4780 9180 4840
rect 9910 4830 9920 4890
rect 9980 4830 9990 4890
rect 9910 4820 9990 4830
rect 10750 4890 10830 4900
rect 10750 4830 10760 4890
rect 10820 4830 10830 4890
rect 10750 4820 10830 4830
rect 11230 4890 11310 4900
rect 11230 4830 11240 4890
rect 11300 4830 11310 4890
rect 8860 4720 8880 4760
rect 8920 4720 8940 4760
rect 8860 4660 8940 4720
rect 8860 4620 8880 4660
rect 8920 4620 8940 4660
rect 8860 4600 8940 4620
rect 8990 4760 9070 4780
rect 8990 4720 9010 4760
rect 9050 4720 9070 4760
rect 8990 4660 9070 4720
rect 8990 4620 9010 4660
rect 9050 4620 9070 4660
rect 8990 4600 9070 4620
rect 9120 4760 9200 4780
rect 9120 4720 9140 4760
rect 9180 4720 9200 4760
rect 9120 4660 9200 4720
rect 9120 4620 9140 4660
rect 9180 4620 9200 4660
rect 9120 4600 9200 4620
rect 9250 4760 9330 4780
rect 9250 4720 9270 4760
rect 9310 4720 9330 4760
rect 9250 4660 9330 4720
rect 9250 4620 9270 4660
rect 9310 4620 9330 4660
rect 9250 4600 9330 4620
rect 9380 4760 9460 4780
rect 9380 4720 9400 4760
rect 9440 4720 9460 4760
rect 9380 4660 9460 4720
rect 9380 4620 9400 4660
rect 9440 4620 9460 4660
rect 9380 4600 9460 4620
rect 7930 4510 8010 4520
rect 7930 4450 7940 4510
rect 8000 4450 8010 4510
rect 7530 4400 7610 4410
rect 7530 4340 7540 4400
rect 7600 4340 7610 4400
rect 7530 4230 7610 4340
rect 7530 4190 7550 4230
rect 7590 4190 7610 4230
rect 7530 4170 7610 4190
rect 7730 4400 7810 4410
rect 7730 4340 7740 4400
rect 7800 4340 7810 4400
rect 7530 4110 7610 4130
rect 7530 4070 7550 4110
rect 7590 4070 7610 4110
rect 7530 4010 7610 4070
rect 7530 3970 7550 4010
rect 7590 3970 7610 4010
rect 7530 3910 7610 3970
rect 7530 3870 7550 3910
rect 7590 3870 7610 3910
rect 7530 3810 7610 3870
rect 7530 3770 7550 3810
rect 7590 3770 7610 3810
rect 7530 3710 7610 3770
rect 7530 3670 7550 3710
rect 7590 3670 7610 3710
rect 7530 3650 7610 3670
rect 7730 4110 7810 4340
rect 7730 4070 7750 4110
rect 7790 4070 7810 4110
rect 7730 4010 7810 4070
rect 7730 3970 7750 4010
rect 7790 3970 7810 4010
rect 7730 3910 7810 3970
rect 7730 3870 7750 3910
rect 7790 3870 7810 3910
rect 7730 3810 7810 3870
rect 7730 3770 7750 3810
rect 7790 3770 7810 3810
rect 7730 3710 7810 3770
rect 7730 3670 7750 3710
rect 7790 3670 7810 3710
rect 7730 3650 7810 3670
rect 7930 4260 8010 4450
rect 7930 4200 7940 4260
rect 8000 4200 8010 4260
rect 7930 4110 8010 4200
rect 7930 4070 7950 4110
rect 7990 4070 8010 4110
rect 7930 4010 8010 4070
rect 7930 3970 7950 4010
rect 7990 3970 8010 4010
rect 7930 3910 8010 3970
rect 7930 3870 7950 3910
rect 7990 3870 8010 3910
rect 7930 3810 8010 3870
rect 7930 3770 7950 3810
rect 7990 3770 8010 3810
rect 7930 3710 8010 3770
rect 7930 3670 7950 3710
rect 7990 3670 8010 3710
rect 7930 3650 8010 3670
rect 8130 4400 8210 4410
rect 8130 4340 8140 4400
rect 8200 4340 8210 4400
rect 8130 4110 8210 4340
rect 8530 4400 8610 4410
rect 8530 4340 8540 4400
rect 8600 4340 8610 4400
rect 8130 4070 8150 4110
rect 8190 4070 8210 4110
rect 8130 4010 8210 4070
rect 8130 3970 8150 4010
rect 8190 3970 8210 4010
rect 8130 3910 8210 3970
rect 8130 3870 8150 3910
rect 8190 3870 8210 3910
rect 8130 3810 8210 3870
rect 8130 3770 8150 3810
rect 8190 3770 8210 3810
rect 8130 3710 8210 3770
rect 8130 3670 8150 3710
rect 8190 3670 8210 3710
rect 8130 3650 8210 3670
rect 8330 4110 8410 4130
rect 8330 4070 8350 4110
rect 8390 4070 8410 4110
rect 8330 4010 8410 4070
rect 8330 3970 8350 4010
rect 8390 3970 8410 4010
rect 8330 3910 8410 3970
rect 8330 3870 8350 3910
rect 8390 3870 8410 3910
rect 8330 3810 8410 3870
rect 8330 3770 8350 3810
rect 8390 3770 8410 3810
rect 8330 3710 8410 3770
rect 8330 3670 8350 3710
rect 8390 3670 8410 3710
rect 7150 3540 7160 3600
rect 7220 3540 7230 3600
rect 7150 3530 7230 3540
rect 8330 3600 8410 3670
rect 8530 4110 8610 4340
rect 8930 4400 9090 4410
rect 8930 4340 8940 4400
rect 9000 4340 9020 4400
rect 9080 4340 9090 4400
rect 8930 4330 9090 4340
rect 9330 4400 9410 4410
rect 9330 4340 9340 4400
rect 9400 4340 9410 4400
rect 8530 4070 8550 4110
rect 8590 4070 8610 4110
rect 8530 4010 8610 4070
rect 8530 3970 8550 4010
rect 8590 3970 8610 4010
rect 8530 3910 8610 3970
rect 8530 3870 8550 3910
rect 8590 3870 8610 3910
rect 8530 3810 8610 3870
rect 8530 3770 8550 3810
rect 8590 3770 8610 3810
rect 8530 3710 8610 3770
rect 8530 3670 8550 3710
rect 8590 3670 8610 3710
rect 8530 3650 8610 3670
rect 8730 4110 8810 4130
rect 8730 4070 8750 4110
rect 8790 4070 8810 4110
rect 8730 4010 8810 4070
rect 8730 3970 8750 4010
rect 8790 3970 8810 4010
rect 8730 3910 8810 3970
rect 8730 3870 8750 3910
rect 8790 3870 8810 3910
rect 8730 3810 8810 3870
rect 8730 3770 8750 3810
rect 8790 3770 8810 3810
rect 8730 3710 8810 3770
rect 8730 3670 8750 3710
rect 8790 3670 8810 3710
rect 8330 3540 8340 3600
rect 8400 3540 8410 3600
rect 8330 3530 8410 3540
rect 8730 3600 8810 3670
rect 8930 4110 9010 4330
rect 8930 4070 8950 4110
rect 8990 4070 9010 4110
rect 8930 4010 9010 4070
rect 8930 3970 8950 4010
rect 8990 3970 9010 4010
rect 8930 3910 9010 3970
rect 8930 3870 8950 3910
rect 8990 3870 9010 3910
rect 8930 3810 9010 3870
rect 8930 3770 8950 3810
rect 8990 3770 9010 3810
rect 8930 3710 9010 3770
rect 8930 3670 8950 3710
rect 8990 3670 9010 3710
rect 8930 3650 9010 3670
rect 9130 4260 9210 4270
rect 9130 4200 9140 4260
rect 9200 4200 9210 4260
rect 9130 4110 9210 4200
rect 9130 4070 9150 4110
rect 9190 4070 9210 4110
rect 9130 4010 9210 4070
rect 9130 3970 9150 4010
rect 9190 3970 9210 4010
rect 9130 3910 9210 3970
rect 9130 3870 9150 3910
rect 9190 3870 9210 3910
rect 9130 3810 9210 3870
rect 9130 3770 9150 3810
rect 9190 3770 9210 3810
rect 9130 3710 9210 3770
rect 9130 3670 9150 3710
rect 9190 3670 9210 3710
rect 9130 3650 9210 3670
rect 9330 4110 9410 4340
rect 9330 4070 9350 4110
rect 9390 4070 9410 4110
rect 9330 4010 9410 4070
rect 9330 3970 9350 4010
rect 9390 3970 9410 4010
rect 9330 3910 9410 3970
rect 9330 3870 9350 3910
rect 9390 3870 9410 3910
rect 9330 3810 9410 3870
rect 9330 3770 9350 3810
rect 9390 3770 9410 3810
rect 9330 3710 9410 3770
rect 9330 3670 9350 3710
rect 9390 3670 9410 3710
rect 9330 3650 9410 3670
rect 9530 4400 9610 4410
rect 9530 4340 9540 4400
rect 9600 4340 9610 4400
rect 9530 4230 9610 4340
rect 10130 4400 10210 4410
rect 10130 4340 10140 4400
rect 10200 4340 10210 4400
rect 10130 4330 10210 4340
rect 9530 4190 9550 4230
rect 9590 4190 9610 4230
rect 9530 4110 9610 4190
rect 9530 4070 9550 4110
rect 9590 4070 9610 4110
rect 9530 4010 9610 4070
rect 9530 3970 9550 4010
rect 9590 3970 9610 4010
rect 9530 3910 9610 3970
rect 9530 3870 9550 3910
rect 9590 3870 9610 3910
rect 9530 3810 9610 3870
rect 11230 4224 11310 4830
rect 11450 4820 11560 4840
rect 11450 4750 11470 4820
rect 11540 4750 11560 4820
rect 11450 4730 11560 4750
rect 11230 3827 11250 4224
rect 11288 3827 11310 4224
rect 11230 3810 11310 3827
rect 9530 3770 9550 3810
rect 9590 3770 9610 3810
rect 9530 3710 9610 3770
rect 9530 3670 9550 3710
rect 9590 3670 9610 3710
rect 9530 3650 9610 3670
rect 8730 3540 8740 3600
rect 8800 3540 8810 3600
rect 8730 3530 8810 3540
rect 11230 3597 11310 3610
rect 11020 3210 11100 3220
rect 11020 3150 11030 3210
rect 11090 3150 11100 3210
rect 11020 3140 11100 3150
rect 11230 3200 11250 3597
rect 11288 3200 11310 3597
rect 6050 2970 6290 2990
rect 6050 2910 6090 2970
rect 6150 2910 6190 2970
rect 6250 2910 6290 2970
rect 6050 2890 6290 2910
rect 11230 2900 11310 3200
rect 5580 -420 5590 -360
rect 5650 -420 5660 -360
rect 5580 -904 5660 -420
rect 5580 -1301 5600 -904
rect 5638 -1301 5660 -904
rect 5580 -1320 5660 -1301
rect 5960 340 6040 350
rect 5960 280 5970 340
rect 6030 280 6040 340
rect 4790 -1520 4870 -1508
rect -420 -1584 -330 -1550
rect -296 -1584 -230 -1550
rect -196 -1584 -130 -1550
rect -96 -1584 -30 -1550
rect 4 -1584 70 -1550
rect 104 -1584 170 -1550
rect 204 -1584 1030 -1550
rect 1064 -1584 1130 -1550
rect 1164 -1584 1230 -1550
rect 1264 -1584 1330 -1550
rect 1364 -1584 1430 -1550
rect 1464 -1584 1530 -1550
rect 1564 -1584 2390 -1550
rect 2424 -1584 2490 -1550
rect 2524 -1584 2590 -1550
rect 2624 -1584 2690 -1550
rect 2724 -1584 2790 -1550
rect 2824 -1584 2890 -1550
rect 2924 -1584 3000 -1550
rect -420 -1650 3000 -1584
rect -420 -1684 -330 -1650
rect -296 -1684 -230 -1650
rect -196 -1684 -130 -1650
rect -96 -1684 -30 -1650
rect 4 -1684 70 -1650
rect 104 -1684 170 -1650
rect 204 -1684 1030 -1650
rect 1064 -1684 1130 -1650
rect 1164 -1684 1230 -1650
rect 1264 -1684 1330 -1650
rect 1364 -1684 1430 -1650
rect 1464 -1684 1530 -1650
rect 1564 -1684 2390 -1650
rect 2424 -1684 2490 -1650
rect 2524 -1684 2590 -1650
rect 2624 -1684 2690 -1650
rect 2724 -1684 2790 -1650
rect 2824 -1684 2890 -1650
rect 2924 -1684 3000 -1650
rect -420 -1750 3000 -1684
rect 4807 -1700 4857 -1698
rect -420 -1784 -330 -1750
rect -296 -1784 -230 -1750
rect -196 -1784 -130 -1750
rect -96 -1784 -30 -1750
rect 4 -1784 70 -1750
rect 104 -1784 170 -1750
rect 204 -1784 1030 -1750
rect 1064 -1784 1130 -1750
rect 1164 -1784 1230 -1750
rect 1264 -1784 1330 -1750
rect 1364 -1784 1430 -1750
rect 1464 -1784 1530 -1750
rect 1564 -1784 2390 -1750
rect 2424 -1784 2490 -1750
rect 2524 -1784 2590 -1750
rect 2624 -1784 2690 -1750
rect 2724 -1784 2790 -1750
rect 2824 -1784 2890 -1750
rect 2924 -1784 3000 -1750
rect -420 -1850 3000 -1784
rect -420 -1884 -330 -1850
rect -296 -1884 -230 -1850
rect -196 -1884 -130 -1850
rect -96 -1884 -30 -1850
rect 4 -1884 70 -1850
rect 104 -1884 170 -1850
rect 204 -1884 1030 -1850
rect 1064 -1884 1130 -1850
rect 1164 -1884 1230 -1850
rect 1264 -1884 1330 -1850
rect 1364 -1884 1430 -1850
rect 1464 -1884 1530 -1850
rect 1564 -1884 2390 -1850
rect 2424 -1884 2490 -1850
rect 2524 -1884 2590 -1850
rect 2624 -1884 2690 -1850
rect 2724 -1884 2790 -1850
rect 2824 -1884 2890 -1850
rect 2924 -1884 3000 -1850
rect -420 -1950 3000 -1884
rect -420 -1984 -330 -1950
rect -296 -1984 -230 -1950
rect -196 -1984 -130 -1950
rect -96 -1984 -30 -1950
rect 4 -1984 70 -1950
rect 104 -1984 170 -1950
rect 204 -1984 1030 -1950
rect 1064 -1984 1130 -1950
rect 1164 -1984 1230 -1950
rect 1264 -1984 1330 -1950
rect 1364 -1984 1430 -1950
rect 1464 -1984 1530 -1950
rect 1564 -1984 2390 -1950
rect 2424 -1984 2490 -1950
rect 2524 -1984 2590 -1950
rect 2624 -1984 2690 -1950
rect 2724 -1984 2790 -1950
rect 2824 -1984 2890 -1950
rect 2924 -1984 3000 -1950
rect -420 -2050 3000 -1984
rect -420 -2084 -330 -2050
rect -296 -2084 -230 -2050
rect -196 -2084 -130 -2050
rect -96 -2084 -30 -2050
rect 4 -2084 70 -2050
rect 104 -2084 170 -2050
rect 204 -2084 1030 -2050
rect 1064 -2084 1130 -2050
rect 1164 -2084 1230 -2050
rect 1264 -2084 1330 -2050
rect 1364 -2084 1430 -2050
rect 1464 -2084 1530 -2050
rect 1564 -2084 2390 -2050
rect 2424 -2084 2490 -2050
rect 2524 -2084 2590 -2050
rect 2624 -2084 2690 -2050
rect 2724 -2084 2790 -2050
rect 2824 -2084 2890 -2050
rect 2924 -2084 3000 -2050
rect -420 -2160 3000 -2084
rect 3680 -1720 3760 -1700
rect 3680 -2110 3700 -1720
rect 3740 -2110 3760 -1720
rect 3680 -2240 3760 -2110
rect 3680 -2280 3700 -2240
rect 3740 -2280 3760 -2240
rect 1250 -2530 1330 -2520
rect 1250 -2590 1260 -2530
rect 1320 -2590 1330 -2530
rect 1250 -2610 1330 -2590
rect 1250 -2670 1260 -2610
rect 1320 -2670 1330 -2610
rect 1250 -2690 1330 -2670
rect 1250 -2750 1260 -2690
rect 1320 -2750 1330 -2690
rect 1250 -2760 1330 -2750
rect 3680 -2530 3760 -2280
rect 3680 -2590 3690 -2530
rect 3750 -2590 3760 -2530
rect 3680 -2610 3760 -2590
rect 3680 -2670 3690 -2610
rect 3750 -2670 3760 -2610
rect 3680 -2690 3760 -2670
rect 3680 -2750 3690 -2690
rect 3750 -2750 3760 -2690
rect 3680 -2760 3760 -2750
rect 4790 -1710 4870 -1700
rect 4790 -2107 4813 -1710
rect 4851 -2107 4870 -1710
rect 4790 -2240 4870 -2107
rect 5580 -1710 5660 -1700
rect 5580 -2110 5590 -1710
rect 5650 -2110 5660 -1710
rect 5580 -2130 5660 -2110
rect 5960 -1720 6040 280
rect 6130 -1060 6210 2890
rect 11220 2880 11320 2900
rect 11220 2820 11240 2880
rect 11300 2820 11320 2880
rect 11220 2800 11320 2820
rect 6130 -1120 6140 -1060
rect 6200 -1120 6210 -1060
rect 6130 -1130 6210 -1120
rect 6660 2010 6740 2020
rect 6660 1950 6670 2010
rect 6730 1950 6740 2010
rect 5960 -1780 5970 -1720
rect 6030 -1780 6040 -1720
rect 6660 -1740 6740 1950
rect 6790 1040 6890 1060
rect 6790 980 6810 1040
rect 6870 980 6890 1040
rect 6790 960 6890 980
rect 6790 -360 6890 -340
rect 6790 -420 6810 -360
rect 6870 -420 6890 -360
rect 6790 -440 6890 -420
rect 5960 -1800 6040 -1780
rect 5960 -1860 5970 -1800
rect 6030 -1860 6040 -1800
rect 6650 -1760 6750 -1740
rect 6650 -1820 6670 -1760
rect 6730 -1820 6750 -1760
rect 6650 -1840 6750 -1820
rect 5960 -1890 6040 -1860
rect 5960 -1950 5970 -1890
rect 6030 -1950 6040 -1890
rect 5960 -1980 6040 -1950
rect 5960 -2040 5970 -1980
rect 6030 -2040 6040 -1980
rect 5960 -2060 6040 -2040
rect 5960 -2120 5970 -2060
rect 6030 -2120 6040 -2060
rect 5960 -2130 6040 -2120
rect 4790 -2280 4810 -2240
rect 4850 -2280 4870 -2240
rect 4790 -2530 4870 -2280
rect 4790 -2590 4800 -2530
rect 4860 -2590 4870 -2530
rect 4790 -2610 4870 -2590
rect 4790 -2670 4800 -2610
rect 4860 -2670 4870 -2610
rect 4790 -2690 4870 -2670
rect 4790 -2750 4800 -2690
rect 4860 -2750 4870 -2690
rect 4790 -2760 4870 -2750
rect 5580 -2240 5660 -2220
rect 5580 -2280 5600 -2240
rect 5640 -2280 5660 -2240
rect 5580 -2530 5660 -2280
rect 5580 -2590 5590 -2530
rect 5650 -2590 5660 -2530
rect 5580 -2610 5660 -2590
rect 5580 -2670 5590 -2610
rect 5650 -2670 5660 -2610
rect 5580 -2690 5660 -2670
rect 5580 -2750 5590 -2690
rect 5650 -2750 5660 -2690
rect 5580 -2760 5660 -2750
rect 6200 -2460 6280 -2450
rect 6200 -2520 6210 -2460
rect 6270 -2520 6280 -2460
rect 6200 -2800 6280 -2520
rect 6200 -2860 6210 -2800
rect 6270 -2860 6280 -2800
rect 6200 -2870 6280 -2860
rect 14010 -3090 14090 7560
rect 3000 -3110 3430 -3100
rect 3000 -3170 3010 -3110
rect 3420 -3170 3430 -3110
rect 3000 -3180 3430 -3170
rect 4910 -3110 5340 -3100
rect 4910 -3170 4920 -3110
rect 5330 -3170 5340 -3110
rect 4910 -3180 5340 -3170
rect 14000 -3110 14100 -3090
rect 14000 -3170 14020 -3110
rect 14080 -3170 14100 -3110
rect 14000 -3190 14100 -3170
rect 4130 -3300 4210 -3290
rect 4130 -3360 4140 -3300
rect 4200 -3360 4210 -3300
rect 4130 -3370 4210 -3360
<< via1 >>
rect 11330 14770 11390 14830
rect 10830 14660 10890 14720
rect 10910 14660 10970 14720
rect 10990 14660 11050 14720
rect 10830 14580 10890 14640
rect 10910 14580 10970 14640
rect 10990 14580 11050 14640
rect 10830 14500 10890 14560
rect 10910 14500 10970 14560
rect 10990 14500 11050 14560
rect 560 13420 620 13430
rect 560 13380 570 13420
rect 570 13380 610 13420
rect 610 13380 620 13420
rect 560 13370 620 13380
rect 780 13420 840 13430
rect 780 13380 790 13420
rect 790 13380 830 13420
rect 830 13380 840 13420
rect 780 13370 840 13380
rect 1250 13420 1310 13430
rect 1250 13380 1260 13420
rect 1260 13380 1300 13420
rect 1300 13380 1310 13420
rect 1250 13370 1310 13380
rect 1590 13420 1650 13430
rect 1590 13380 1600 13420
rect 1600 13380 1640 13420
rect 1640 13380 1650 13420
rect 1590 13370 1650 13380
rect 1810 13420 1870 13430
rect 1810 13380 1820 13420
rect 1820 13380 1860 13420
rect 1860 13380 1870 13420
rect 1810 13370 1870 13380
rect 2250 13420 2310 13430
rect 2250 13380 2260 13420
rect 2260 13380 2300 13420
rect 2300 13380 2310 13420
rect 2250 13370 2310 13380
rect 2930 13420 2990 13430
rect 2930 13380 2940 13420
rect 2940 13380 2980 13420
rect 2980 13380 2990 13420
rect 2930 13370 2990 13380
rect 3150 13420 3210 13430
rect 3150 13380 3160 13420
rect 3160 13380 3200 13420
rect 3200 13380 3210 13420
rect 3150 13370 3210 13380
rect 3620 13420 3680 13430
rect 3620 13380 3630 13420
rect 3630 13380 3670 13420
rect 3670 13380 3680 13420
rect 3620 13370 3680 13380
rect 4080 13420 4140 13430
rect 4080 13380 4090 13420
rect 4090 13380 4130 13420
rect 4130 13380 4140 13420
rect 4080 13370 4140 13380
rect 4430 13420 4490 13430
rect 4430 13380 4440 13420
rect 4440 13380 4480 13420
rect 4480 13380 4490 13420
rect 4430 13370 4490 13380
rect 4680 13420 4740 13430
rect 4680 13380 4690 13420
rect 4690 13380 4730 13420
rect 4730 13380 4740 13420
rect 4680 13370 4740 13380
rect 4900 13420 4960 13430
rect 4900 13380 4910 13420
rect 4910 13380 4950 13420
rect 4950 13380 4960 13420
rect 4900 13370 4960 13380
rect 5230 13420 5290 13430
rect 5230 13380 5240 13420
rect 5240 13380 5280 13420
rect 5280 13380 5290 13420
rect 5230 13370 5290 13380
rect 5890 13420 5950 13430
rect 5890 13380 5900 13420
rect 5900 13380 5940 13420
rect 5940 13380 5950 13420
rect 5890 13370 5950 13380
rect 6110 13420 6170 13430
rect 6110 13380 6120 13420
rect 6120 13380 6160 13420
rect 6160 13380 6170 13420
rect 6110 13370 6170 13380
rect 6680 13420 6740 13430
rect 6680 13380 6690 13420
rect 6690 13380 6730 13420
rect 6730 13380 6740 13420
rect 6680 13370 6740 13380
rect 6940 13420 7000 13430
rect 6940 13380 6950 13420
rect 6950 13380 6990 13420
rect 6990 13380 7000 13420
rect 6940 13370 7000 13380
rect 7190 13420 7250 13430
rect 7190 13380 7200 13420
rect 7200 13380 7240 13420
rect 7240 13380 7250 13420
rect 7190 13370 7250 13380
rect 7410 13420 7470 13430
rect 7410 13380 7420 13420
rect 7420 13380 7460 13420
rect 7460 13380 7470 13420
rect 7410 13370 7470 13380
rect 7960 13420 8020 13430
rect 7960 13380 7970 13420
rect 7970 13380 8010 13420
rect 8010 13380 8020 13420
rect 7960 13370 8020 13380
rect 8240 13420 8300 13430
rect 8240 13380 8250 13420
rect 8250 13380 8290 13420
rect 8290 13380 8300 13420
rect 8240 13370 8300 13380
rect 8490 13420 8550 13430
rect 8490 13380 8500 13420
rect 8500 13380 8540 13420
rect 8540 13380 8550 13420
rect 8490 13370 8550 13380
rect 8710 13420 8770 13430
rect 8710 13380 8720 13420
rect 8720 13380 8760 13420
rect 8760 13380 8770 13420
rect 8710 13370 8770 13380
rect 9260 13420 9320 13430
rect 9260 13380 9270 13420
rect 9270 13380 9310 13420
rect 9310 13380 9320 13420
rect 9260 13370 9320 13380
rect 9540 13420 9600 13430
rect 9540 13380 9550 13420
rect 9550 13380 9590 13420
rect 9590 13380 9600 13420
rect 9540 13370 9600 13380
rect 9790 13420 9850 13430
rect 9790 13380 9800 13420
rect 9800 13380 9840 13420
rect 9840 13380 9850 13420
rect 9790 13370 9850 13380
rect 10010 13420 10070 13430
rect 10010 13380 10020 13420
rect 10020 13380 10060 13420
rect 10060 13380 10070 13420
rect 10010 13370 10070 13380
rect 10560 13420 10620 13430
rect 10560 13380 10570 13420
rect 10570 13380 10610 13420
rect 10610 13380 10620 13420
rect 10560 13370 10620 13380
rect 130 12990 190 13050
rect 340 13040 400 13050
rect 340 13000 350 13040
rect 350 13000 390 13040
rect 390 13000 400 13040
rect 340 12990 400 13000
rect 11850 14770 11910 14830
rect 12370 14770 12430 14830
rect 12860 14770 12920 14830
rect 13190 14660 13250 14720
rect 13270 14660 13330 14720
rect 13350 14660 13410 14720
rect 13190 14580 13250 14640
rect 13270 14580 13330 14640
rect 13350 14580 13410 14640
rect 13190 14500 13250 14560
rect 13270 14500 13330 14560
rect 13350 14500 13410 14560
rect 11280 14102 11332 14112
rect 11280 14068 11288 14102
rect 11288 14068 11322 14102
rect 11322 14068 11332 14102
rect 11280 14060 11332 14068
rect 11800 14102 11852 14112
rect 11800 14068 11808 14102
rect 11808 14068 11842 14102
rect 11842 14068 11852 14102
rect 11800 14060 11852 14068
rect 11330 13740 11390 13750
rect 11330 13700 11340 13740
rect 11340 13700 11380 13740
rect 11380 13700 11390 13740
rect 11330 13690 11390 13700
rect 11540 13690 11600 13750
rect 11294 13622 11346 13632
rect 11294 13588 11302 13622
rect 11302 13588 11336 13622
rect 11336 13588 11346 13622
rect 11294 13580 11346 13588
rect 11430 13570 11490 13630
rect 10830 13080 10890 13140
rect 10910 13080 10970 13140
rect 10990 13080 11050 13140
rect 10766 13042 10818 13052
rect 10766 13008 10774 13042
rect 10774 13008 10808 13042
rect 10808 13008 10818 13042
rect 10766 13000 10818 13008
rect 10830 13000 10890 13060
rect 10910 13000 10970 13060
rect 10990 13000 11050 13060
rect 10830 12920 10890 12980
rect 10910 12920 10970 12980
rect 10990 12920 11050 12980
rect 11260 13080 11320 13140
rect 11260 13000 11320 13060
rect 11260 12920 11320 12980
rect 11350 13080 11410 13140
rect 11350 13000 11410 13060
rect 11350 12920 11410 12980
rect 720 12640 780 12650
rect 720 12600 730 12640
rect 730 12600 770 12640
rect 770 12600 780 12640
rect 720 12590 780 12600
rect 1140 12640 1200 12650
rect 1140 12600 1150 12640
rect 1150 12600 1190 12640
rect 1190 12600 1200 12640
rect 1140 12590 1200 12600
rect 1810 12640 1870 12650
rect 1810 12600 1820 12640
rect 1820 12600 1860 12640
rect 1860 12600 1870 12640
rect 1810 12590 1870 12600
rect 2380 12640 2440 12650
rect 2380 12600 2390 12640
rect 2390 12600 2430 12640
rect 2430 12600 2440 12640
rect 2380 12590 2440 12600
rect 3090 12640 3150 12650
rect 3090 12600 3100 12640
rect 3100 12600 3140 12640
rect 3140 12600 3150 12640
rect 3090 12590 3150 12600
rect 3520 12640 3580 12650
rect 3520 12600 3530 12640
rect 3530 12600 3570 12640
rect 3570 12600 3580 12640
rect 3520 12590 3580 12600
rect 3960 12640 4020 12650
rect 3960 12600 3970 12640
rect 3970 12600 4010 12640
rect 4010 12600 4020 12640
rect 3960 12590 4020 12600
rect 4210 12640 4270 12650
rect 4210 12600 4220 12640
rect 4220 12600 4260 12640
rect 4260 12600 4270 12640
rect 4210 12590 4270 12600
rect 4430 12640 4490 12650
rect 4430 12600 4440 12640
rect 4440 12600 4480 12640
rect 4480 12600 4490 12640
rect 4430 12590 4490 12600
rect 4900 12640 4960 12650
rect 4900 12600 4910 12640
rect 4910 12600 4950 12640
rect 4950 12600 4960 12640
rect 4900 12590 4960 12600
rect 5340 12640 5400 12650
rect 5340 12600 5350 12640
rect 5350 12600 5390 12640
rect 5390 12600 5400 12640
rect 5340 12590 5400 12600
rect 5960 12640 6020 12650
rect 5960 12600 5970 12640
rect 5970 12600 6010 12640
rect 6010 12600 6020 12640
rect 5960 12590 6020 12600
rect 6300 12640 6360 12650
rect 6300 12600 6310 12640
rect 6310 12600 6350 12640
rect 6350 12600 6360 12640
rect 6300 12590 6360 12600
rect 6660 12640 6720 12650
rect 6660 12600 6670 12640
rect 6670 12600 6710 12640
rect 6710 12600 6720 12640
rect 6660 12590 6720 12600
rect 7260 12640 7320 12650
rect 7260 12600 7270 12640
rect 7270 12600 7310 12640
rect 7310 12600 7320 12640
rect 7260 12590 7320 12600
rect 7600 12640 7660 12650
rect 7600 12600 7610 12640
rect 7610 12600 7650 12640
rect 7650 12600 7660 12640
rect 7600 12590 7660 12600
rect 7960 12640 8020 12650
rect 7960 12600 7970 12640
rect 7970 12600 8010 12640
rect 8010 12600 8020 12640
rect 7960 12590 8020 12600
rect 8560 12640 8620 12650
rect 8560 12600 8570 12640
rect 8570 12600 8610 12640
rect 8610 12600 8620 12640
rect 8560 12590 8620 12600
rect 8900 12640 8960 12650
rect 8900 12600 8910 12640
rect 8910 12600 8950 12640
rect 8950 12600 8960 12640
rect 8900 12590 8960 12600
rect 9260 12640 9320 12650
rect 9260 12600 9270 12640
rect 9270 12600 9310 12640
rect 9310 12600 9320 12640
rect 9260 12590 9320 12600
rect 9860 12640 9920 12650
rect 9860 12600 9870 12640
rect 9870 12600 9910 12640
rect 9910 12600 9920 12640
rect 9860 12590 9920 12600
rect 10200 12640 10260 12650
rect 10200 12600 10210 12640
rect 10210 12600 10250 12640
rect 10250 12600 10260 12640
rect 10200 12590 10260 12600
rect 10560 12640 10620 12650
rect 10560 12600 10570 12640
rect 10570 12600 10610 12640
rect 10610 12600 10620 12640
rect 10560 12590 10620 12600
rect 11294 12272 11346 12282
rect 11294 12238 11302 12272
rect 11302 12238 11336 12272
rect 11336 12238 11346 12272
rect 11294 12230 11346 12238
rect 12320 14102 12372 14112
rect 12320 14068 12328 14102
rect 12328 14068 12362 14102
rect 12362 14068 12372 14102
rect 12320 14060 12372 14068
rect 12886 14102 12938 14112
rect 12886 14068 12896 14102
rect 12896 14068 12930 14102
rect 12930 14068 12938 14102
rect 12886 14060 12938 14068
rect 11850 13740 11910 13750
rect 11850 13700 11860 13740
rect 11860 13700 11900 13740
rect 11900 13700 11910 13740
rect 11850 13690 11910 13700
rect 12060 13690 12120 13750
rect 11814 13622 11866 13632
rect 11814 13588 11822 13622
rect 11822 13588 11856 13622
rect 11856 13588 11866 13622
rect 11814 13580 11866 13588
rect 11950 13570 12010 13630
rect 11780 13080 11840 13140
rect 11780 13000 11840 13060
rect 11780 12920 11840 12980
rect 11870 13080 11930 13140
rect 11870 13000 11930 13060
rect 11870 12920 11930 12980
rect 11540 12230 11600 12290
rect 11330 12160 11390 12170
rect 11330 12120 11340 12160
rect 11340 12120 11380 12160
rect 11380 12120 11390 12160
rect 11330 12110 11390 12120
rect 11430 12110 11490 12170
rect 11814 12272 11866 12282
rect 11814 12238 11822 12272
rect 11822 12238 11856 12272
rect 11856 12238 11866 12272
rect 11814 12230 11866 12238
rect 12370 13740 12430 13750
rect 12370 13700 12380 13740
rect 12380 13700 12420 13740
rect 12420 13700 12430 13740
rect 12370 13690 12430 13700
rect 12580 13690 12640 13750
rect 12334 13622 12386 13632
rect 12334 13588 12342 13622
rect 12342 13588 12376 13622
rect 12376 13588 12386 13622
rect 12334 13580 12386 13588
rect 12470 13570 12530 13630
rect 12300 13080 12360 13140
rect 12300 13000 12360 13060
rect 12300 12920 12360 12980
rect 12390 13080 12450 13140
rect 12390 13000 12450 13060
rect 12390 12920 12450 12980
rect 12060 12230 12120 12290
rect 11330 11520 11390 11580
rect 11600 11520 11660 11580
rect 11410 11390 11470 11400
rect 11410 11350 11420 11390
rect 11420 11350 11460 11390
rect 11460 11350 11470 11390
rect 11410 11340 11470 11350
rect 11850 12160 11910 12170
rect 11850 12120 11860 12160
rect 11860 12120 11900 12160
rect 11900 12120 11910 12160
rect 11850 12110 11910 12120
rect 11950 12110 12010 12170
rect 12334 12272 12386 12282
rect 12334 12238 12342 12272
rect 12342 12238 12376 12272
rect 12376 12238 12386 12272
rect 12334 12230 12386 12238
rect 12580 12230 12640 12290
rect 11850 11520 11910 11580
rect 12120 11520 12180 11580
rect 11930 11390 11990 11400
rect 11930 11350 11940 11390
rect 11940 11350 11980 11390
rect 11980 11350 11990 11390
rect 11930 11340 11990 11350
rect 12370 12160 12430 12170
rect 12370 12120 12380 12160
rect 12380 12120 12420 12160
rect 12420 12120 12430 12160
rect 12370 12110 12430 12120
rect 12470 12110 12530 12170
rect 12370 11520 12430 11580
rect 12640 11520 12700 11580
rect 12450 11390 12510 11400
rect 12450 11350 12460 11390
rect 12460 11350 12500 11390
rect 12500 11350 12510 11390
rect 12450 11340 12510 11350
rect 12780 11340 12840 11400
rect 13190 13080 13250 13140
rect 13270 13080 13330 13140
rect 13350 13080 13410 13140
rect 13190 13000 13250 13060
rect 13270 13000 13330 13060
rect 13350 13000 13410 13060
rect 13190 12920 13250 12980
rect 13270 12920 13330 12980
rect 13350 12920 13410 12980
rect 14020 14050 14080 14110
rect 12970 11390 13030 11400
rect 12970 11350 12980 11390
rect 12980 11350 13020 11390
rect 13020 11350 13030 11390
rect 12970 11340 13030 11350
rect 11600 10690 11660 10750
rect 12120 10690 12180 10750
rect 12640 10690 12700 10750
rect 13160 10690 13220 10750
rect 1270 10440 1330 10450
rect 1270 10400 1280 10440
rect 1280 10400 1320 10440
rect 1320 10400 1330 10440
rect 1270 10390 1330 10400
rect 1490 10440 1550 10450
rect 1490 10400 1500 10440
rect 1500 10400 1540 10440
rect 1540 10400 1550 10440
rect 1490 10390 1550 10400
rect 1790 10440 1850 10450
rect 1790 10400 1800 10440
rect 1800 10400 1840 10440
rect 1840 10400 1850 10440
rect 1790 10390 1850 10400
rect 2010 10440 2070 10450
rect 2010 10400 2020 10440
rect 2020 10400 2060 10440
rect 2060 10400 2070 10440
rect 2010 10390 2070 10400
rect 2170 10440 2230 10450
rect 2170 10400 2180 10440
rect 2180 10400 2220 10440
rect 2220 10400 2230 10440
rect 2170 10390 2230 10400
rect 2390 10440 2450 10450
rect 2390 10400 2400 10440
rect 2400 10400 2440 10440
rect 2440 10400 2450 10440
rect 2390 10390 2450 10400
rect 2690 10440 2750 10450
rect 2690 10400 2700 10440
rect 2700 10400 2740 10440
rect 2740 10400 2750 10440
rect 2690 10390 2750 10400
rect 2910 10440 2970 10450
rect 2910 10400 2920 10440
rect 2920 10400 2960 10440
rect 2960 10400 2970 10440
rect 2910 10390 2970 10400
rect 3210 10440 3270 10450
rect 3210 10400 3220 10440
rect 3220 10400 3260 10440
rect 3260 10400 3270 10440
rect 3210 10390 3270 10400
rect 3650 10440 3710 10450
rect 3650 10400 3660 10440
rect 3660 10400 3700 10440
rect 3700 10400 3710 10440
rect 3650 10390 3710 10400
rect 3980 10440 4040 10450
rect 3980 10400 3990 10440
rect 3990 10400 4030 10440
rect 4030 10400 4040 10440
rect 3980 10390 4040 10400
rect 4410 10440 4470 10450
rect 4410 10400 4420 10440
rect 4420 10400 4460 10440
rect 4460 10400 4470 10440
rect 4410 10390 4470 10400
rect 4800 10440 4860 10450
rect 4800 10400 4810 10440
rect 4810 10400 4850 10440
rect 4850 10400 4860 10440
rect 4800 10390 4860 10400
rect 5190 10440 5250 10450
rect 5190 10400 5200 10440
rect 5200 10400 5240 10440
rect 5240 10400 5250 10440
rect 5190 10390 5250 10400
rect 5710 10450 5770 10510
rect 1680 10330 1740 10340
rect 1680 10290 1690 10330
rect 1690 10290 1730 10330
rect 1730 10290 1740 10330
rect 1680 10280 1740 10290
rect 3400 10330 3460 10340
rect 3400 10290 3410 10330
rect 3410 10290 3450 10330
rect 3450 10290 3460 10330
rect 3400 10280 3460 10290
rect 4250 10260 4310 10320
rect 5480 10330 5540 10340
rect 5480 10290 5490 10330
rect 5490 10290 5530 10330
rect 5530 10290 5540 10330
rect 5480 10280 5540 10290
rect 1150 9950 1210 9960
rect 1150 9910 1160 9950
rect 1160 9910 1200 9950
rect 1200 9910 1210 9950
rect 1150 9900 1210 9910
rect 3050 9980 3110 9990
rect 3050 9940 3060 9980
rect 3060 9940 3100 9980
rect 3100 9940 3110 9980
rect 3050 9930 3110 9940
rect 1270 9260 1330 9270
rect 1270 9220 1280 9260
rect 1280 9220 1320 9260
rect 1320 9220 1330 9260
rect 1270 9210 1330 9220
rect 2010 9260 2070 9270
rect 2010 9220 2020 9260
rect 2020 9220 2060 9260
rect 2060 9220 2070 9260
rect 2010 9210 2070 9220
rect 2170 9260 2230 9270
rect 2170 9220 2180 9260
rect 2180 9220 2220 9260
rect 2220 9220 2230 9260
rect 2170 9210 2230 9220
rect 2910 9260 2970 9270
rect 2910 9220 2920 9260
rect 2920 9220 2960 9260
rect 2960 9220 2970 9260
rect 2910 9210 2970 9220
rect 1720 9150 1780 9160
rect 1720 9110 1730 9150
rect 1730 9110 1770 9150
rect 1770 9110 1780 9150
rect 1720 9100 1780 9110
rect 4140 9940 4200 9950
rect 4140 9900 4150 9940
rect 4150 9900 4190 9940
rect 4190 9900 4200 9940
rect 4140 9890 4200 9900
rect 11010 10450 11080 10520
rect 6420 10280 6480 10340
rect 6020 9990 6080 10000
rect 6020 9950 6030 9990
rect 6030 9950 6070 9990
rect 6070 9950 6080 9990
rect 6020 9940 6080 9950
rect 6310 9940 6370 10000
rect 3270 9370 3330 9380
rect 3270 9330 3280 9370
rect 3280 9330 3320 9370
rect 3320 9330 3330 9370
rect 3270 9320 3330 9330
rect 3160 9260 3220 9270
rect 3160 9220 3170 9260
rect 3170 9220 3210 9260
rect 3210 9220 3220 9260
rect 3160 9210 3220 9220
rect 3350 9260 3410 9270
rect 3350 9220 3360 9260
rect 3360 9220 3400 9260
rect 3400 9220 3410 9260
rect 3350 9210 3410 9220
rect 3430 9260 3490 9270
rect 3430 9220 3440 9260
rect 3440 9220 3480 9260
rect 3480 9220 3490 9260
rect 3430 9210 3490 9220
rect 3640 9260 3700 9270
rect 3640 9220 3650 9260
rect 3650 9220 3690 9260
rect 3690 9220 3700 9260
rect 3640 9210 3700 9220
rect 3970 9260 4030 9270
rect 3970 9220 3980 9260
rect 3980 9220 4020 9260
rect 4020 9220 4030 9260
rect 3970 9210 4030 9220
rect 3250 9100 3310 9160
rect 5710 9910 5770 9920
rect 5710 9870 5720 9910
rect 5720 9870 5760 9910
rect 5760 9870 5770 9910
rect 5710 9860 5770 9870
rect 4410 9260 4470 9270
rect 4410 9220 4420 9260
rect 4420 9220 4460 9260
rect 4460 9220 4470 9260
rect 4410 9210 4470 9220
rect 4800 9260 4860 9270
rect 4800 9220 4810 9260
rect 4810 9220 4850 9260
rect 4850 9220 4860 9260
rect 4800 9210 4860 9220
rect 5010 9210 5070 9270
rect 5190 9260 5250 9270
rect 5190 9220 5200 9260
rect 5200 9220 5240 9260
rect 5240 9220 5250 9260
rect 5190 9210 5250 9220
rect 5870 9260 5930 9270
rect 5870 9220 5880 9260
rect 5880 9220 5920 9260
rect 5920 9220 5930 9260
rect 5870 9210 5930 9220
rect 130 8520 190 8580
rect 1150 8570 1210 8580
rect 1150 8530 1160 8570
rect 1160 8530 1200 8570
rect 1200 8530 1210 8570
rect 1150 8520 1210 8530
rect 3070 8580 3130 8590
rect 3070 8540 3080 8580
rect 3080 8540 3120 8580
rect 3120 8540 3130 8580
rect 3070 8530 3130 8540
rect 4100 8580 4160 8590
rect 4100 8540 4110 8580
rect 4110 8540 4150 8580
rect 4150 8540 4160 8580
rect 4100 8530 4160 8540
rect 4250 9090 4310 9150
rect 4670 9100 4730 9160
rect 4840 9150 4900 9160
rect 4840 9110 4850 9150
rect 4850 9110 4890 9150
rect 4890 9110 4900 9150
rect 4840 9100 4900 9110
rect 5480 9150 5540 9160
rect 5480 9110 5490 9150
rect 5490 9110 5530 9150
rect 5530 9110 5540 9150
rect 5480 9100 5540 9110
rect 6200 9100 6260 9160
rect 7560 9940 7620 10000
rect 7780 9940 7840 10000
rect 8220 9940 8280 10000
rect 6420 9170 6480 9230
rect 6940 9290 7000 9350
rect 6310 9060 6370 9120
rect 6200 8950 6260 9010
rect 6670 8950 6730 9010
rect 6750 8950 6810 9010
rect 6830 8950 6890 9010
rect 6200 8840 6260 8900
rect 6020 8530 6080 8540
rect 6020 8490 6030 8530
rect 6030 8490 6070 8530
rect 6070 8490 6080 8530
rect 6020 8480 6080 8490
rect 6200 8480 6260 8540
rect 4920 8190 4980 8200
rect 4920 8150 4930 8190
rect 4930 8150 4970 8190
rect 4970 8150 4980 8190
rect 4920 8140 4980 8150
rect 5550 8190 5610 8200
rect 5550 8150 5560 8190
rect 5560 8150 5600 8190
rect 5600 8150 5610 8190
rect 5550 8140 5610 8150
rect 6120 8140 6180 8200
rect 1270 8080 1330 8090
rect 1270 8040 1280 8080
rect 1280 8040 1320 8080
rect 1320 8040 1330 8080
rect 1270 8030 1330 8040
rect 1490 8080 1550 8090
rect 1490 8040 1500 8080
rect 1500 8040 1540 8080
rect 1540 8040 1550 8080
rect 1490 8030 1550 8040
rect 1790 8080 1850 8090
rect 1790 8040 1800 8080
rect 1800 8040 1840 8080
rect 1840 8040 1850 8080
rect 1790 8030 1850 8040
rect 2020 8080 2080 8090
rect 2020 8040 2030 8080
rect 2030 8040 2070 8080
rect 2070 8040 2080 8080
rect 2020 8030 2080 8040
rect 2170 8080 2230 8090
rect 2170 8040 2180 8080
rect 2180 8040 2220 8080
rect 2220 8040 2230 8080
rect 2170 8030 2230 8040
rect 2390 8080 2450 8090
rect 2390 8040 2400 8080
rect 2400 8040 2440 8080
rect 2440 8040 2450 8080
rect 2390 8030 2450 8040
rect 2690 8080 2750 8090
rect 2690 8040 2700 8080
rect 2700 8040 2740 8080
rect 2740 8040 2750 8080
rect 2690 8030 2750 8040
rect 2910 8080 2970 8090
rect 2910 8040 2920 8080
rect 2920 8040 2960 8080
rect 2960 8040 2970 8080
rect 2910 8030 2970 8040
rect 3310 8080 3370 8090
rect 3310 8040 3320 8080
rect 3320 8040 3360 8080
rect 3360 8040 3370 8080
rect 3310 8030 3370 8040
rect 3640 8080 3700 8090
rect 3640 8040 3650 8080
rect 3650 8040 3690 8080
rect 3690 8040 3700 8080
rect 3640 8030 3700 8040
rect 3970 8080 4030 8090
rect 3970 8040 3980 8080
rect 3980 8040 4020 8080
rect 4020 8040 4030 8080
rect 3970 8030 4030 8040
rect 4410 8080 4470 8090
rect 4410 8040 4420 8080
rect 4420 8040 4460 8080
rect 4460 8040 4470 8080
rect 4410 8030 4470 8040
rect 4670 8030 4730 8090
rect 5190 8080 5250 8090
rect 5190 8040 5200 8080
rect 5200 8040 5240 8080
rect 5240 8040 5250 8080
rect 5190 8030 5250 8040
rect 5870 8080 5930 8090
rect 5870 8040 5880 8080
rect 5880 8040 5920 8080
rect 5920 8040 5930 8080
rect 5870 8030 5930 8040
rect 6120 7960 6180 8020
rect 1660 7190 1720 7250
rect 1660 7110 1720 7170
rect -2300 7020 -2240 7080
rect -3530 6570 -3470 6630
rect -3530 4750 -3470 4810
rect -2520 5240 -2460 5300
rect -2520 2120 -2460 2180
rect -2410 5130 -2350 5190
rect -2410 3810 -2350 3870
rect -240 7020 -180 7080
rect -20 7020 40 7080
rect 200 7020 260 7080
rect 420 7020 480 7080
rect 640 7020 700 7080
rect 860 7020 920 7080
rect 1660 7030 1720 7090
rect 1880 7190 1940 7250
rect 1880 7110 1940 7170
rect 1880 7030 1940 7090
rect 2100 7190 2160 7250
rect 2100 7110 2160 7170
rect 2100 7030 2160 7090
rect 2320 7190 2380 7250
rect 2320 7110 2380 7170
rect 2320 7030 2380 7090
rect 2540 7190 2600 7250
rect 2540 7110 2600 7170
rect 2540 7030 2600 7090
rect 2760 7190 2820 7250
rect 2760 7110 2820 7170
rect 2760 7030 2820 7090
rect 6670 7190 6730 7250
rect 6750 7190 6810 7250
rect 6830 7190 6890 7250
rect 6670 7110 6730 7170
rect 6750 7110 6810 7170
rect 6830 7110 6890 7170
rect 6670 7030 6730 7090
rect 6750 7030 6810 7090
rect 6830 7030 6890 7090
rect -350 6960 -290 6970
rect -350 6920 -340 6960
rect -340 6920 -300 6960
rect -300 6920 -290 6960
rect -350 6910 -290 6920
rect -130 6910 -70 6970
rect 90 6910 150 6970
rect 310 6910 370 6970
rect 530 6910 590 6970
rect 750 6910 810 6970
rect 970 6960 1030 6970
rect 970 6920 980 6960
rect 980 6920 1020 6960
rect 1020 6920 1030 6960
rect 970 6910 1030 6920
rect 1550 6960 1610 6970
rect 1550 6920 1560 6960
rect 1560 6920 1600 6960
rect 1600 6920 1610 6960
rect 1550 6910 1610 6920
rect 1770 6910 1830 6970
rect 1990 6910 2050 6970
rect 2210 6910 2270 6970
rect 2430 6910 2490 6970
rect 2650 6910 2710 6970
rect 2870 6960 2930 6970
rect 2870 6920 2880 6960
rect 2880 6920 2920 6960
rect 2920 6920 2930 6960
rect 2870 6910 2930 6920
rect -182 6622 -130 6632
rect -182 6588 -172 6622
rect -172 6588 -138 6622
rect -138 6588 -130 6622
rect -182 6580 -130 6588
rect -72 6622 -20 6632
rect -72 6588 -62 6622
rect -62 6588 -28 6622
rect -28 6588 -20 6622
rect -72 6580 -20 6588
rect 38 6622 90 6632
rect 38 6588 48 6622
rect 48 6588 82 6622
rect 82 6588 90 6622
rect 38 6580 90 6588
rect 148 6622 200 6632
rect 148 6588 158 6622
rect 158 6588 192 6622
rect 192 6588 200 6622
rect 148 6580 200 6588
rect 258 6622 310 6632
rect 258 6588 268 6622
rect 268 6588 302 6622
rect 302 6588 310 6622
rect 258 6580 310 6588
rect 368 6622 420 6632
rect 368 6588 378 6622
rect 378 6588 412 6622
rect 412 6588 420 6622
rect 368 6580 420 6588
rect 478 6622 530 6632
rect 478 6588 488 6622
rect 488 6588 522 6622
rect 522 6588 530 6622
rect 478 6580 530 6588
rect 588 6622 640 6632
rect 588 6588 598 6622
rect 598 6588 632 6622
rect 632 6588 640 6622
rect 588 6580 640 6588
rect 698 6622 750 6632
rect 698 6588 708 6622
rect 708 6588 742 6622
rect 742 6588 750 6622
rect 698 6580 750 6588
rect 808 6622 860 6632
rect 808 6588 818 6622
rect 818 6588 852 6622
rect 852 6588 860 6622
rect 808 6580 860 6588
rect 1718 6622 1770 6632
rect 1718 6588 1728 6622
rect 1728 6588 1762 6622
rect 1762 6588 1770 6622
rect 1718 6580 1770 6588
rect 1828 6622 1880 6632
rect 1828 6588 1838 6622
rect 1838 6588 1872 6622
rect 1872 6588 1880 6622
rect 1828 6580 1880 6588
rect 1938 6622 1990 6632
rect 1938 6588 1948 6622
rect 1948 6588 1982 6622
rect 1982 6588 1990 6622
rect 1938 6580 1990 6588
rect 2048 6622 2100 6632
rect 2048 6588 2058 6622
rect 2058 6588 2092 6622
rect 2092 6588 2100 6622
rect 2048 6580 2100 6588
rect 2158 6622 2210 6632
rect 2158 6588 2168 6622
rect 2168 6588 2202 6622
rect 2202 6588 2210 6622
rect 2158 6580 2210 6588
rect 2268 6622 2320 6632
rect 2268 6588 2278 6622
rect 2278 6588 2312 6622
rect 2312 6588 2320 6622
rect 2268 6580 2320 6588
rect 2378 6622 2430 6632
rect 2378 6588 2388 6622
rect 2388 6588 2422 6622
rect 2422 6588 2430 6622
rect 2378 6580 2430 6588
rect 2488 6622 2540 6632
rect 2488 6588 2498 6622
rect 2498 6588 2532 6622
rect 2532 6588 2540 6622
rect 2488 6580 2540 6588
rect 2598 6622 2650 6632
rect 2598 6588 2608 6622
rect 2608 6588 2642 6622
rect 2642 6588 2650 6622
rect 2598 6580 2650 6588
rect 2708 6622 2760 6632
rect 2708 6588 2718 6622
rect 2718 6588 2752 6622
rect 2752 6588 2760 6622
rect 2708 6580 2760 6588
rect -360 6470 -300 6530
rect -360 6390 -300 6450
rect -360 6360 -300 6370
rect -360 6320 -350 6360
rect -350 6320 -310 6360
rect -310 6320 -300 6360
rect -360 6310 -300 6320
rect 0 6470 60 6530
rect 0 6390 60 6450
rect 0 6360 60 6370
rect 0 6320 10 6360
rect 10 6320 50 6360
rect 50 6320 60 6360
rect 0 6310 60 6320
rect 360 6470 420 6530
rect 360 6390 420 6450
rect 360 6360 420 6370
rect 360 6320 370 6360
rect 370 6320 410 6360
rect 410 6320 420 6360
rect 360 6310 420 6320
rect 720 6470 780 6530
rect 720 6390 780 6450
rect 720 6360 780 6370
rect 720 6320 730 6360
rect 730 6320 770 6360
rect 770 6320 780 6360
rect 720 6310 780 6320
rect 1080 6470 1140 6530
rect 1080 6390 1140 6450
rect 1080 6360 1140 6370
rect 1080 6320 1090 6360
rect 1090 6320 1130 6360
rect 1130 6320 1140 6360
rect 1080 6310 1140 6320
rect 1440 6470 1500 6530
rect 1440 6390 1500 6450
rect 1440 6360 1500 6370
rect 1440 6320 1450 6360
rect 1450 6320 1490 6360
rect 1490 6320 1500 6360
rect 1440 6310 1500 6320
rect 1800 6470 1860 6530
rect 1800 6390 1860 6450
rect 1800 6360 1860 6370
rect 1800 6320 1810 6360
rect 1810 6320 1850 6360
rect 1850 6320 1860 6360
rect 1800 6310 1860 6320
rect 2160 6470 2220 6530
rect 2160 6390 2220 6450
rect 2160 6360 2220 6370
rect 2160 6320 2170 6360
rect 2170 6320 2210 6360
rect 2210 6320 2220 6360
rect 2160 6310 2220 6320
rect 2520 6470 2580 6530
rect 2520 6390 2580 6450
rect 2520 6360 2580 6370
rect 2520 6320 2530 6360
rect 2530 6320 2570 6360
rect 2570 6320 2580 6360
rect 2520 6310 2580 6320
rect 2880 6470 2940 6530
rect 2880 6390 2940 6450
rect 2880 6360 2940 6370
rect 2880 6320 2890 6360
rect 2890 6320 2930 6360
rect 2930 6320 2940 6360
rect 2880 6310 2940 6320
rect 3510 6470 3570 6530
rect 3510 6390 3570 6450
rect 3510 6310 3570 6370
rect 3950 6470 4010 6530
rect 3950 6390 4010 6450
rect 3950 6310 4010 6370
rect -90 5620 -30 5630
rect -90 5580 -80 5620
rect -80 5580 -40 5620
rect -40 5580 -30 5620
rect -90 5570 -30 5580
rect 90 5620 150 5630
rect 90 5580 100 5620
rect 100 5580 140 5620
rect 140 5580 150 5620
rect 90 5570 150 5580
rect 270 5620 330 5630
rect 270 5580 280 5620
rect 280 5580 320 5620
rect 320 5580 330 5620
rect 270 5570 330 5580
rect 450 5620 510 5630
rect 450 5580 460 5620
rect 460 5580 500 5620
rect 500 5580 510 5620
rect 450 5570 510 5580
rect 630 5620 690 5630
rect 630 5580 640 5620
rect 640 5580 680 5620
rect 680 5580 690 5620
rect 630 5570 690 5580
rect 810 5620 870 5630
rect 810 5580 820 5620
rect 820 5580 860 5620
rect 860 5580 870 5620
rect 810 5570 870 5580
rect 990 5620 1050 5630
rect 990 5580 1000 5620
rect 1000 5580 1040 5620
rect 1040 5580 1050 5620
rect 990 5570 1050 5580
rect 1170 5620 1230 5630
rect 1170 5580 1180 5620
rect 1180 5580 1220 5620
rect 1220 5580 1230 5620
rect 1170 5570 1230 5580
rect 900 5460 960 5520
rect 540 5350 600 5410
rect 180 5240 240 5300
rect 1350 5620 1410 5630
rect 1350 5580 1360 5620
rect 1360 5580 1400 5620
rect 1400 5580 1410 5620
rect 1350 5570 1410 5580
rect 1440 5570 1500 5630
rect 1530 5620 1590 5630
rect 1530 5580 1540 5620
rect 1540 5580 1580 5620
rect 1580 5580 1590 5620
rect 1530 5570 1590 5580
rect -180 5130 -120 5190
rect 1260 5130 1320 5190
rect -1460 5020 -1400 5080
rect -1460 4940 -1400 5000
rect -1460 4860 -1400 4920
rect -1220 5020 -1160 5080
rect -1220 4940 -1160 5000
rect -1220 4860 -1160 4920
rect -980 5020 -920 5080
rect -980 4940 -920 5000
rect -980 4860 -920 4920
rect -740 5020 -680 5080
rect -740 4940 -680 5000
rect -740 4860 -680 4920
rect -500 5020 -440 5080
rect -500 4940 -440 5000
rect -500 4860 -440 4920
rect -260 5020 -200 5080
rect -260 4940 -200 5000
rect -260 4860 -200 4920
rect -20 5020 40 5080
rect -20 4940 40 5000
rect -20 4860 40 4920
rect 220 5020 280 5080
rect 220 4940 280 5000
rect 220 4860 280 4920
rect 460 5020 520 5080
rect 460 4940 520 5000
rect 460 4860 520 4920
rect 700 5020 760 5080
rect 700 4940 760 5000
rect 700 4860 760 4920
rect 940 5020 1000 5080
rect 940 4940 1000 5000
rect 940 4860 1000 4920
rect -1340 4750 -1280 4810
rect -1100 4460 -1040 4470
rect -1100 4420 -1090 4460
rect -1090 4420 -1050 4460
rect -1050 4420 -1040 4460
rect -1100 4410 -1040 4420
rect -620 4750 -560 4810
rect -380 4460 -320 4470
rect -380 4420 -370 4460
rect -370 4420 -330 4460
rect -330 4420 -320 4460
rect -380 4410 -320 4420
rect -2300 3580 -2240 3640
rect -1360 4290 -1300 4350
rect -1280 4290 -1220 4350
rect -860 4290 -800 4350
rect -620 4290 -560 4350
rect -620 4020 -560 4080
rect 100 4750 160 4810
rect 340 4460 400 4470
rect 340 4420 350 4460
rect 350 4420 390 4460
rect 390 4420 400 4460
rect 340 4410 400 4420
rect 820 4750 880 4810
rect 1080 4750 1140 4810
rect 1710 5620 1770 5630
rect 1710 5580 1720 5620
rect 1720 5580 1760 5620
rect 1760 5580 1770 5620
rect 1710 5570 1770 5580
rect 1890 5620 1950 5630
rect 1890 5580 1900 5620
rect 1900 5580 1940 5620
rect 1940 5580 1950 5620
rect 1890 5570 1950 5580
rect 1620 5460 1680 5520
rect 2070 5620 2130 5630
rect 2070 5580 2080 5620
rect 2080 5580 2120 5620
rect 2120 5580 2130 5620
rect 2070 5570 2130 5580
rect 2250 5620 2310 5630
rect 2250 5580 2260 5620
rect 2260 5580 2300 5620
rect 2300 5580 2310 5620
rect 2250 5570 2310 5580
rect 1980 5350 2040 5410
rect 2430 5620 2490 5630
rect 2430 5580 2440 5620
rect 2440 5580 2480 5620
rect 2480 5580 2490 5620
rect 2430 5570 2490 5580
rect 2610 5620 2670 5630
rect 2610 5580 2620 5620
rect 2620 5580 2660 5620
rect 2660 5580 2670 5620
rect 2610 5570 2670 5580
rect 2340 5240 2400 5300
rect 3260 6110 3320 6170
rect 3730 6160 3790 6170
rect 3730 6120 3740 6160
rect 3740 6120 3780 6160
rect 3780 6120 3790 6160
rect 3730 6110 3790 6120
rect 3610 5820 3670 5830
rect 3610 5780 3620 5820
rect 3620 5780 3660 5820
rect 3660 5780 3670 5820
rect 3610 5770 3670 5780
rect 3260 5350 3320 5410
rect 3850 5820 3910 5830
rect 3850 5780 3860 5820
rect 3860 5780 3900 5820
rect 3900 5780 3910 5820
rect 3850 5770 3910 5780
rect 3730 5240 3790 5300
rect 2700 5130 2760 5190
rect 1580 5020 1640 5080
rect 1580 4940 1640 5000
rect 1580 4860 1640 4920
rect 1820 5020 1880 5080
rect 1820 4940 1880 5000
rect 1820 4860 1880 4920
rect 2060 5020 2120 5080
rect 2060 4940 2120 5000
rect 2060 4860 2120 4920
rect 2300 5020 2360 5080
rect 2300 4940 2360 5000
rect 2300 4860 2360 4920
rect 2540 5020 2600 5080
rect 2540 4940 2600 5000
rect 2540 4860 2600 4920
rect 2780 5020 2840 5080
rect 2780 4940 2840 5000
rect 2780 4860 2840 4920
rect 3020 5020 3080 5080
rect 3020 4940 3080 5000
rect 3020 4860 3080 4920
rect 3260 5020 3320 5080
rect 3260 4940 3320 5000
rect 3260 4860 3320 4920
rect 3500 5020 3560 5080
rect 3500 4940 3560 5000
rect 3500 4860 3560 4920
rect 3740 5020 3800 5080
rect 3740 4940 3800 5000
rect 3740 4860 3800 4920
rect 1440 4750 1500 4810
rect -140 4290 -80 4350
rect 100 4290 160 4350
rect 580 4290 640 4350
rect 760 4290 820 4350
rect -140 4020 -80 4080
rect 340 4020 400 4080
rect -380 3910 -320 3970
rect -454 3852 -402 3860
rect -454 3818 -446 3852
rect -446 3818 -412 3852
rect -412 3818 -402 3852
rect -454 3808 -402 3818
rect -296 3852 -244 3860
rect -296 3818 -288 3852
rect -288 3818 -254 3852
rect -254 3818 -244 3852
rect -296 3808 -244 3818
rect 100 3910 160 3970
rect 28 3852 80 3860
rect 28 3818 36 3852
rect 36 3818 70 3852
rect 70 3818 80 3852
rect 28 3808 80 3818
rect 182 3852 234 3860
rect 182 3818 190 3852
rect 190 3818 224 3852
rect 224 3818 234 3852
rect 182 3808 234 3818
rect 580 3910 640 3970
rect 506 3852 558 3860
rect 506 3818 514 3852
rect 514 3818 548 3852
rect 548 3818 558 3852
rect 506 3808 558 3818
rect 820 3810 880 3820
rect 820 3770 830 3810
rect 830 3770 870 3810
rect 870 3770 880 3810
rect 820 3760 880 3770
rect 820 3730 880 3740
rect 820 3690 830 3730
rect 830 3690 870 3730
rect 870 3690 880 3730
rect 820 3680 880 3690
rect -557 3622 -505 3632
rect -557 3588 -547 3622
rect -547 3588 -513 3622
rect -513 3588 -505 3622
rect -557 3580 -505 3588
rect -197 3622 -145 3632
rect -197 3588 -187 3622
rect -187 3588 -153 3622
rect -153 3588 -145 3622
rect -197 3580 -145 3588
rect -77 3622 -25 3632
rect -77 3588 -67 3622
rect -67 3588 -33 3622
rect -33 3588 -25 3622
rect -77 3580 -25 3588
rect 283 3622 335 3632
rect 283 3588 293 3622
rect 293 3588 327 3622
rect 327 3588 335 3622
rect 283 3580 335 3588
rect 403 3622 455 3632
rect 403 3588 413 3622
rect 413 3588 447 3622
rect 447 3588 455 3622
rect 403 3580 455 3588
rect 820 3650 880 3660
rect 820 3610 830 3650
rect 830 3610 870 3650
rect 870 3610 880 3650
rect 820 3600 880 3610
rect -1240 3470 -1180 3530
rect -490 3470 -430 3530
rect -270 3470 -210 3530
rect -10 3470 50 3530
rect 210 3470 270 3530
rect 470 3470 530 3530
rect -1060 3360 -1000 3420
rect -1060 3280 -1000 3340
rect -1060 3250 -1000 3260
rect -1060 3210 -1050 3250
rect -1050 3210 -1010 3250
rect -1010 3210 -1000 3250
rect -1060 3200 -1000 3210
rect -820 3360 -760 3420
rect -820 3280 -760 3340
rect -820 3250 -760 3260
rect -820 3210 -810 3250
rect -810 3210 -770 3250
rect -770 3210 -760 3250
rect -820 3200 -760 3210
rect -580 3360 -520 3420
rect -580 3280 -520 3340
rect -580 3250 -520 3260
rect -580 3210 -570 3250
rect -570 3210 -530 3250
rect -530 3210 -520 3250
rect -580 3200 -520 3210
rect -340 3360 -280 3420
rect -340 3280 -280 3340
rect -340 3250 -280 3260
rect -340 3210 -330 3250
rect -330 3210 -290 3250
rect -290 3210 -280 3250
rect -340 3200 -280 3210
rect 300 3360 360 3420
rect 300 3280 360 3340
rect 300 3250 360 3260
rect 300 3210 310 3250
rect 310 3210 350 3250
rect 350 3210 360 3250
rect 300 3200 360 3210
rect 540 3360 600 3420
rect 540 3280 600 3340
rect 540 3250 600 3260
rect 540 3210 550 3250
rect 550 3210 590 3250
rect 590 3210 600 3250
rect 540 3200 600 3210
rect 780 3360 840 3420
rect 780 3280 840 3340
rect 780 3250 840 3260
rect 780 3210 790 3250
rect 790 3210 830 3250
rect 830 3210 840 3250
rect 780 3200 840 3210
rect 1180 3760 1240 3820
rect 1260 3760 1320 3820
rect 1340 3760 1400 3820
rect 1180 3680 1240 3740
rect 1260 3680 1320 3740
rect 1340 3680 1400 3740
rect 1180 3600 1240 3660
rect 1260 3600 1320 3660
rect 1340 3600 1400 3660
rect -80 2610 -20 2620
rect -80 2570 -70 2610
rect -70 2570 -30 2610
rect -30 2570 -20 2610
rect -80 2560 -20 2570
rect -80 2480 -20 2540
rect -80 2400 -20 2460
rect 1700 4750 1760 4810
rect 2420 4750 2480 4810
rect 2180 4460 2240 4470
rect 2180 4420 2190 4460
rect 2190 4420 2230 4460
rect 2230 4420 2240 4460
rect 2180 4410 2240 4420
rect 3140 4750 3200 4810
rect 2900 4460 2960 4470
rect 2900 4420 2910 4460
rect 2910 4420 2950 4460
rect 2950 4420 2960 4460
rect 2900 4410 2960 4420
rect 1760 4290 1820 4350
rect 1760 4210 1820 4270
rect 1760 4130 1820 4190
rect 1940 4290 2000 4350
rect 1940 4210 2000 4270
rect 1940 4130 2000 4190
rect 2180 4290 2240 4350
rect 2180 4210 2240 4270
rect 2180 4130 2240 4190
rect 2420 4290 2480 4350
rect 2420 4210 2480 4270
rect 2420 4130 2480 4190
rect 2660 4290 2720 4350
rect 2660 4210 2720 4270
rect 2660 4130 2720 4190
rect 2180 4020 2240 4080
rect 2660 4020 2720 4080
rect 1940 3910 2000 3970
rect 1700 3810 1760 3820
rect 1700 3770 1710 3810
rect 1710 3770 1750 3810
rect 1750 3770 1760 3810
rect 1700 3760 1760 3770
rect 2022 3852 2074 3860
rect 2022 3818 2032 3852
rect 2032 3818 2066 3852
rect 2066 3818 2074 3852
rect 2022 3808 2074 3818
rect 2420 3910 2480 3970
rect 2346 3852 2398 3860
rect 2346 3818 2356 3852
rect 2356 3818 2390 3852
rect 2390 3818 2398 3852
rect 2346 3808 2398 3818
rect 2500 3852 2552 3860
rect 2500 3818 2510 3852
rect 2510 3818 2544 3852
rect 2544 3818 2552 3852
rect 2500 3808 2552 3818
rect 4170 5460 4230 5520
rect 3980 5020 4040 5080
rect 3980 4940 4040 5000
rect 3980 4860 4040 4920
rect 3860 4750 3920 4810
rect 3620 4460 3680 4470
rect 3620 4420 3630 4460
rect 3630 4420 3670 4460
rect 3670 4420 3680 4460
rect 3620 4410 3680 4420
rect 3140 4290 3200 4350
rect 3140 4210 3200 4270
rect 3140 4130 3200 4190
rect 3380 4290 3440 4350
rect 3380 4210 3440 4270
rect 3380 4130 3440 4190
rect 3800 4290 3860 4350
rect 3800 4210 3860 4270
rect 3800 4130 3860 4190
rect 3140 4020 3200 4080
rect 2900 3910 2960 3970
rect 2824 3852 2876 3860
rect 2824 3818 2834 3852
rect 2834 3818 2868 3852
rect 2868 3818 2876 3852
rect 2824 3808 2876 3818
rect 2982 3852 3034 3860
rect 2982 3818 2992 3852
rect 2992 3818 3026 3852
rect 3026 3818 3034 3852
rect 2982 3808 3034 3818
rect 1700 3730 1760 3740
rect 1700 3690 1710 3730
rect 1710 3690 1750 3730
rect 1750 3690 1760 3730
rect 1700 3680 1760 3690
rect 1700 3650 1760 3660
rect 1700 3610 1710 3650
rect 1710 3610 1750 3650
rect 1750 3610 1760 3650
rect 1700 3600 1760 3610
rect 2125 3622 2177 3632
rect 2125 3588 2133 3622
rect 2133 3588 2167 3622
rect 2167 3588 2177 3622
rect 2125 3580 2177 3588
rect 2245 3622 2297 3632
rect 2245 3588 2253 3622
rect 2253 3588 2287 3622
rect 2287 3588 2297 3622
rect 2245 3580 2297 3588
rect 2605 3622 2657 3632
rect 2605 3588 2613 3622
rect 2613 3588 2647 3622
rect 2647 3588 2657 3622
rect 2605 3580 2657 3588
rect 2725 3622 2777 3632
rect 2725 3588 2733 3622
rect 2733 3588 2767 3622
rect 2767 3588 2777 3622
rect 2725 3580 2777 3588
rect 4260 5350 4320 5410
rect 8660 9940 8720 10000
rect 8000 9290 8060 9350
rect 7160 9170 7220 9230
rect 8980 9940 9040 10000
rect 9300 9940 9360 10000
rect 9740 9940 9800 10000
rect 8440 9290 8500 9350
rect 8880 9290 8940 9350
rect 10180 9940 10240 10000
rect 8220 9170 8280 9230
rect 7800 8950 7860 9010
rect 7360 8100 7420 8160
rect 7580 8100 7640 8160
rect 8020 8100 8080 8160
rect 8340 8100 8400 8160
rect 9390 9310 9450 9320
rect 9390 9270 9400 9310
rect 9400 9270 9440 9310
rect 9440 9270 9450 9310
rect 9390 9260 9450 9270
rect 9520 9290 9580 9350
rect 10400 9940 10460 10000
rect 9960 9290 10020 9350
rect 9390 9060 9450 9120
rect 10090 9310 10150 9320
rect 10090 9270 10100 9310
rect 10100 9270 10140 9310
rect 10140 9270 10150 9310
rect 10090 9260 10150 9270
rect 10770 9270 10840 9340
rect 9960 9010 10020 9070
rect 9830 8810 9890 8820
rect 9830 8770 9840 8810
rect 9840 8770 9880 8810
rect 9880 8770 9890 8810
rect 9830 8760 9890 8770
rect 8660 8100 8720 8160
rect 9100 8100 9160 8160
rect 9420 8100 9480 8160
rect 14020 9010 14080 9070
rect 10090 8810 10150 8820
rect 10090 8770 10100 8810
rect 10100 8770 10140 8810
rect 10140 8770 10150 8810
rect 10090 8760 10150 8770
rect 10770 8740 10840 8810
rect 9740 8100 9800 8160
rect 10180 8100 10240 8160
rect 10400 8100 10460 8160
rect 11120 7950 11190 8020
rect 7160 7830 7220 7890
rect 13910 7830 13970 7890
rect 6940 5080 7000 5140
rect 7050 7720 7110 7780
rect 7050 7640 7110 7700
rect 7050 7560 7110 7620
rect 11240 7200 11300 7260
rect 11030 6730 11090 6740
rect 11030 6690 11040 6730
rect 11040 6690 11080 6730
rect 11080 6690 11090 6730
rect 11030 6680 11090 6690
rect 7050 4920 7110 4980
rect 5590 4750 5650 4810
rect 4370 4290 4430 4350
rect 4450 4290 4510 4350
rect 4530 4290 4590 4350
rect 4370 4210 4430 4270
rect 4450 4210 4510 4270
rect 4530 4210 4590 4270
rect 4370 4130 4430 4190
rect 4450 4130 4510 4190
rect 4530 4130 4590 4190
rect 4260 3810 4320 3870
rect 3085 3622 3137 3632
rect 3085 3588 3093 3622
rect 3093 3588 3127 3622
rect 3127 3588 3137 3622
rect 3085 3580 3137 3588
rect 4170 3580 4230 3640
rect 2050 3470 2110 3530
rect 2310 3470 2370 3530
rect 2530 3470 2590 3530
rect 2790 3470 2850 3530
rect 3010 3470 3070 3530
rect 3760 3470 3820 3530
rect 1740 3360 1800 3420
rect 1740 3280 1800 3340
rect 1740 3250 1800 3260
rect 1740 3210 1750 3250
rect 1750 3210 1790 3250
rect 1790 3210 1800 3250
rect 1740 3200 1800 3210
rect 1980 3360 2040 3420
rect 1980 3280 2040 3340
rect 1980 3250 2040 3260
rect 1980 3210 1990 3250
rect 1990 3210 2030 3250
rect 2030 3210 2040 3250
rect 1980 3200 2040 3210
rect 2220 3360 2280 3420
rect 2220 3280 2280 3340
rect 2220 3250 2280 3260
rect 2220 3210 2230 3250
rect 2230 3210 2270 3250
rect 2270 3210 2280 3250
rect 2220 3200 2280 3210
rect 2860 3360 2920 3420
rect 2860 3280 2920 3340
rect 2860 3250 2920 3260
rect 2860 3210 2870 3250
rect 2870 3210 2910 3250
rect 2910 3210 2920 3250
rect 2860 3200 2920 3210
rect 3100 3360 3160 3420
rect 3100 3280 3160 3340
rect 3100 3250 3160 3260
rect 3100 3210 3110 3250
rect 3110 3210 3150 3250
rect 3150 3210 3160 3250
rect 3100 3200 3160 3210
rect 3340 3360 3400 3420
rect 3340 3280 3400 3340
rect 3340 3250 3400 3260
rect 3340 3210 3350 3250
rect 3350 3210 3390 3250
rect 3390 3210 3400 3250
rect 3340 3200 3400 3210
rect 3580 3360 3640 3420
rect 3580 3280 3640 3340
rect 3580 3250 3640 3260
rect 3580 3210 3590 3250
rect 3590 3210 3630 3250
rect 3630 3210 3640 3250
rect 3580 3200 3640 3210
rect 1180 2560 1240 2620
rect 1260 2560 1320 2620
rect 1340 2560 1400 2620
rect 1180 2480 1240 2540
rect 1260 2480 1320 2540
rect 1340 2480 1400 2540
rect 1180 2400 1240 2460
rect 1260 2400 1320 2460
rect 1340 2400 1400 2460
rect 2600 2610 2660 2620
rect 2600 2570 2610 2610
rect 2610 2570 2650 2610
rect 2650 2570 2660 2610
rect 2600 2560 2660 2570
rect 2600 2480 2660 2540
rect 2600 2400 2660 2460
rect -820 2340 -760 2350
rect -820 2300 -810 2340
rect -810 2300 -770 2340
rect -770 2300 -760 2340
rect -820 2290 -760 2300
rect -660 2340 -600 2350
rect -660 2300 -650 2340
rect -650 2300 -610 2340
rect -610 2300 -600 2340
rect -660 2290 -600 2300
rect -500 2340 -440 2350
rect -500 2300 -490 2340
rect -490 2300 -450 2340
rect -450 2300 -440 2340
rect -500 2290 -440 2300
rect -340 2340 -280 2350
rect -340 2300 -330 2340
rect -330 2300 -290 2340
rect -290 2300 -280 2340
rect -340 2290 -280 2300
rect -180 2340 -120 2350
rect -180 2300 -170 2340
rect -170 2300 -130 2340
rect -130 2300 -120 2340
rect -180 2290 -120 2300
rect -20 2340 40 2350
rect -20 2300 -10 2340
rect -10 2300 30 2340
rect 30 2300 40 2340
rect -20 2290 40 2300
rect 140 2340 200 2350
rect 140 2300 150 2340
rect 150 2300 190 2340
rect 190 2300 200 2340
rect 140 2290 200 2300
rect 300 2340 360 2350
rect 300 2300 310 2340
rect 310 2300 350 2340
rect 350 2300 360 2340
rect 300 2290 360 2300
rect 460 2340 520 2350
rect 460 2300 470 2340
rect 470 2300 510 2340
rect 510 2300 520 2340
rect 460 2290 520 2300
rect 620 2340 680 2350
rect 620 2300 630 2340
rect 630 2300 670 2340
rect 670 2300 680 2340
rect 620 2290 680 2300
rect 780 2340 840 2350
rect 780 2300 790 2340
rect 790 2300 830 2340
rect 830 2300 840 2340
rect 780 2290 840 2300
rect 940 2340 1000 2350
rect 940 2300 950 2340
rect 950 2300 990 2340
rect 990 2300 1000 2340
rect 940 2290 1000 2300
rect 1100 2340 1160 2350
rect 1100 2300 1110 2340
rect 1110 2300 1150 2340
rect 1150 2300 1160 2340
rect 1100 2290 1160 2300
rect 1260 2340 1320 2350
rect 1260 2300 1270 2340
rect 1270 2300 1310 2340
rect 1310 2300 1320 2340
rect 1260 2290 1320 2300
rect 1420 2340 1480 2350
rect 1420 2300 1430 2340
rect 1430 2300 1470 2340
rect 1470 2300 1480 2340
rect 1420 2290 1480 2300
rect 1580 2340 1640 2350
rect 1580 2300 1590 2340
rect 1590 2300 1630 2340
rect 1630 2300 1640 2340
rect 1580 2290 1640 2300
rect 1740 2340 1800 2350
rect 1740 2300 1750 2340
rect 1750 2300 1790 2340
rect 1790 2300 1800 2340
rect 1740 2290 1800 2300
rect 1900 2340 1960 2350
rect 1900 2300 1910 2340
rect 1910 2300 1950 2340
rect 1950 2300 1960 2340
rect 1900 2290 1960 2300
rect 2060 2340 2120 2350
rect 2060 2300 2070 2340
rect 2070 2300 2110 2340
rect 2110 2300 2120 2340
rect 2060 2290 2120 2300
rect 2220 2340 2280 2350
rect 2220 2300 2230 2340
rect 2230 2300 2270 2340
rect 2270 2300 2280 2340
rect 2220 2290 2280 2300
rect 2380 2340 2440 2350
rect 2380 2300 2390 2340
rect 2390 2300 2430 2340
rect 2430 2300 2440 2340
rect 2380 2290 2440 2300
rect 2540 2340 2600 2350
rect 2540 2300 2550 2340
rect 2550 2300 2590 2340
rect 2590 2300 2600 2340
rect 2540 2290 2600 2300
rect 2700 2340 2760 2350
rect 2700 2300 2710 2340
rect 2710 2300 2750 2340
rect 2750 2300 2760 2340
rect 2700 2290 2760 2300
rect 2860 2340 2920 2350
rect 2860 2300 2870 2340
rect 2870 2300 2910 2340
rect 2910 2300 2920 2340
rect 2860 2290 2920 2300
rect 3020 2340 3080 2350
rect 3020 2300 3030 2340
rect 3030 2300 3070 2340
rect 3070 2300 3080 2340
rect 3020 2290 3080 2300
rect 3180 2340 3240 2350
rect 3180 2300 3190 2340
rect 3190 2300 3230 2340
rect 3230 2300 3240 2340
rect 3180 2290 3240 2300
rect -900 2170 -840 2180
rect -900 2130 -890 2170
rect -890 2130 -850 2170
rect -850 2130 -840 2170
rect -900 2120 -840 2130
rect 3490 2210 3550 2220
rect 3490 2170 3500 2210
rect 3500 2170 3540 2210
rect 3540 2170 3550 2210
rect 3490 2160 3550 2170
rect 3490 2130 3550 2140
rect 3490 2090 3500 2130
rect 3500 2090 3540 2130
rect 3540 2090 3550 2130
rect 3490 2080 3550 2090
rect -1360 1950 -1300 2010
rect -950 1950 -890 2010
rect -2300 1840 -2240 1900
rect -1630 1610 -1570 1670
rect -3530 -1713 -3470 -1710
rect -3530 -2110 -3520 -1713
rect -3520 -2110 -3482 -1713
rect -3482 -2110 -3470 -1713
rect -3110 -1780 -3050 -1720
rect -3110 -1860 -3050 -1800
rect -3110 -1950 -3050 -1890
rect -3110 -2040 -3050 -1980
rect -3110 -2120 -3050 -2060
rect -3530 -2590 -3470 -2530
rect -3530 -2670 -3470 -2610
rect -3530 -2750 -3470 -2690
rect -2740 -2590 -2680 -2530
rect -2740 -2670 -2680 -2610
rect -2740 -2750 -2680 -2690
rect -1300 -2590 -1240 -2530
rect -1300 -2670 -1240 -2610
rect -1300 -2750 -1240 -2690
rect -3110 -2860 -3050 -2800
rect -840 1720 -780 1780
rect 562 1780 632 1790
rect 562 1730 572 1780
rect 572 1730 622 1780
rect 622 1730 632 1780
rect 562 1720 632 1730
rect 1960 1780 2030 1790
rect 1960 1730 1970 1780
rect 1970 1730 2020 1780
rect 2020 1730 2030 1780
rect 1960 1720 2030 1730
rect 4170 1730 4230 1790
rect 1970 1610 2030 1670
rect 3360 1530 3420 1590
rect -840 -480 -780 -420
rect -410 -480 -350 -420
rect 1260 -424 1264 -420
rect 1264 -424 1320 -420
rect 1260 -480 1320 -424
rect 4020 1530 4080 1590
rect 4260 1530 4320 1590
rect 4370 980 4430 1040
rect 4450 980 4510 1040
rect 4530 980 4590 1040
rect 4800 1840 4860 1900
rect 3360 -480 3420 -420
rect 7420 5560 7480 5620
rect 7620 5560 7680 5620
rect 7860 5610 7920 5620
rect 7860 5570 7870 5610
rect 7870 5570 7910 5610
rect 7910 5570 7920 5610
rect 7860 5560 7920 5570
rect 8020 5560 8080 5620
rect 8420 5560 8480 5620
rect 8820 5560 8880 5620
rect 9000 5720 9060 5730
rect 9000 5680 9010 5720
rect 9010 5680 9050 5720
rect 9050 5680 9060 5720
rect 9000 5670 9060 5680
rect 9220 5560 9280 5620
rect 9420 5560 9480 5620
rect 10140 5610 10200 5620
rect 10140 5570 10150 5610
rect 10150 5570 10190 5610
rect 10190 5570 10200 5610
rect 10140 5560 10200 5570
rect 9000 5500 9060 5510
rect 9000 5460 9010 5500
rect 9010 5460 9050 5500
rect 9050 5460 9060 5500
rect 9000 5450 9060 5460
rect 7640 4880 7700 4890
rect 7640 4840 7650 4880
rect 7650 4840 7690 4880
rect 7690 4840 7700 4880
rect 7640 4830 7700 4840
rect 8780 5220 8840 5230
rect 8780 5180 8790 5220
rect 8790 5180 8830 5220
rect 8830 5180 8840 5220
rect 8780 5170 8840 5180
rect 8080 5100 8140 5160
rect 7990 5000 8050 5060
rect 8740 4920 8800 4980
rect 9220 5220 9280 5230
rect 9220 5180 9230 5220
rect 9230 5180 9270 5220
rect 9270 5180 9280 5220
rect 9220 5170 9280 5180
rect 10760 5220 10820 5230
rect 10760 5180 10770 5220
rect 10770 5180 10810 5220
rect 10810 5180 10820 5220
rect 10760 5170 10820 5180
rect 11470 5260 11540 5330
rect 11240 5170 11300 5230
rect 9920 5100 9980 5110
rect 9920 5060 9930 5100
rect 9930 5060 9970 5100
rect 9970 5060 9980 5100
rect 9920 5050 9980 5060
rect 11630 5050 11690 5060
rect 11630 5010 11640 5050
rect 11640 5010 11680 5050
rect 11680 5010 11690 5050
rect 11630 5000 11690 5010
rect 13910 5000 13970 5060
rect 14020 7720 14080 7780
rect 14020 7640 14080 7700
rect 14020 7560 14080 7620
rect 8080 4880 8140 4890
rect 8080 4840 8090 4880
rect 8090 4840 8130 4880
rect 8130 4840 8140 4880
rect 8080 4830 8140 4840
rect 9150 4850 9210 4910
rect 9920 4880 9980 4890
rect 9920 4840 9930 4880
rect 9930 4840 9970 4880
rect 9970 4840 9980 4880
rect 9920 4830 9980 4840
rect 10760 4880 10820 4890
rect 10760 4840 10770 4880
rect 10770 4840 10810 4880
rect 10810 4840 10820 4880
rect 10760 4830 10820 4840
rect 11240 4830 11300 4890
rect 7940 4500 8000 4510
rect 7940 4460 7950 4500
rect 7950 4460 7990 4500
rect 7990 4460 8000 4500
rect 7940 4450 8000 4460
rect 7540 4340 7600 4400
rect 7740 4340 7800 4400
rect 7940 4200 8000 4260
rect 8140 4340 8200 4400
rect 8540 4340 8600 4400
rect 7160 3540 7220 3600
rect 8940 4340 9000 4400
rect 9020 4390 9080 4400
rect 9020 4350 9030 4390
rect 9030 4350 9070 4390
rect 9070 4350 9080 4390
rect 9020 4340 9080 4350
rect 9340 4340 9400 4400
rect 8340 3590 8400 3600
rect 8340 3550 8350 3590
rect 8350 3550 8390 3590
rect 8390 3550 8400 3590
rect 8340 3540 8400 3550
rect 9140 4200 9200 4260
rect 9540 4340 9600 4400
rect 10140 4390 10200 4400
rect 10140 4350 10150 4390
rect 10150 4350 10190 4390
rect 10190 4350 10200 4390
rect 10140 4340 10200 4350
rect 11470 4750 11540 4820
rect 8740 3590 8800 3600
rect 8740 3550 8750 3590
rect 8750 3550 8790 3590
rect 8790 3550 8800 3590
rect 8740 3540 8800 3550
rect 11030 3200 11090 3210
rect 11030 3160 11040 3200
rect 11040 3160 11080 3200
rect 11080 3160 11090 3200
rect 11030 3150 11090 3160
rect 6090 2910 6150 2970
rect 6190 2910 6250 2970
rect 5590 -420 5650 -360
rect 5970 280 6030 340
rect 1260 -2540 1320 -2530
rect 1260 -2580 1270 -2540
rect 1270 -2580 1310 -2540
rect 1310 -2580 1320 -2540
rect 1260 -2590 1320 -2580
rect 1260 -2620 1320 -2610
rect 1260 -2660 1270 -2620
rect 1270 -2660 1310 -2620
rect 1310 -2660 1320 -2620
rect 1260 -2670 1320 -2660
rect 1260 -2700 1320 -2690
rect 1260 -2740 1270 -2700
rect 1270 -2740 1310 -2700
rect 1310 -2740 1320 -2700
rect 1260 -2750 1320 -2740
rect 3690 -2590 3750 -2530
rect 3690 -2670 3750 -2610
rect 3690 -2750 3750 -2690
rect 5590 -1713 5650 -1710
rect 5590 -2110 5600 -1713
rect 5600 -2110 5638 -1713
rect 5638 -2110 5650 -1713
rect 11240 2820 11300 2880
rect 6140 -1120 6200 -1060
rect 6670 1950 6730 2010
rect 5970 -1780 6030 -1720
rect 6810 980 6870 1040
rect 6810 -420 6870 -360
rect 5970 -1860 6030 -1800
rect 6670 -1820 6730 -1760
rect 5970 -1950 6030 -1890
rect 5970 -2040 6030 -1980
rect 5970 -2120 6030 -2060
rect 4800 -2590 4860 -2530
rect 4800 -2670 4860 -2610
rect 4800 -2750 4860 -2690
rect 5590 -2590 5650 -2530
rect 5590 -2670 5650 -2610
rect 5590 -2750 5650 -2690
rect 6210 -2520 6270 -2460
rect 6210 -2860 6270 -2800
rect 3010 -3122 3420 -3110
rect 3010 -3160 3020 -3122
rect 3020 -3160 3417 -3122
rect 3417 -3160 3420 -3122
rect 3010 -3170 3420 -3160
rect 4920 -3122 5330 -3110
rect 4920 -3160 4923 -3122
rect 4923 -3160 5320 -3122
rect 5320 -3160 5330 -3122
rect 4920 -3170 5330 -3160
rect 14020 -3170 14080 -3110
rect 4140 -3310 4200 -3300
rect 4140 -3350 4150 -3310
rect 4150 -3350 4190 -3310
rect 4190 -3350 4200 -3310
rect 4140 -3360 4200 -3350
<< metal2 >>
rect 10600 14880 10700 14920
rect 10600 14820 10620 14880
rect 10680 14840 10700 14880
rect 10680 14830 12930 14840
rect 10680 14820 11330 14830
rect 10600 14780 11330 14820
rect 10600 14720 10620 14780
rect 10680 14770 11330 14780
rect 11390 14770 11850 14830
rect 11910 14770 12370 14830
rect 12430 14770 12860 14830
rect 12920 14770 12930 14830
rect 10680 14760 12930 14770
rect 10680 14720 10700 14760
rect 10600 14680 10700 14720
rect 10820 14720 13420 14730
rect 10820 14660 10830 14720
rect 10890 14660 10910 14720
rect 10970 14660 10990 14720
rect 11050 14660 13190 14720
rect 13250 14660 13270 14720
rect 13330 14660 13350 14720
rect 13410 14660 13420 14720
rect 10820 14640 13420 14660
rect 10820 14580 10830 14640
rect 10890 14580 10910 14640
rect 10970 14580 10990 14640
rect 11050 14580 13190 14640
rect 13250 14580 13270 14640
rect 13330 14580 13350 14640
rect 13410 14580 13420 14640
rect 10820 14560 13420 14580
rect 10820 14500 10830 14560
rect 10890 14500 10910 14560
rect 10970 14500 10990 14560
rect 11050 14500 13190 14560
rect 13250 14500 13270 14560
rect 13330 14500 13350 14560
rect 13410 14500 13420 14560
rect 10820 14490 13420 14500
rect 11275 14112 14090 14120
rect 11275 14060 11280 14112
rect 11332 14060 11800 14112
rect 11852 14060 12320 14112
rect 12372 14060 12886 14112
rect 12938 14110 14090 14112
rect 12938 14060 14020 14110
rect 11275 14050 14020 14060
rect 14080 14050 14090 14110
rect 11330 13750 11610 13760
rect 11390 13690 11540 13750
rect 11600 13690 11610 13750
rect 11330 13680 11610 13690
rect 11850 13750 12130 13760
rect 11910 13690 12060 13750
rect 12120 13690 12130 13750
rect 11850 13680 12130 13690
rect 12370 13750 12650 13760
rect 12430 13690 12580 13750
rect 12640 13690 12650 13750
rect 12370 13680 12650 13690
rect 11290 13632 11500 13640
rect 11290 13580 11294 13632
rect 11346 13630 11500 13632
rect 11346 13580 11430 13630
rect 11290 13570 11430 13580
rect 11490 13570 11500 13630
rect 11810 13632 12020 13640
rect 11810 13580 11814 13632
rect 11866 13630 12020 13632
rect 11866 13580 11950 13630
rect 11810 13570 11950 13580
rect 12010 13570 12020 13630
rect 12330 13632 12540 13640
rect 12330 13580 12334 13632
rect 12386 13630 12540 13632
rect 12386 13580 12470 13630
rect 12330 13570 12470 13580
rect 12530 13570 12540 13630
rect 11420 13560 11500 13570
rect 11940 13560 12020 13570
rect 12460 13560 12540 13570
rect 230 13480 330 13520
rect 230 13420 250 13480
rect 310 13440 330 13480
rect 310 13430 10630 13440
rect 310 13420 560 13430
rect 230 13380 560 13420
rect 230 13320 250 13380
rect 310 13370 560 13380
rect 620 13370 780 13430
rect 840 13370 1250 13430
rect 1310 13370 1590 13430
rect 1650 13370 1810 13430
rect 1870 13370 2250 13430
rect 2310 13370 2930 13430
rect 2990 13370 3150 13430
rect 3210 13370 3620 13430
rect 3680 13370 4080 13430
rect 4140 13370 4430 13430
rect 4490 13370 4680 13430
rect 4740 13370 4900 13430
rect 4960 13370 5230 13430
rect 5290 13370 5890 13430
rect 5950 13370 6110 13430
rect 6170 13370 6680 13430
rect 6740 13370 6940 13430
rect 7000 13370 7190 13430
rect 7250 13370 7410 13430
rect 7470 13370 7960 13430
rect 8020 13370 8240 13430
rect 8300 13370 8490 13430
rect 8550 13370 8710 13430
rect 8770 13370 9260 13430
rect 9320 13370 9540 13430
rect 9600 13370 9790 13430
rect 9850 13370 10010 13430
rect 10070 13370 10560 13430
rect 10620 13370 10630 13430
rect 310 13360 10630 13370
rect 310 13320 330 13360
rect 230 13280 330 13320
rect 10820 13140 11320 13150
rect 10820 13080 10830 13140
rect 10890 13080 10910 13140
rect 10970 13080 10990 13140
rect 11050 13080 11260 13140
rect 10820 13070 11320 13080
rect 10762 13060 11320 13070
rect 120 13050 410 13060
rect 120 12990 130 13050
rect 190 12990 340 13050
rect 400 12990 410 13050
rect 10762 13052 10830 13060
rect 10762 13000 10766 13052
rect 10818 13000 10830 13052
rect 10890 13000 10910 13060
rect 10970 13000 10990 13060
rect 11050 13000 11260 13060
rect 10762 12990 11320 13000
rect 120 12980 410 12990
rect 10820 12980 11320 12990
rect 10820 12920 10830 12980
rect 10890 12920 10910 12980
rect 10970 12920 10990 12980
rect 11050 12920 11260 12980
rect 10820 12910 11320 12920
rect 11350 13140 11840 13150
rect 11410 13080 11780 13140
rect 11350 13060 11840 13080
rect 11410 13000 11780 13060
rect 11350 12980 11840 13000
rect 11410 12920 11780 12980
rect 11350 12910 11840 12920
rect 11870 13140 12360 13150
rect 11930 13080 12300 13140
rect 11870 13060 12360 13080
rect 11930 13000 12300 13060
rect 11870 12980 12360 13000
rect 11930 12920 12300 12980
rect 11870 12910 12360 12920
rect 12390 13140 13420 13150
rect 12450 13080 13190 13140
rect 13250 13080 13270 13140
rect 13330 13080 13350 13140
rect 13410 13080 13420 13140
rect 12390 13060 13420 13080
rect 12450 13000 13190 13060
rect 13250 13000 13270 13060
rect 13330 13000 13350 13060
rect 13410 13000 13420 13060
rect 12390 12980 13420 13000
rect 12450 12920 13190 12980
rect 13250 12920 13270 12980
rect 13330 12920 13350 12980
rect 13410 12920 13420 12980
rect 12390 12910 13420 12920
rect 230 12700 330 12740
rect 230 12640 250 12700
rect 310 12660 330 12700
rect 310 12650 10630 12660
rect 310 12640 720 12650
rect 230 12600 720 12640
rect 230 12540 250 12600
rect 310 12590 720 12600
rect 780 12590 1140 12650
rect 1200 12590 1810 12650
rect 1870 12590 2380 12650
rect 2440 12590 3090 12650
rect 3150 12590 3520 12650
rect 3580 12590 3960 12650
rect 4020 12590 4210 12650
rect 4270 12590 4430 12650
rect 4490 12590 4900 12650
rect 4960 12590 5340 12650
rect 5400 12590 5960 12650
rect 6020 12590 6300 12650
rect 6360 12590 6660 12650
rect 6720 12590 7260 12650
rect 7320 12590 7600 12650
rect 7660 12590 7960 12650
rect 8020 12590 8560 12650
rect 8620 12590 8900 12650
rect 8960 12590 9260 12650
rect 9320 12590 9860 12650
rect 9920 12590 10200 12650
rect 10260 12590 10560 12650
rect 10620 12590 10630 12650
rect 310 12580 10630 12590
rect 310 12540 330 12580
rect 230 12500 330 12540
rect 11530 12290 11610 12300
rect 12050 12290 12130 12300
rect 12570 12290 12650 12300
rect 11290 12282 11540 12290
rect 11290 12230 11294 12282
rect 11346 12230 11540 12282
rect 11600 12230 11610 12290
rect 11290 12220 11610 12230
rect 11810 12282 12060 12290
rect 11810 12230 11814 12282
rect 11866 12230 12060 12282
rect 12120 12230 12130 12290
rect 11810 12220 12130 12230
rect 12330 12282 12580 12290
rect 12330 12230 12334 12282
rect 12386 12230 12580 12282
rect 12640 12230 12650 12290
rect 12330 12220 12650 12230
rect 11330 12170 11500 12180
rect 11390 12110 11430 12170
rect 11490 12110 11500 12170
rect 11330 12100 11500 12110
rect 11850 12170 12020 12180
rect 11910 12110 11950 12170
rect 12010 12110 12020 12170
rect 11850 12100 12020 12110
rect 12370 12170 12540 12180
rect 12430 12110 12470 12170
rect 12530 12110 12540 12170
rect 12370 12100 12540 12110
rect 11320 11580 11670 11590
rect 11320 11520 11330 11580
rect 11390 11520 11600 11580
rect 11660 11520 11670 11580
rect 11320 11510 11670 11520
rect 11840 11580 12190 11590
rect 11840 11520 11850 11580
rect 11910 11520 12120 11580
rect 12180 11520 12190 11580
rect 11840 11510 12190 11520
rect 12360 11580 12710 11590
rect 12360 11520 12370 11580
rect 12430 11520 12640 11580
rect 12700 11520 12710 11580
rect 12360 11510 12710 11520
rect 11400 11400 13030 11410
rect 11400 11340 11410 11400
rect 11470 11340 11930 11400
rect 11990 11340 12450 11400
rect 12510 11340 12780 11400
rect 12840 11340 12970 11400
rect 11400 11330 13030 11340
rect 10600 10800 10700 10840
rect 10600 10740 10620 10800
rect 10680 10760 10700 10800
rect 10680 10750 13230 10760
rect 10680 10740 11600 10750
rect 10600 10700 11600 10740
rect 10600 10640 10620 10700
rect 10680 10690 11600 10700
rect 11660 10690 12120 10750
rect 12180 10690 12640 10750
rect 12700 10690 13160 10750
rect 13220 10690 13230 10750
rect 10680 10680 13230 10690
rect 10680 10640 10700 10680
rect 10600 10600 10700 10640
rect 920 10500 1020 10540
rect 10990 10520 11100 10540
rect 920 10440 940 10500
rect 1000 10460 1020 10500
rect 5700 10510 11010 10520
rect 1000 10450 5260 10460
rect 1000 10440 1270 10450
rect 920 10400 1270 10440
rect 920 10340 940 10400
rect 1000 10390 1270 10400
rect 1330 10390 1490 10450
rect 1550 10390 1790 10450
rect 1850 10390 2010 10450
rect 2070 10390 2170 10450
rect 2230 10390 2390 10450
rect 2450 10390 2690 10450
rect 2750 10390 2910 10450
rect 2970 10390 3210 10450
rect 3270 10390 3650 10450
rect 3710 10390 3980 10450
rect 4040 10390 4410 10450
rect 4470 10390 4800 10450
rect 4860 10390 5190 10450
rect 5250 10390 5260 10450
rect 5700 10450 5710 10510
rect 5770 10450 11010 10510
rect 11080 10450 11100 10520
rect 5700 10440 11100 10450
rect 10990 10430 11100 10440
rect 1000 10380 5260 10390
rect 1000 10340 1020 10380
rect 920 10300 1020 10340
rect 1670 10340 1750 10350
rect 1670 10280 1680 10340
rect 1740 10310 1750 10340
rect 3390 10340 3470 10350
rect 3390 10310 3400 10340
rect 1740 10280 3400 10310
rect 3460 10310 3470 10340
rect 5470 10340 6490 10350
rect 4240 10320 4320 10330
rect 4240 10310 4250 10320
rect 3460 10280 4250 10310
rect 1670 10270 4250 10280
rect 4240 10260 4250 10270
rect 4310 10260 4320 10320
rect 5470 10280 5480 10340
rect 5540 10280 6420 10340
rect 6480 10280 6490 10340
rect 5470 10270 6490 10280
rect 4240 10250 4320 10260
rect 6010 10000 6380 10010
rect 3040 9990 3120 10000
rect 10 9960 1220 9970
rect 10 9900 1150 9960
rect 1210 9900 1220 9960
rect 3040 9930 3050 9990
rect 3110 9930 3120 9990
rect 3040 9920 3120 9930
rect 4130 9950 4210 9960
rect 10 9890 1220 9900
rect 4130 9890 4140 9950
rect 4200 9890 4210 9950
rect 6010 9940 6020 10000
rect 6080 9940 6310 10000
rect 6370 9940 6380 10000
rect 6010 9930 6380 9940
rect 7250 10000 10470 10010
rect 7250 9940 7290 10000
rect 7350 9940 7390 10000
rect 7450 9940 7560 10000
rect 7620 9940 7780 10000
rect 7840 9940 8220 10000
rect 8280 9940 8660 10000
rect 8720 9940 8980 10000
rect 9040 9940 9300 10000
rect 9360 9940 9740 10000
rect 9800 9940 10180 10000
rect 10240 9940 10400 10000
rect 10460 9940 10470 10000
rect 7250 9930 10470 9940
rect 4130 9880 4210 9890
rect 5700 9920 5780 9930
rect 5700 9860 5710 9920
rect 5770 9860 5780 9920
rect 5700 9850 5780 9860
rect 3260 9380 3340 9390
rect 920 9320 1020 9360
rect 3260 9320 3270 9380
rect 3330 9320 3340 9380
rect 6930 9350 8950 9360
rect 920 9260 940 9320
rect 1000 9280 1020 9320
rect 6930 9290 6940 9350
rect 7000 9290 8000 9350
rect 8060 9290 8440 9350
rect 8500 9290 8880 9350
rect 8940 9290 8950 9350
rect 9510 9350 10030 9360
rect 6930 9280 8950 9290
rect 9380 9320 9460 9330
rect 1000 9270 5940 9280
rect 1000 9260 1270 9270
rect 920 9220 1270 9260
rect 920 9160 940 9220
rect 1000 9210 1270 9220
rect 1330 9210 2010 9270
rect 2070 9210 2170 9270
rect 2230 9210 2910 9270
rect 2970 9210 3160 9270
rect 3220 9210 3350 9270
rect 3410 9210 3430 9270
rect 3490 9210 3640 9270
rect 3700 9210 3970 9270
rect 4030 9210 4410 9270
rect 4470 9210 4800 9270
rect 4860 9210 5010 9270
rect 5070 9210 5190 9270
rect 5250 9210 5870 9270
rect 5930 9210 5940 9270
rect 9380 9260 9390 9320
rect 9450 9260 9460 9320
rect 9510 9290 9520 9350
rect 9580 9290 9960 9350
rect 10020 9290 10030 9350
rect 10750 9340 10860 9360
rect 10750 9330 10770 9340
rect 9510 9280 10030 9290
rect 10080 9320 10770 9330
rect 9380 9250 9460 9260
rect 10080 9260 10090 9320
rect 10150 9270 10770 9320
rect 10840 9270 10860 9340
rect 10150 9260 10860 9270
rect 10080 9250 10860 9260
rect 1000 9200 5940 9210
rect 6410 9230 8290 9240
rect 1000 9160 1020 9200
rect 6410 9170 6420 9230
rect 6480 9170 7160 9230
rect 7220 9170 8220 9230
rect 8280 9170 8290 9230
rect 920 9120 1020 9160
rect 1710 9160 1790 9170
rect 1710 9100 1720 9160
rect 1780 9150 1790 9160
rect 3240 9160 3320 9170
rect 5470 9160 6270 9170
rect 6410 9160 8290 9170
rect 3240 9150 3250 9160
rect 1780 9110 3250 9150
rect 1780 9100 1790 9110
rect 1710 9090 1790 9100
rect 3240 9100 3250 9110
rect 3310 9140 3320 9160
rect 4240 9150 4320 9160
rect 4240 9140 4250 9150
rect 3310 9100 4250 9140
rect 3240 9090 3320 9100
rect 4240 9090 4250 9100
rect 4310 9090 4320 9150
rect 4660 9100 4670 9160
rect 4730 9150 4740 9160
rect 4830 9150 4840 9160
rect 4730 9110 4840 9150
rect 4730 9100 4740 9110
rect 4830 9100 4840 9110
rect 4900 9100 4910 9160
rect 4830 9090 4910 9100
rect 5470 9100 5480 9160
rect 5540 9100 6200 9160
rect 6260 9100 6270 9160
rect 5470 9090 6270 9100
rect 6300 9120 9460 9130
rect 4240 9080 4320 9090
rect 6300 9060 6310 9120
rect 6370 9060 9390 9120
rect 9450 9060 9460 9120
rect 6300 9050 9460 9060
rect 9950 9070 14090 9080
rect 6190 9010 7870 9020
rect 6190 8950 6200 9010
rect 6260 8950 6670 9010
rect 6730 8950 6750 9010
rect 6810 8950 6830 9010
rect 6890 8950 7800 9010
rect 7860 8950 7870 9010
rect 9950 9010 9960 9070
rect 10020 9010 14020 9070
rect 14080 9010 14090 9070
rect 9950 9000 14090 9010
rect 6190 8940 7870 8950
rect 6190 8900 9900 8910
rect 6190 8840 6200 8900
rect 6260 8840 9900 8900
rect 6190 8830 9900 8840
rect 9820 8820 9900 8830
rect 9820 8760 9830 8820
rect 9890 8760 9900 8820
rect 9820 8750 9900 8760
rect 10080 8820 10860 8830
rect 10080 8760 10090 8820
rect 10150 8810 10860 8820
rect 10150 8760 10770 8810
rect 10080 8750 10770 8760
rect 10750 8740 10770 8750
rect 10840 8740 10860 8810
rect 10750 8720 10860 8740
rect 3060 8590 3140 8600
rect 120 8580 1220 8590
rect 120 8520 130 8580
rect 190 8520 1150 8580
rect 1210 8520 1220 8580
rect 3060 8530 3070 8590
rect 3130 8530 3140 8590
rect 3060 8520 3140 8530
rect 4090 8590 4170 8600
rect 4090 8530 4100 8590
rect 4160 8530 4170 8590
rect 4090 8520 4170 8530
rect 6010 8540 6270 8550
rect 120 8510 1220 8520
rect 6010 8480 6020 8540
rect 6080 8480 6200 8540
rect 6260 8480 6270 8540
rect 6010 8470 6270 8480
rect 4910 8200 4990 8210
rect 920 8140 1020 8180
rect 920 8080 940 8140
rect 1000 8100 1020 8140
rect 4910 8140 4920 8200
rect 4980 8140 4990 8200
rect 4910 8130 4990 8140
rect 5540 8200 6190 8210
rect 5540 8140 5550 8200
rect 5610 8140 6120 8200
rect 6180 8140 6190 8200
rect 5540 8130 6190 8140
rect 6350 8160 10470 8170
rect 6350 8100 6390 8160
rect 6450 8100 6490 8160
rect 6550 8100 7360 8160
rect 7420 8100 7580 8160
rect 7640 8100 8020 8160
rect 8080 8100 8340 8160
rect 8400 8100 8660 8160
rect 8720 8100 9100 8160
rect 9160 8100 9420 8160
rect 9480 8100 9740 8160
rect 9800 8100 10180 8160
rect 10240 8100 10400 8160
rect 10460 8100 10470 8160
rect 1000 8090 5940 8100
rect 6350 8090 10470 8100
rect 1000 8080 1270 8090
rect 920 8040 1270 8080
rect 920 7980 940 8040
rect 1000 8030 1270 8040
rect 1330 8030 1490 8090
rect 1550 8030 1790 8090
rect 1850 8030 2020 8090
rect 2080 8030 2170 8090
rect 2230 8030 2390 8090
rect 2450 8030 2690 8090
rect 2750 8030 2910 8090
rect 2970 8030 3310 8090
rect 3370 8030 3640 8090
rect 3700 8030 3970 8090
rect 4030 8030 4410 8090
rect 4470 8030 4670 8090
rect 4730 8030 5190 8090
rect 5250 8030 5870 8090
rect 5930 8030 5940 8090
rect 11100 8030 11210 8040
rect 1000 8020 5940 8030
rect 6110 8020 11210 8030
rect 1000 7980 1020 8020
rect 920 7940 1020 7980
rect 6110 7960 6120 8020
rect 6180 7960 11120 8020
rect 6110 7950 11120 7960
rect 11190 7950 11210 8020
rect 11100 7930 11210 7950
rect 7150 7890 13980 7900
rect 7150 7830 7160 7890
rect 7220 7830 13910 7890
rect 13970 7830 13980 7890
rect 7150 7820 13980 7830
rect 7040 7780 14090 7790
rect 7040 7720 7050 7780
rect 7110 7720 14020 7780
rect 14080 7720 14090 7780
rect 7040 7700 14090 7720
rect 7040 7640 7050 7700
rect 7110 7640 14020 7700
rect 14080 7640 14090 7700
rect 7040 7620 14090 7640
rect 7040 7560 7050 7620
rect 7110 7560 14020 7620
rect 14080 7560 14090 7620
rect 7040 7550 14090 7560
rect 11220 7260 11320 7280
rect 1650 7250 6900 7260
rect 1650 7190 1660 7250
rect 1720 7190 1880 7250
rect 1940 7190 2100 7250
rect 2160 7190 2320 7250
rect 2380 7190 2540 7250
rect 2600 7190 2760 7250
rect 2820 7190 6670 7250
rect 6730 7190 6750 7250
rect 6810 7190 6830 7250
rect 6890 7190 6900 7250
rect 1650 7170 6900 7190
rect 11220 7200 11240 7260
rect 11300 7200 11320 7260
rect 11220 7180 11320 7200
rect 1650 7110 1660 7170
rect 1720 7110 1880 7170
rect 1940 7110 2100 7170
rect 2160 7110 2320 7170
rect 2380 7110 2540 7170
rect 2600 7110 2760 7170
rect 2820 7110 6670 7170
rect 6730 7110 6750 7170
rect 6810 7110 6830 7170
rect 6890 7110 6900 7170
rect 1650 7090 6900 7110
rect -2310 7080 930 7090
rect -2310 7020 -2300 7080
rect -2240 7020 -240 7080
rect -180 7020 -20 7080
rect 40 7020 200 7080
rect 260 7020 420 7080
rect 480 7020 640 7080
rect 700 7020 860 7080
rect 920 7020 930 7080
rect 1650 7030 1660 7090
rect 1720 7030 1880 7090
rect 1940 7030 2100 7090
rect 2160 7030 2320 7090
rect 2380 7030 2540 7090
rect 2600 7030 2760 7090
rect 2820 7030 6670 7090
rect 6730 7030 6750 7090
rect 6810 7030 6830 7090
rect 6890 7030 6900 7090
rect 1650 7020 6900 7030
rect -2310 7010 930 7020
rect 6050 6980 6290 6990
rect -360 6970 6290 6980
rect -360 6910 -350 6970
rect -290 6910 -130 6970
rect -70 6910 90 6970
rect 150 6910 310 6970
rect 370 6910 530 6970
rect 590 6910 750 6970
rect 810 6910 970 6970
rect 1030 6910 1550 6970
rect 1610 6910 1770 6970
rect 1830 6910 1990 6970
rect 2050 6910 2210 6970
rect 2270 6910 2430 6970
rect 2490 6910 2650 6970
rect 2710 6910 2870 6970
rect 2930 6910 6090 6970
rect 6150 6910 6190 6970
rect 6250 6910 6290 6970
rect -360 6900 6290 6910
rect 6050 6890 6290 6900
rect 6350 6740 11100 6750
rect 6350 6680 6390 6740
rect 6450 6680 6490 6740
rect 6550 6680 11030 6740
rect 11090 6680 11100 6740
rect 6350 6670 11100 6680
rect -3540 6632 2764 6640
rect -3540 6630 -182 6632
rect -3540 6570 -3530 6630
rect -3470 6580 -182 6630
rect -130 6580 -72 6632
rect -20 6580 38 6632
rect 90 6580 148 6632
rect 200 6580 258 6632
rect 310 6580 368 6632
rect 420 6580 478 6632
rect 530 6580 588 6632
rect 640 6580 698 6632
rect 750 6580 808 6632
rect 860 6580 1718 6632
rect 1770 6580 1828 6632
rect 1880 6580 1938 6632
rect 1990 6580 2048 6632
rect 2100 6580 2158 6632
rect 2210 6580 2268 6632
rect 2320 6580 2378 6632
rect 2430 6580 2488 6632
rect 2540 6580 2598 6632
rect 2650 6580 2708 6632
rect 2760 6580 2764 6632
rect -3470 6570 2764 6580
rect -370 6530 6290 6540
rect -370 6470 -360 6530
rect -300 6470 0 6530
rect 60 6470 360 6530
rect 420 6470 720 6530
rect 780 6470 1080 6530
rect 1140 6470 1440 6530
rect 1500 6470 1800 6530
rect 1860 6470 2160 6530
rect 2220 6470 2520 6530
rect 2580 6470 2880 6530
rect 2940 6470 3510 6530
rect 3570 6470 3950 6530
rect 4010 6500 6290 6530
rect 4010 6470 6090 6500
rect -370 6450 6090 6470
rect -370 6390 -360 6450
rect -300 6390 0 6450
rect 60 6390 360 6450
rect 420 6390 720 6450
rect 780 6390 1080 6450
rect 1140 6390 1440 6450
rect 1500 6390 1800 6450
rect 1860 6390 2160 6450
rect 2220 6390 2520 6450
rect 2580 6390 2880 6450
rect 2940 6390 3510 6450
rect 3570 6390 3950 6450
rect 4010 6440 6090 6450
rect 6150 6440 6190 6500
rect 6250 6440 6290 6500
rect 4010 6400 6290 6440
rect 4010 6390 6090 6400
rect -370 6370 6090 6390
rect -370 6310 -360 6370
rect -300 6310 0 6370
rect 60 6310 360 6370
rect 420 6310 720 6370
rect 780 6310 1080 6370
rect 1140 6310 1440 6370
rect 1500 6310 1800 6370
rect 1860 6310 2160 6370
rect 2220 6310 2520 6370
rect 2580 6310 2880 6370
rect 2940 6310 3510 6370
rect 3570 6310 3950 6370
rect 4010 6340 6090 6370
rect 6150 6340 6190 6400
rect 6250 6340 6290 6400
rect 4010 6310 6290 6340
rect -370 6300 6290 6310
rect 3250 6170 3330 6180
rect 3250 6110 3260 6170
rect 3320 6160 3330 6170
rect 3720 6170 3800 6180
rect 3720 6160 3730 6170
rect 3320 6120 3730 6160
rect 3320 6110 3330 6120
rect 3250 6100 3330 6110
rect 3720 6110 3730 6120
rect 3790 6110 3800 6170
rect 3720 6100 3800 6110
rect 3600 5830 3920 5840
rect 3600 5770 3610 5830
rect 3670 5770 3850 5830
rect 3910 5770 3920 5830
rect 3600 5760 3920 5770
rect 8990 5730 9070 5740
rect 8990 5670 9000 5730
rect 9060 5670 9070 5730
rect 8990 5660 9070 5670
rect -90 5630 2670 5640
rect -30 5570 90 5630
rect 150 5570 270 5630
rect 330 5570 450 5630
rect 510 5570 630 5630
rect 690 5570 810 5630
rect 870 5570 990 5630
rect 1050 5570 1170 5630
rect 1230 5570 1350 5630
rect 1410 5570 1440 5630
rect 1500 5570 1530 5630
rect 1590 5570 1710 5630
rect 1770 5570 1890 5630
rect 1950 5570 2070 5630
rect 2130 5570 2250 5630
rect 2310 5570 2430 5630
rect 2490 5570 2610 5630
rect -90 5560 2670 5570
rect 6350 5630 6590 5640
rect 6350 5620 10210 5630
rect 6350 5560 6390 5620
rect 6450 5560 6490 5620
rect 6550 5560 7420 5620
rect 7480 5560 7620 5620
rect 7680 5560 7860 5620
rect 7920 5560 8020 5620
rect 8080 5560 8420 5620
rect 8480 5560 8820 5620
rect 8880 5560 9220 5620
rect 9280 5560 9420 5620
rect 9480 5560 10140 5620
rect 10200 5560 10210 5620
rect 6350 5550 10210 5560
rect 6350 5540 6590 5550
rect 890 5520 4240 5530
rect 890 5460 900 5520
rect 960 5460 1620 5520
rect 1680 5460 4170 5520
rect 4230 5460 4240 5520
rect 890 5450 4240 5460
rect 8990 5510 9070 5520
rect 8990 5450 9000 5510
rect 9060 5450 9070 5510
rect 8990 5440 9070 5450
rect 530 5410 4330 5420
rect 530 5350 540 5410
rect 600 5350 1980 5410
rect 2040 5350 3260 5410
rect 3320 5350 4260 5410
rect 4320 5350 4330 5410
rect 530 5340 4330 5350
rect 11450 5330 11560 5350
rect -2530 5300 3800 5310
rect -2530 5240 -2520 5300
rect -2460 5240 180 5300
rect 240 5240 2340 5300
rect 2400 5240 3730 5300
rect 3790 5240 3800 5300
rect 11450 5260 11470 5330
rect 11540 5260 11560 5330
rect 11450 5240 11560 5260
rect -2530 5230 3800 5240
rect 8770 5230 8850 5240
rect -2420 5190 2770 5200
rect -2420 5130 -2410 5190
rect -2350 5130 -180 5190
rect -120 5130 1260 5190
rect 1320 5130 2700 5190
rect 2760 5130 2770 5190
rect 8770 5170 8780 5230
rect 8840 5170 8850 5230
rect 8070 5160 8150 5170
rect 8770 5160 8850 5170
rect 9210 5230 9290 5240
rect 9210 5170 9220 5230
rect 9280 5170 9290 5230
rect -2420 5120 2770 5130
rect 6930 5140 7010 5150
rect -1470 5080 6290 5090
rect -1470 5020 -1460 5080
rect -1400 5020 -1220 5080
rect -1160 5020 -980 5080
rect -920 5020 -740 5080
rect -680 5020 -500 5080
rect -440 5020 -260 5080
rect -200 5020 -20 5080
rect 40 5020 220 5080
rect 280 5020 460 5080
rect 520 5020 700 5080
rect 760 5020 940 5080
rect 1000 5020 1580 5080
rect 1640 5020 1820 5080
rect 1880 5020 2060 5080
rect 2120 5020 2300 5080
rect 2360 5020 2540 5080
rect 2600 5020 2780 5080
rect 2840 5020 3020 5080
rect 3080 5020 3260 5080
rect 3320 5020 3500 5080
rect 3560 5020 3740 5080
rect 3800 5020 3980 5080
rect 4040 5050 6290 5080
rect 6930 5080 6940 5140
rect 7000 5130 7010 5140
rect 8070 5130 8080 5160
rect 7000 5100 8080 5130
rect 8140 5130 8150 5160
rect 9210 5130 9290 5170
rect 10750 5230 11310 5240
rect 10750 5170 10760 5230
rect 10820 5170 11240 5230
rect 11300 5170 11310 5230
rect 10750 5160 11310 5170
rect 8140 5100 9290 5130
rect 7000 5090 9290 5100
rect 9910 5110 9990 5120
rect 7000 5080 7010 5090
rect 6930 5070 7010 5080
rect 4040 5020 6090 5050
rect -1470 5000 6090 5020
rect -1470 4940 -1460 5000
rect -1400 4940 -1220 5000
rect -1160 4940 -980 5000
rect -920 4940 -740 5000
rect -680 4940 -500 5000
rect -440 4940 -260 5000
rect -200 4940 -20 5000
rect 40 4940 220 5000
rect 280 4940 460 5000
rect 520 4940 700 5000
rect 760 4940 940 5000
rect 1000 4940 1580 5000
rect 1640 4940 1820 5000
rect 1880 4940 2060 5000
rect 2120 4940 2300 5000
rect 2360 4940 2540 5000
rect 2600 4940 2780 5000
rect 2840 4940 3020 5000
rect 3080 4940 3260 5000
rect 3320 4940 3500 5000
rect 3560 4940 3740 5000
rect 3800 4940 3980 5000
rect 4040 4990 6090 5000
rect 6150 4990 6190 5050
rect 6250 4990 6290 5050
rect 7980 5000 7990 5060
rect 8050 5050 8060 5060
rect 9910 5050 9920 5110
rect 9980 5050 9990 5110
rect 8050 5010 9990 5050
rect 11620 5060 13980 5070
rect 8050 5000 8060 5010
rect 11620 5000 11630 5060
rect 11690 5000 13910 5060
rect 13970 5000 13980 5060
rect 11620 4990 13980 5000
rect 4040 4950 6290 4990
rect 4040 4940 6090 4950
rect -1470 4920 6090 4940
rect -1470 4860 -1460 4920
rect -1400 4860 -1220 4920
rect -1160 4860 -980 4920
rect -920 4860 -740 4920
rect -680 4860 -500 4920
rect -440 4860 -260 4920
rect -200 4860 -20 4920
rect 40 4860 220 4920
rect 280 4860 460 4920
rect 520 4860 700 4920
rect 760 4860 940 4920
rect 1000 4860 1580 4920
rect 1640 4860 1820 4920
rect 1880 4860 2060 4920
rect 2120 4860 2300 4920
rect 2360 4860 2540 4920
rect 2600 4860 2780 4920
rect 2840 4860 3020 4920
rect 3080 4860 3260 4920
rect 3320 4860 3500 4920
rect 3560 4860 3740 4920
rect 3800 4860 3980 4920
rect 4040 4890 6090 4920
rect 6150 4890 6190 4950
rect 6250 4890 6290 4950
rect 7040 4980 7120 4990
rect 7040 4920 7050 4980
rect 7110 4970 7120 4980
rect 8730 4970 8740 4980
rect 7110 4930 8740 4970
rect 7110 4920 7120 4930
rect 7040 4910 7120 4920
rect 4040 4860 6290 4890
rect -1470 4850 6290 4860
rect 7630 4890 7710 4930
rect 8730 4920 8740 4930
rect 8800 4920 8810 4980
rect 9140 4910 9220 4920
rect 7630 4830 7640 4890
rect 7700 4830 7710 4890
rect 7630 4820 7710 4830
rect 8070 4890 8150 4900
rect 8070 4830 8080 4890
rect 8140 4830 8150 4890
rect 9140 4850 9150 4910
rect 9210 4900 9220 4910
rect 9210 4890 9990 4900
rect 9210 4860 9920 4890
rect 9210 4850 9220 4860
rect 9140 4840 9220 4850
rect 8070 4820 8150 4830
rect 9910 4830 9920 4860
rect 9980 4830 9990 4890
rect 9910 4820 9990 4830
rect 10750 4890 11310 4900
rect 10750 4830 10760 4890
rect 10820 4830 11240 4890
rect 11300 4830 11310 4890
rect 10750 4820 11310 4830
rect 11450 4820 11560 4840
rect -3540 4810 1150 4820
rect -3540 4750 -3530 4810
rect -3470 4750 -1340 4810
rect -1280 4750 -620 4810
rect -560 4750 100 4810
rect 160 4750 820 4810
rect 880 4750 1080 4810
rect 1140 4750 1150 4810
rect -3540 4740 1150 4750
rect 1430 4810 5660 4820
rect 1430 4750 1440 4810
rect 1500 4750 1700 4810
rect 1760 4750 2420 4810
rect 2480 4750 3140 4810
rect 3200 4750 3860 4810
rect 3920 4750 5590 4810
rect 5650 4750 5660 4810
rect 1430 4740 5660 4750
rect 11450 4750 11470 4820
rect 11540 4750 11560 4820
rect -620 4710 -560 4740
rect 3140 4700 3200 4740
rect 11450 4730 11560 4750
rect 7930 4510 8010 4520
rect -1110 4470 -1030 4480
rect -1110 4410 -1100 4470
rect -1040 4460 -1030 4470
rect -390 4470 -310 4480
rect -390 4460 -380 4470
rect -1040 4420 -380 4460
rect -1040 4410 -1030 4420
rect -1110 4400 -1030 4410
rect -390 4410 -380 4420
rect -320 4460 -310 4470
rect 330 4470 410 4480
rect 330 4460 340 4470
rect -320 4420 340 4460
rect -320 4410 -310 4420
rect -390 4400 -310 4410
rect 330 4410 340 4420
rect 400 4410 410 4470
rect 330 4400 410 4410
rect 2170 4470 2250 4480
rect 2170 4410 2180 4470
rect 2240 4460 2250 4470
rect 2890 4470 2970 4480
rect 2890 4460 2900 4470
rect 2240 4420 2900 4460
rect 2240 4410 2250 4420
rect 2170 4400 2250 4410
rect 2890 4410 2900 4420
rect 2960 4460 2970 4470
rect 3610 4470 3690 4480
rect 3610 4460 3620 4470
rect 2960 4420 3620 4460
rect 2960 4410 2970 4420
rect 2890 4400 2970 4410
rect 3610 4410 3620 4420
rect 3680 4410 3690 4470
rect 7930 4450 7940 4510
rect 8000 4450 8010 4510
rect 7930 4440 8010 4450
rect 3610 4400 3690 4410
rect 6050 4410 6290 4420
rect 6050 4400 10210 4410
rect -1370 4350 830 4360
rect -1370 4290 -1360 4350
rect -1300 4290 -1280 4350
rect -1220 4290 -860 4350
rect -800 4290 -620 4350
rect -560 4290 -140 4350
rect -80 4290 100 4350
rect 160 4290 580 4350
rect 640 4290 760 4350
rect 820 4290 830 4350
rect -1370 4280 830 4290
rect 1750 4350 4600 4360
rect 1750 4290 1760 4350
rect 1820 4290 1940 4350
rect 2000 4290 2180 4350
rect 2240 4290 2420 4350
rect 2480 4290 2660 4350
rect 2720 4290 3140 4350
rect 3200 4290 3380 4350
rect 3440 4290 3800 4350
rect 3860 4290 4370 4350
rect 4430 4290 4450 4350
rect 4510 4290 4530 4350
rect 4590 4290 4600 4350
rect 6050 4340 6090 4400
rect 6150 4340 6190 4400
rect 6250 4340 7540 4400
rect 7600 4340 7740 4400
rect 7800 4340 8140 4400
rect 8200 4340 8540 4400
rect 8600 4340 8940 4400
rect 9000 4340 9020 4400
rect 9080 4340 9340 4400
rect 9400 4340 9540 4400
rect 9600 4340 10140 4400
rect 10200 4340 10210 4400
rect 6050 4330 10210 4340
rect 6050 4320 6290 4330
rect 1750 4270 4600 4290
rect 1750 4210 1760 4270
rect 1820 4210 1940 4270
rect 2000 4210 2180 4270
rect 2240 4210 2420 4270
rect 2480 4210 2660 4270
rect 2720 4210 3140 4270
rect 3200 4210 3380 4270
rect 3440 4210 3800 4270
rect 3860 4210 4370 4270
rect 4430 4210 4450 4270
rect 4510 4210 4530 4270
rect 4590 4210 4600 4270
rect 1750 4190 4600 4210
rect 7930 4260 9210 4270
rect 7930 4200 7940 4260
rect 8000 4200 9140 4260
rect 9200 4200 9210 4260
rect 7930 4190 9210 4200
rect 1750 4130 1760 4190
rect 1820 4130 1940 4190
rect 2000 4130 2180 4190
rect 2240 4130 2420 4190
rect 2480 4130 2660 4190
rect 2720 4130 3140 4190
rect 3200 4130 3380 4190
rect 3440 4130 3800 4190
rect 3860 4130 4370 4190
rect 4430 4130 4450 4190
rect 4510 4130 4530 4190
rect 4590 4130 4600 4190
rect 1750 4120 4600 4130
rect -630 4080 410 4090
rect -630 4020 -620 4080
rect -560 4020 -140 4080
rect -80 4020 340 4080
rect 400 4020 410 4080
rect -630 4010 410 4020
rect 2170 4080 3210 4090
rect 2170 4020 2180 4080
rect 2240 4020 2660 4080
rect 2720 4020 3140 4080
rect 3200 4020 3210 4080
rect 2170 4010 3210 4020
rect -390 3970 650 3980
rect -390 3910 -380 3970
rect -320 3910 100 3970
rect 160 3910 580 3970
rect 640 3910 650 3970
rect -390 3900 650 3910
rect 1930 3970 2970 3980
rect 1930 3910 1940 3970
rect 2000 3910 2420 3970
rect 2480 3910 2900 3970
rect 2960 3910 2970 3970
rect 1930 3900 2970 3910
rect -2420 3870 -2340 3880
rect 4250 3870 4330 3880
rect -2420 3810 -2410 3870
rect -2350 3860 560 3870
rect -2350 3810 -454 3860
rect -2420 3808 -454 3810
rect -402 3808 -296 3860
rect -244 3808 28 3860
rect 80 3808 182 3860
rect 234 3808 506 3860
rect 558 3808 560 3860
rect 2020 3860 4260 3870
rect -2420 3800 560 3808
rect 810 3820 1770 3830
rect 810 3760 820 3820
rect 880 3760 1180 3820
rect 1240 3760 1260 3820
rect 1320 3760 1340 3820
rect 1400 3760 1700 3820
rect 1760 3760 1770 3820
rect 2020 3808 2022 3860
rect 2074 3808 2346 3860
rect 2398 3808 2500 3860
rect 2552 3808 2824 3860
rect 2876 3808 2982 3860
rect 3034 3810 4260 3860
rect 4320 3810 4330 3870
rect 3034 3808 4330 3810
rect 2020 3800 4330 3808
rect 810 3740 1770 3760
rect 810 3680 820 3740
rect 880 3680 1180 3740
rect 1240 3680 1260 3740
rect 1320 3680 1340 3740
rect 1400 3680 1700 3740
rect 1760 3680 1770 3740
rect 810 3660 1770 3680
rect -2310 3640 -2230 3650
rect -2310 3580 -2300 3640
rect -2240 3632 459 3640
rect -2240 3580 -557 3632
rect -505 3580 -197 3632
rect -145 3580 -77 3632
rect -25 3580 283 3632
rect 335 3580 403 3632
rect 455 3580 459 3632
rect 810 3600 820 3660
rect 880 3600 1180 3660
rect 1240 3600 1260 3660
rect 1320 3600 1340 3660
rect 1400 3600 1700 3660
rect 1760 3600 1770 3660
rect 4160 3640 4240 3650
rect 810 3590 1770 3600
rect 2121 3632 4170 3640
rect -2310 3570 459 3580
rect 2121 3580 2125 3632
rect 2177 3580 2245 3632
rect 2297 3580 2605 3632
rect 2657 3580 2725 3632
rect 2777 3580 3085 3632
rect 3137 3580 4170 3632
rect 4230 3580 4240 3640
rect 2121 3570 4240 3580
rect 7150 3600 8810 3610
rect 7150 3540 7160 3600
rect 7220 3540 8340 3600
rect 8400 3540 8740 3600
rect 8800 3540 8810 3600
rect -1250 3530 540 3540
rect -1250 3470 -1240 3530
rect -1180 3470 -490 3530
rect -430 3470 -270 3530
rect -210 3470 -10 3530
rect 50 3470 210 3530
rect 270 3470 470 3530
rect 530 3470 540 3530
rect -1250 3460 540 3470
rect 2040 3530 3830 3540
rect 7150 3530 8810 3540
rect 2040 3470 2050 3530
rect 2110 3470 2310 3530
rect 2370 3470 2530 3530
rect 2590 3470 2790 3530
rect 2850 3470 3010 3530
rect 3070 3470 3760 3530
rect 3820 3470 3830 3530
rect 2040 3460 3830 3470
rect -1070 3420 6290 3430
rect -1070 3360 -1060 3420
rect -1000 3360 -820 3420
rect -760 3360 -580 3420
rect -520 3360 -340 3420
rect -280 3360 300 3420
rect 360 3360 540 3420
rect 600 3360 780 3420
rect 840 3360 1740 3420
rect 1800 3360 1980 3420
rect 2040 3360 2220 3420
rect 2280 3360 2860 3420
rect 2920 3360 3100 3420
rect 3160 3360 3340 3420
rect 3400 3360 3580 3420
rect 3640 3390 6290 3420
rect 3640 3360 6090 3390
rect -1070 3340 6090 3360
rect -1070 3280 -1060 3340
rect -1000 3280 -820 3340
rect -760 3280 -580 3340
rect -520 3280 -340 3340
rect -280 3280 300 3340
rect 360 3280 540 3340
rect 600 3280 780 3340
rect 840 3280 1740 3340
rect 1800 3280 1980 3340
rect 2040 3280 2220 3340
rect 2280 3280 2860 3340
rect 2920 3280 3100 3340
rect 3160 3280 3340 3340
rect 3400 3280 3580 3340
rect 3640 3330 6090 3340
rect 6150 3330 6190 3390
rect 6250 3330 6290 3390
rect 3640 3290 6290 3330
rect 3640 3280 6090 3290
rect -1070 3260 6090 3280
rect -1070 3200 -1060 3260
rect -1000 3200 -820 3260
rect -760 3200 -580 3260
rect -520 3200 -340 3260
rect -280 3200 300 3260
rect 360 3200 540 3260
rect 600 3200 780 3260
rect 840 3200 1740 3260
rect 1800 3200 1980 3260
rect 2040 3200 2220 3260
rect 2280 3200 2860 3260
rect 2920 3200 3100 3260
rect 3160 3200 3340 3260
rect 3400 3200 3580 3260
rect 3640 3230 6090 3260
rect 6150 3230 6190 3290
rect 6250 3230 6290 3290
rect 3640 3200 6290 3230
rect -1070 3190 6290 3200
rect 6350 3210 11100 3220
rect 6350 3150 6390 3210
rect 6450 3150 6490 3210
rect 6550 3150 11030 3210
rect 11090 3150 11100 3210
rect 6350 3140 11100 3150
rect 6050 2970 6290 2990
rect 6050 2910 6090 2970
rect 6150 2910 6190 2970
rect 6250 2910 6290 2970
rect 6050 2890 6290 2910
rect 11220 2880 11320 2900
rect 11220 2820 11240 2880
rect 11300 2820 11320 2880
rect 11220 2800 11320 2820
rect -90 2620 6590 2630
rect -90 2560 -80 2620
rect -20 2560 1180 2620
rect 1240 2560 1260 2620
rect 1320 2560 1340 2620
rect 1400 2560 2600 2620
rect 2660 2590 6590 2620
rect 2660 2560 6390 2590
rect -90 2540 6390 2560
rect -90 2480 -80 2540
rect -20 2480 1180 2540
rect 1240 2480 1260 2540
rect 1320 2480 1340 2540
rect 1400 2480 2600 2540
rect 2660 2530 6390 2540
rect 6450 2530 6490 2590
rect 6550 2530 6590 2590
rect 2660 2490 6590 2530
rect 2660 2480 6390 2490
rect -90 2460 6390 2480
rect -90 2400 -80 2460
rect -20 2400 1180 2460
rect 1240 2400 1260 2460
rect 1320 2400 1340 2460
rect 1400 2400 2600 2460
rect 2660 2430 6390 2460
rect 6450 2430 6490 2490
rect 6550 2430 6590 2490
rect 2660 2400 6590 2430
rect -90 2390 6590 2400
rect -830 2350 -750 2360
rect -830 2290 -820 2350
rect -760 2340 -750 2350
rect -670 2350 -590 2360
rect -670 2340 -660 2350
rect -760 2300 -660 2340
rect -760 2290 -750 2300
rect -830 2280 -750 2290
rect -670 2290 -660 2300
rect -600 2340 -590 2350
rect -510 2350 -430 2360
rect -510 2340 -500 2350
rect -600 2300 -500 2340
rect -600 2290 -590 2300
rect -670 2280 -590 2290
rect -510 2290 -500 2300
rect -440 2340 -430 2350
rect -350 2350 -270 2360
rect -350 2340 -340 2350
rect -440 2300 -340 2340
rect -440 2290 -430 2300
rect -510 2280 -430 2290
rect -350 2290 -340 2300
rect -280 2340 -270 2350
rect -190 2350 -110 2360
rect -190 2340 -180 2350
rect -280 2300 -180 2340
rect -280 2290 -270 2300
rect -350 2280 -270 2290
rect -190 2290 -180 2300
rect -120 2340 -110 2350
rect -30 2350 50 2360
rect -30 2340 -20 2350
rect -120 2300 -20 2340
rect -120 2290 -110 2300
rect -190 2280 -110 2290
rect -30 2290 -20 2300
rect 40 2340 50 2350
rect 130 2350 210 2360
rect 130 2340 140 2350
rect 40 2300 140 2340
rect 40 2290 50 2300
rect -30 2280 50 2290
rect 130 2290 140 2300
rect 200 2340 210 2350
rect 290 2350 370 2360
rect 290 2340 300 2350
rect 200 2300 300 2340
rect 200 2290 210 2300
rect 130 2280 210 2290
rect 290 2290 300 2300
rect 360 2340 370 2350
rect 450 2350 530 2360
rect 450 2340 460 2350
rect 360 2300 460 2340
rect 360 2290 370 2300
rect 290 2280 370 2290
rect 450 2290 460 2300
rect 520 2340 530 2350
rect 610 2350 690 2360
rect 610 2340 620 2350
rect 520 2300 620 2340
rect 520 2290 530 2300
rect 450 2280 530 2290
rect 610 2290 620 2300
rect 680 2340 690 2350
rect 770 2350 850 2360
rect 770 2340 780 2350
rect 680 2300 780 2340
rect 680 2290 690 2300
rect 610 2280 690 2290
rect 770 2290 780 2300
rect 840 2340 850 2350
rect 930 2350 1010 2360
rect 930 2340 940 2350
rect 840 2300 940 2340
rect 840 2290 850 2300
rect 770 2280 850 2290
rect 930 2290 940 2300
rect 1000 2340 1010 2350
rect 1090 2350 1170 2360
rect 1090 2340 1100 2350
rect 1000 2300 1100 2340
rect 1000 2290 1010 2300
rect 930 2280 1010 2290
rect 1090 2290 1100 2300
rect 1160 2290 1170 2350
rect 1090 2280 1170 2290
rect 1250 2350 1330 2360
rect 1250 2290 1260 2350
rect 1320 2340 1330 2350
rect 1410 2350 1490 2360
rect 1410 2340 1420 2350
rect 1320 2300 1420 2340
rect 1320 2290 1330 2300
rect 1250 2280 1330 2290
rect 1410 2290 1420 2300
rect 1480 2340 1490 2350
rect 1570 2350 1650 2360
rect 1570 2340 1580 2350
rect 1480 2300 1580 2340
rect 1480 2290 1490 2300
rect 1410 2280 1490 2290
rect 1570 2290 1580 2300
rect 1640 2340 1650 2350
rect 1730 2350 1810 2360
rect 1730 2340 1740 2350
rect 1640 2300 1740 2340
rect 1640 2290 1650 2300
rect 1570 2280 1650 2290
rect 1730 2290 1740 2300
rect 1800 2340 1810 2350
rect 1890 2350 1970 2360
rect 1890 2340 1900 2350
rect 1800 2300 1900 2340
rect 1800 2290 1810 2300
rect 1730 2280 1810 2290
rect 1890 2290 1900 2300
rect 1960 2340 1970 2350
rect 2050 2350 2130 2360
rect 2050 2340 2060 2350
rect 1960 2300 2060 2340
rect 1960 2290 1970 2300
rect 1890 2280 1970 2290
rect 2050 2290 2060 2300
rect 2120 2340 2130 2350
rect 2210 2350 2290 2360
rect 2210 2340 2220 2350
rect 2120 2300 2220 2340
rect 2120 2290 2130 2300
rect 2050 2280 2130 2290
rect 2210 2290 2220 2300
rect 2280 2340 2290 2350
rect 2370 2350 2450 2360
rect 2370 2340 2380 2350
rect 2280 2300 2380 2340
rect 2280 2290 2290 2300
rect 2210 2280 2290 2290
rect 2370 2290 2380 2300
rect 2440 2340 2450 2350
rect 2530 2350 2610 2360
rect 2530 2340 2540 2350
rect 2440 2300 2540 2340
rect 2440 2290 2450 2300
rect 2370 2280 2450 2290
rect 2530 2290 2540 2300
rect 2600 2340 2610 2350
rect 2690 2350 2770 2360
rect 2690 2340 2700 2350
rect 2600 2300 2700 2340
rect 2600 2290 2610 2300
rect 2530 2280 2610 2290
rect 2690 2290 2700 2300
rect 2760 2340 2770 2350
rect 2850 2350 2930 2360
rect 2850 2340 2860 2350
rect 2760 2300 2860 2340
rect 2760 2290 2770 2300
rect 2690 2280 2770 2290
rect 2850 2290 2860 2300
rect 2920 2340 2930 2350
rect 3010 2350 3090 2360
rect 3010 2340 3020 2350
rect 2920 2300 3020 2340
rect 2920 2290 2930 2300
rect 2850 2280 2930 2290
rect 3010 2290 3020 2300
rect 3080 2340 3090 2350
rect 3170 2350 3250 2360
rect 3170 2340 3180 2350
rect 3080 2300 3180 2340
rect 3080 2290 3090 2300
rect 3010 2280 3090 2290
rect 3170 2290 3180 2300
rect 3240 2290 3250 2350
rect 3170 2280 3250 2290
rect 3480 2220 6590 2230
rect -2530 2180 -830 2190
rect -2530 2120 -2520 2180
rect -2460 2120 -900 2180
rect -840 2120 -830 2180
rect -2530 2110 -830 2120
rect 3480 2160 3490 2220
rect 3550 2180 6590 2220
rect 3550 2160 6390 2180
rect 3480 2140 6390 2160
rect 3480 2080 3490 2140
rect 3550 2120 6390 2140
rect 6450 2120 6490 2180
rect 6550 2120 6590 2180
rect 3550 2080 6590 2120
rect 3480 2070 6590 2080
rect -1370 2010 6740 2020
rect -1370 1950 -1360 2010
rect -1300 1950 -950 2010
rect -890 1950 6670 2010
rect 6730 1950 6740 2010
rect -1370 1940 6740 1950
rect -2310 1900 4870 1910
rect -2310 1840 -2300 1900
rect -2240 1840 4800 1900
rect 4860 1840 4870 1900
rect -2310 1830 4870 1840
rect 4160 1790 4240 1800
rect -850 1780 562 1790
rect -850 1720 -840 1780
rect -780 1720 562 1780
rect 632 1720 642 1790
rect 1950 1720 1960 1790
rect 2030 1780 2040 1790
rect 4160 1780 4170 1790
rect 2030 1740 4170 1780
rect 2030 1720 2040 1740
rect 4160 1730 4170 1740
rect 4230 1730 4240 1790
rect 4160 1720 4240 1730
rect -850 1710 560 1720
rect -1640 1670 2040 1680
rect -1640 1610 -1630 1670
rect -1570 1610 1970 1670
rect 2030 1610 2040 1670
rect -1640 1600 2040 1610
rect 3350 1590 4330 1600
rect 3350 1530 3360 1590
rect 3420 1530 4020 1590
rect 4080 1530 4260 1590
rect 4320 1530 4330 1590
rect 3350 1520 4330 1530
rect 4360 1040 6890 1060
rect 4360 980 4370 1040
rect 4430 980 4450 1040
rect 4510 980 4530 1040
rect 4590 980 6810 1040
rect 6870 980 6890 1040
rect 4360 960 6890 980
rect 5960 340 7080 350
rect 5960 280 5970 340
rect 6030 280 7010 340
rect 7070 280 7080 340
rect 5960 270 7080 280
rect 5580 -360 6890 -340
rect -850 -420 -340 -410
rect -850 -480 -840 -420
rect -780 -480 -410 -420
rect -350 -480 -340 -420
rect -850 -490 -340 -480
rect 1250 -420 3430 -410
rect 1250 -480 1260 -420
rect 1320 -480 3360 -420
rect 3420 -480 3430 -420
rect 5580 -420 5590 -360
rect 5650 -420 6810 -360
rect 6870 -420 6890 -360
rect 5580 -440 6890 -420
rect 1250 -490 3430 -480
rect 6130 -1060 6210 -1050
rect 6130 -1120 6140 -1060
rect 6200 -1120 6210 -1060
rect 6130 -1130 6210 -1120
rect -3540 -1710 -3040 -1700
rect -3540 -2110 -3530 -1710
rect -3470 -1720 -3040 -1710
rect -3470 -1780 -3110 -1720
rect -3050 -1780 -3040 -1720
rect -3470 -1800 -3040 -1780
rect -3470 -1860 -3110 -1800
rect -3050 -1860 -3040 -1800
rect -3470 -1890 -3040 -1860
rect -3470 -1950 -3110 -1890
rect -3050 -1950 -3040 -1890
rect -3470 -1980 -3040 -1950
rect -3470 -2040 -3110 -1980
rect -3050 -2040 -3040 -1980
rect -3470 -2060 -3040 -2040
rect -3470 -2110 -3110 -2060
rect -3540 -2120 -3110 -2110
rect -3050 -2120 -3040 -2060
rect -3540 -2130 -3040 -2120
rect 5580 -1710 6040 -1700
rect 5580 -2110 5590 -1710
rect 5650 -1720 6040 -1710
rect 5650 -1780 5970 -1720
rect 6030 -1780 6040 -1720
rect 5650 -1800 6040 -1780
rect 5650 -1860 5970 -1800
rect 6030 -1860 6040 -1800
rect 6650 -1760 6750 -1740
rect 6650 -1820 6670 -1760
rect 6730 -1820 6750 -1760
rect 6650 -1840 6750 -1820
rect 5650 -1890 6040 -1860
rect 5650 -1950 5970 -1890
rect 6030 -1950 6040 -1890
rect 5650 -1980 6040 -1950
rect 5650 -2040 5970 -1980
rect 6030 -2040 6040 -1980
rect 5650 -2060 6040 -2040
rect 5650 -2110 5970 -2060
rect 5580 -2120 5970 -2110
rect 6030 -2120 6040 -2060
rect 5580 -2130 6040 -2120
rect 6200 -2460 6280 -2450
rect 6200 -2520 6210 -2460
rect 6270 -2520 6280 -2460
rect -3540 -2530 5660 -2520
rect 6200 -2530 6280 -2520
rect -3540 -2590 -3530 -2530
rect -3470 -2590 -2740 -2530
rect -2680 -2590 -1300 -2530
rect -1240 -2590 1260 -2530
rect 1320 -2590 3690 -2530
rect 3750 -2590 4800 -2530
rect 4860 -2590 5590 -2530
rect 5650 -2590 5660 -2530
rect -3540 -2610 5660 -2590
rect -3540 -2670 -3530 -2610
rect -3470 -2670 -2740 -2610
rect -2680 -2670 -1300 -2610
rect -1240 -2670 1260 -2610
rect 1320 -2670 3690 -2610
rect 3750 -2670 4800 -2610
rect 4860 -2670 5590 -2610
rect 5650 -2670 5660 -2610
rect -3540 -2690 5660 -2670
rect -3540 -2750 -3530 -2690
rect -3470 -2750 -2740 -2690
rect -2680 -2750 -1300 -2690
rect -1240 -2750 1260 -2690
rect 1320 -2750 3690 -2690
rect 3750 -2750 4800 -2690
rect 4860 -2750 5590 -2690
rect 5650 -2750 5660 -2690
rect -3540 -2760 5660 -2750
rect -3120 -2800 6280 -2790
rect -3120 -2860 -3110 -2800
rect -3050 -2860 6210 -2800
rect 6270 -2860 6280 -2800
rect -3120 -2870 6280 -2860
rect -3070 -3100 -2970 -3090
rect 14000 -3100 14100 -3090
rect -3070 -3110 3430 -3100
rect -3070 -3170 -3050 -3110
rect -2990 -3170 3010 -3110
rect 3420 -3170 3430 -3110
rect -3070 -3180 3430 -3170
rect 4910 -3110 14100 -3100
rect 4910 -3170 4920 -3110
rect 5330 -3170 14020 -3110
rect 14080 -3170 14100 -3110
rect 4910 -3180 14100 -3170
rect -3070 -3190 -2970 -3180
rect 14000 -3190 14100 -3180
rect 4130 -3300 4210 -3290
rect 4130 -3360 4140 -3300
rect 4200 -3360 4210 -3300
rect 4130 -3370 4210 -3360
rect -4270 -3390 11420 -3370
rect -4270 -3460 10830 -3390
rect 10900 -3460 11330 -3390
rect 11400 -3460 11420 -3390
rect -4270 -3480 11420 -3460
<< via2 >>
rect 10620 14820 10680 14880
rect 10620 14720 10680 14780
rect 250 13420 310 13480
rect 250 13320 310 13380
rect 250 12640 310 12700
rect 250 12540 310 12600
rect 10620 10740 10680 10800
rect 10620 10640 10680 10700
rect 940 10440 1000 10500
rect 940 10340 1000 10400
rect 11010 10450 11080 10520
rect 7290 9940 7350 10000
rect 7390 9940 7450 10000
rect 940 9260 1000 9320
rect 940 9160 1000 9220
rect 10770 9270 10840 9340
rect 10770 8740 10840 8810
rect 940 8080 1000 8140
rect 6390 8100 6450 8160
rect 6490 8100 6550 8160
rect 940 7980 1000 8040
rect 11120 7950 11190 8020
rect 11240 7200 11300 7260
rect 6090 6910 6150 6970
rect 6190 6910 6250 6970
rect 6390 6680 6450 6740
rect 6490 6680 6550 6740
rect 6090 6440 6150 6500
rect 6190 6440 6250 6500
rect 6090 6340 6150 6400
rect 6190 6340 6250 6400
rect 6390 5560 6450 5620
rect 6490 5560 6550 5620
rect 11470 5260 11540 5330
rect 6090 4990 6150 5050
rect 6190 4990 6250 5050
rect 6090 4890 6150 4950
rect 6190 4890 6250 4950
rect 11470 4750 11540 4820
rect 6090 4340 6150 4400
rect 6190 4340 6250 4400
rect 6090 3330 6150 3390
rect 6190 3330 6250 3390
rect 6090 3230 6150 3290
rect 6190 3230 6250 3290
rect 6390 3150 6450 3210
rect 6490 3150 6550 3210
rect 6090 2910 6150 2970
rect 6190 2910 6250 2970
rect 11240 2820 11300 2880
rect 6390 2530 6450 2590
rect 6490 2530 6550 2590
rect 6390 2430 6450 2490
rect 6490 2430 6550 2490
rect 6390 2120 6450 2180
rect 6490 2120 6550 2180
rect 6810 980 6870 1040
rect 7010 280 7070 340
rect 6810 -420 6870 -360
rect 6140 -1120 6200 -1060
rect 6670 -1820 6730 -1760
rect 6210 -2520 6270 -2460
rect -3050 -3170 -2990 -3110
rect 14020 -3170 14080 -3110
rect 10830 -3460 10900 -3390
rect 11330 -3460 11400 -3390
<< metal3 >>
rect -4270 14880 10700 14920
rect -4270 14820 10620 14880
rect 10680 14820 10700 14880
rect -4270 14780 10700 14820
rect -4270 14720 10620 14780
rect 10680 14720 10700 14780
rect -4270 14680 10700 14720
rect -4270 13480 330 13520
rect -4270 13420 250 13480
rect 310 13420 330 13480
rect -4270 13380 330 13420
rect -4270 13320 250 13380
rect 310 13320 330 13380
rect -4270 13280 330 13320
rect -4270 12700 330 12740
rect -4270 12640 250 12700
rect 310 12640 330 12700
rect -4270 12600 330 12640
rect -4270 12540 250 12600
rect 310 12540 330 12600
rect -4270 12500 330 12540
rect -4270 10800 10700 10840
rect -4270 10740 10620 10800
rect 10680 10740 10700 10800
rect -4270 10700 10700 10740
rect -4270 10640 10620 10700
rect 10680 10640 10700 10700
rect -4270 10600 10700 10640
rect -4270 10500 1020 10540
rect -4270 10440 940 10500
rect 1000 10440 1020 10500
rect -4270 10400 1020 10440
rect -4270 10340 940 10400
rect 1000 10340 1020 10400
rect -4270 10300 1020 10340
rect 7250 10000 7490 10600
rect 10990 10520 12200 10540
rect 10990 10450 11010 10520
rect 11080 10450 12200 10520
rect 10990 10430 12200 10450
rect 7250 9940 7290 10000
rect 7350 9940 7390 10000
rect 7450 9940 7490 10000
rect 7250 9930 7490 9940
rect -4270 9320 1020 9360
rect -4270 9260 940 9320
rect 1000 9260 1020 9320
rect -4270 9220 1020 9260
rect 10750 9340 10860 9360
rect 10750 9270 10770 9340
rect 10840 9270 10860 9340
rect 10750 9250 10860 9270
rect 11100 9220 12200 10430
rect -4270 9160 940 9220
rect 1000 9160 1020 9220
rect -4270 9120 1020 9160
rect 10750 8810 10860 8830
rect 10750 8740 10770 8810
rect 10840 8740 10860 8810
rect 10750 8720 10860 8740
rect -4270 8140 1020 8180
rect -4270 8080 940 8140
rect 1000 8080 1020 8140
rect -4270 8040 1020 8080
rect -4270 7980 940 8040
rect 1000 7980 1020 8040
rect -4270 7940 1020 7980
rect 6350 8160 6590 8170
rect 6350 8100 6390 8160
rect 6450 8100 6490 8160
rect 6550 8100 6590 8160
rect 6350 7830 6590 8100
rect 11100 8040 11700 8860
rect 11100 8020 11210 8040
rect 11100 7950 11120 8020
rect 11190 7950 11210 8020
rect 11100 7930 11210 7950
rect -4270 7590 6590 7830
rect -4270 7290 6290 7530
rect 6050 6970 6290 7290
rect 6050 6910 6090 6970
rect 6150 6910 6190 6970
rect 6250 6910 6290 6970
rect 6050 6500 6290 6910
rect 6050 6440 6090 6500
rect 6150 6440 6190 6500
rect 6250 6440 6290 6500
rect 6050 6400 6290 6440
rect 6050 6340 6090 6400
rect 6150 6340 6190 6400
rect 6250 6340 6290 6400
rect 6050 5050 6290 6340
rect 6050 4990 6090 5050
rect 6150 4990 6190 5050
rect 6250 4990 6290 5050
rect 6050 4950 6290 4990
rect 6050 4890 6090 4950
rect 6150 4890 6190 4950
rect 6250 4890 6290 4950
rect 6050 4400 6290 4890
rect 6050 4340 6090 4400
rect 6150 4340 6190 4400
rect 6250 4340 6290 4400
rect 6050 3390 6290 4340
rect 6050 3330 6090 3390
rect 6150 3330 6190 3390
rect 6250 3330 6290 3390
rect 6050 3290 6290 3330
rect 6050 3230 6090 3290
rect 6150 3230 6190 3290
rect 6250 3230 6290 3290
rect 6050 2970 6290 3230
rect 6050 2910 6090 2970
rect 6150 2910 6190 2970
rect 6250 2910 6290 2970
rect 6050 2890 6290 2910
rect 6350 6740 6590 7590
rect 11220 7270 11320 7280
rect 11220 7260 13860 7270
rect 11220 7200 11240 7260
rect 11300 7200 13860 7260
rect 11220 7180 13860 7200
rect 6350 6680 6390 6740
rect 6450 6680 6490 6740
rect 6550 6680 6590 6740
rect 6350 5620 6590 6680
rect 6350 5560 6390 5620
rect 6450 5560 6490 5620
rect 6550 5560 6590 5620
rect 6350 3210 6590 5560
rect 11450 5330 11560 5350
rect 11450 5260 11470 5330
rect 11540 5260 11560 5330
rect 11450 5240 11560 5260
rect 11800 5210 13860 7180
rect 11450 4820 11560 4840
rect 11450 4750 11470 4820
rect 11540 4750 11560 4820
rect 11450 4730 11560 4750
rect 6350 3150 6390 3210
rect 6450 3150 6490 3210
rect 6550 3150 6590 3210
rect 6350 2590 6590 3150
rect 11800 2900 13860 4870
rect 11220 2880 13860 2900
rect 11220 2820 11240 2880
rect 11300 2820 13860 2880
rect 11220 2810 13860 2820
rect 11220 2800 11320 2810
rect 6350 2530 6390 2590
rect 6450 2530 6490 2590
rect 6550 2530 6590 2590
rect 6350 2490 6590 2530
rect 6350 2430 6390 2490
rect 6450 2430 6490 2490
rect 6550 2430 6590 2490
rect 6350 2180 6590 2430
rect 6350 2120 6390 2180
rect 6450 2120 6490 2180
rect 6550 2120 6590 2180
rect 6350 2070 6590 2120
rect 7130 1060 7590 1250
rect 7830 1060 8290 1250
rect 8530 1060 8990 1250
rect 9230 1060 9690 1250
rect 9930 1060 10390 1250
rect 10630 1060 11090 1250
rect 11330 1060 11790 1250
rect 12030 1060 12490 1250
rect 12730 1060 13190 1250
rect 13430 1060 13890 1250
rect 6790 1050 6890 1060
rect 6790 970 6800 1050
rect 6880 970 6890 1050
rect 6790 960 6890 970
rect 7130 960 13890 1060
rect 7130 790 7590 960
rect 7830 790 8290 960
rect 8530 790 8990 960
rect 9230 790 9690 960
rect 9930 790 10390 960
rect 10630 790 11090 960
rect 11330 790 11790 960
rect 12030 790 12490 960
rect 12730 790 13190 960
rect 13430 790 13890 960
rect 13610 550 13710 790
rect 7130 360 7590 550
rect 7830 360 8290 550
rect 8530 360 8990 550
rect 9230 360 9690 550
rect 9930 360 10390 550
rect 10630 360 11090 550
rect 11330 360 11790 550
rect 12030 360 12490 550
rect 12730 360 13190 550
rect 13430 360 13890 550
rect 7130 350 13890 360
rect 7000 340 13890 350
rect 7000 280 7010 340
rect 7070 280 13890 340
rect 7000 270 13890 280
rect 7130 260 13890 270
rect 7130 90 7590 260
rect 7830 90 8290 260
rect 8530 90 8990 260
rect 9230 90 9690 260
rect 9930 90 10390 260
rect 10630 90 11090 260
rect 11330 90 11790 260
rect 12030 90 12490 260
rect 12730 90 13190 260
rect 13430 90 13890 260
rect 7130 -340 7590 -150
rect 7830 -340 8290 -150
rect 8530 -340 8990 -150
rect 9230 -340 9690 -150
rect 9930 -340 10390 -150
rect 10630 -340 11090 -150
rect 11330 -340 11790 -150
rect 12030 -340 12490 -150
rect 12730 -340 13190 -150
rect 13430 -340 13890 -150
rect 6790 -350 6890 -340
rect 6790 -430 6800 -350
rect 6880 -430 6890 -350
rect 6790 -440 6890 -430
rect 7130 -440 13890 -340
rect 7130 -610 7590 -440
rect 7830 -610 8290 -440
rect 8530 -610 8990 -440
rect 9230 -610 9690 -440
rect 9930 -610 10390 -440
rect 10630 -610 11090 -440
rect 11330 -610 11790 -440
rect 12030 -610 12490 -440
rect 12730 -610 13190 -440
rect 13430 -610 13890 -440
rect 13610 -850 13710 -610
rect 7130 -1040 7590 -850
rect 7830 -1040 8290 -850
rect 8530 -1040 8990 -850
rect 9230 -1040 9690 -850
rect 9930 -1040 10390 -850
rect 10630 -1040 11090 -850
rect 11330 -1040 11790 -850
rect 12030 -1040 12490 -850
rect 12730 -1040 13190 -850
rect 13430 -1040 13890 -850
rect 7130 -1050 13890 -1040
rect 6130 -1060 13890 -1050
rect 6130 -1120 6140 -1060
rect 6200 -1120 13890 -1060
rect 6130 -1130 13890 -1120
rect 7130 -1140 13890 -1130
rect 7130 -1310 7590 -1140
rect 7830 -1310 8290 -1140
rect 8530 -1310 8990 -1140
rect 9230 -1310 9690 -1140
rect 9930 -1310 10390 -1140
rect 10630 -1310 11090 -1140
rect 11330 -1310 11790 -1140
rect 12030 -1310 12490 -1140
rect 12730 -1310 13190 -1140
rect 13430 -1310 13890 -1140
rect 7130 -1740 7590 -1550
rect 7830 -1740 8290 -1550
rect 8530 -1740 8990 -1550
rect 9230 -1740 9690 -1550
rect 9930 -1740 10390 -1550
rect 10630 -1740 11090 -1550
rect 11330 -1740 11790 -1550
rect 12030 -1740 12490 -1550
rect 12730 -1740 13190 -1550
rect 13430 -1740 13890 -1550
rect 6650 -1750 6750 -1740
rect 6650 -1830 6660 -1750
rect 6740 -1830 6750 -1750
rect 6650 -1840 6750 -1830
rect 7130 -1840 13890 -1740
rect 7130 -2010 7590 -1840
rect 7830 -2010 8290 -1840
rect 8530 -2010 8990 -1840
rect 9230 -2010 9690 -1840
rect 9930 -2010 10390 -1840
rect 10630 -2010 11090 -1840
rect 11330 -2010 11790 -1840
rect 12030 -2010 12490 -1840
rect 12730 -2010 13190 -1840
rect 13430 -2010 13890 -1840
rect 13610 -2250 13710 -2010
rect 7130 -2440 7590 -2250
rect 7830 -2440 8290 -2250
rect 8530 -2440 8990 -2250
rect 9230 -2440 9690 -2250
rect 9930 -2440 10390 -2250
rect 10630 -2440 11090 -2250
rect 11330 -2440 11790 -2250
rect 12030 -2440 12490 -2250
rect 12730 -2440 13190 -2250
rect 13430 -2440 13890 -2250
rect 7130 -2450 13890 -2440
rect 6200 -2460 13890 -2450
rect 6200 -2520 6210 -2460
rect 6270 -2520 13890 -2460
rect 6200 -2530 13890 -2520
rect 7130 -2540 13890 -2530
rect 7130 -2710 7590 -2540
rect 7830 -2710 8290 -2540
rect 8530 -2710 8990 -2540
rect 9230 -2710 9690 -2540
rect 9930 -2710 10390 -2540
rect 10630 -2710 11090 -2540
rect 11330 -2710 11790 -2540
rect 12030 -2710 12490 -2540
rect 12730 -2710 13190 -2540
rect 13430 -2710 13890 -2540
rect -3070 -3110 -2970 -3090
rect -3070 -3170 -3050 -3110
rect -2990 -3170 -2970 -3110
rect -3070 -3720 -2970 -3170
rect 14000 -3110 14100 -3090
rect 14000 -3170 14020 -3110
rect 14080 -3170 14100 -3110
rect 10810 -3390 10920 -3370
rect 10810 -3460 10830 -3390
rect 10900 -3460 10920 -3390
rect 10810 -3480 10920 -3460
rect 11310 -3390 11420 -3370
rect 11310 -3460 11330 -3390
rect 11400 -3460 11420 -3390
rect 11310 -3480 11420 -3460
rect 14000 -3720 14100 -3170
rect -3070 -15780 10950 -3720
rect 11280 -15780 14100 -3720
<< via3 >>
rect 10770 9270 10840 9340
rect 10770 8740 10840 8810
rect 11470 5260 11540 5330
rect 11470 4750 11540 4820
rect 6800 1040 6880 1050
rect 6800 980 6810 1040
rect 6810 980 6870 1040
rect 6870 980 6880 1040
rect 6800 970 6880 980
rect 6800 -360 6880 -350
rect 6800 -420 6810 -360
rect 6810 -420 6870 -360
rect 6870 -420 6880 -360
rect 6800 -430 6880 -420
rect 6660 -1760 6740 -1750
rect 6660 -1820 6670 -1760
rect 6670 -1820 6730 -1760
rect 6730 -1820 6740 -1760
rect 6660 -1830 6740 -1820
rect 10830 -3460 10900 -3390
rect 11330 -3460 11400 -3390
<< mimcap >>
rect 11130 9340 12170 10510
rect 11130 9270 11150 9340
rect 11220 9270 12170 9340
rect 11130 9250 12170 9270
rect 11130 8810 11670 8830
rect 11130 8740 11150 8810
rect 11220 8740 11670 8810
rect 11130 8070 11670 8740
rect 11830 5330 13830 7240
rect 11830 5260 11850 5330
rect 11920 5260 13830 5330
rect 11830 5240 13830 5260
rect 11830 4820 13830 4840
rect 11830 4750 11850 4820
rect 11920 4750 13830 4820
rect 11830 2840 13830 4750
rect 7160 1050 7560 1220
rect 7160 970 7330 1050
rect 7410 970 7560 1050
rect 7160 820 7560 970
rect 7860 1050 8260 1220
rect 7860 970 8020 1050
rect 8100 970 8260 1050
rect 7860 820 8260 970
rect 8560 1050 8960 1220
rect 8560 970 8720 1050
rect 8800 970 8960 1050
rect 8560 820 8960 970
rect 9260 1050 9660 1220
rect 9260 970 9420 1050
rect 9500 970 9660 1050
rect 9260 820 9660 970
rect 9960 1050 10360 1220
rect 9960 970 10120 1050
rect 10200 970 10360 1050
rect 9960 820 10360 970
rect 10660 1050 11060 1220
rect 10660 970 10820 1050
rect 10900 970 11060 1050
rect 10660 820 11060 970
rect 11360 1050 11760 1220
rect 11360 970 11520 1050
rect 11600 970 11760 1050
rect 11360 820 11760 970
rect 12060 1050 12460 1220
rect 12060 970 12220 1050
rect 12300 970 12460 1050
rect 12060 820 12460 970
rect 12760 1050 13160 1220
rect 12760 970 12920 1050
rect 13000 970 13160 1050
rect 12760 820 13160 970
rect 13460 1050 13860 1220
rect 13460 970 13620 1050
rect 13700 970 13860 1050
rect 13460 820 13860 970
rect 7160 350 7560 520
rect 7160 270 7330 350
rect 7410 270 7560 350
rect 7160 120 7560 270
rect 7860 350 8260 520
rect 7860 270 8020 350
rect 8100 270 8260 350
rect 7860 120 8260 270
rect 8560 350 8960 520
rect 8560 270 8720 350
rect 8800 270 8960 350
rect 8560 120 8960 270
rect 9260 350 9660 520
rect 9260 270 9420 350
rect 9500 270 9660 350
rect 9260 120 9660 270
rect 9960 350 10360 520
rect 9960 270 10120 350
rect 10200 270 10360 350
rect 9960 120 10360 270
rect 10660 350 11060 520
rect 10660 270 10820 350
rect 10900 270 11060 350
rect 10660 120 11060 270
rect 11360 350 11760 520
rect 11360 270 11520 350
rect 11600 270 11760 350
rect 11360 120 11760 270
rect 12060 350 12460 520
rect 12060 270 12220 350
rect 12300 270 12460 350
rect 12060 120 12460 270
rect 12760 350 13160 520
rect 12760 270 12920 350
rect 13000 270 13160 350
rect 12760 120 13160 270
rect 13460 350 13860 520
rect 13460 270 13620 350
rect 13700 270 13860 350
rect 13460 120 13860 270
rect 7160 -350 7560 -180
rect 7160 -430 7330 -350
rect 7410 -430 7560 -350
rect 7160 -580 7560 -430
rect 7860 -350 8260 -180
rect 7860 -430 8020 -350
rect 8100 -430 8260 -350
rect 7860 -580 8260 -430
rect 8560 -350 8960 -180
rect 8560 -430 8720 -350
rect 8800 -430 8960 -350
rect 8560 -580 8960 -430
rect 9260 -350 9660 -180
rect 9260 -430 9420 -350
rect 9500 -430 9660 -350
rect 9260 -580 9660 -430
rect 9960 -350 10360 -180
rect 9960 -430 10120 -350
rect 10200 -430 10360 -350
rect 9960 -580 10360 -430
rect 10660 -350 11060 -180
rect 10660 -430 10820 -350
rect 10900 -430 11060 -350
rect 10660 -580 11060 -430
rect 11360 -350 11760 -180
rect 11360 -430 11520 -350
rect 11600 -430 11760 -350
rect 11360 -580 11760 -430
rect 12060 -350 12460 -180
rect 12060 -430 12220 -350
rect 12300 -430 12460 -350
rect 12060 -580 12460 -430
rect 12760 -350 13160 -180
rect 12760 -430 12920 -350
rect 13000 -430 13160 -350
rect 12760 -580 13160 -430
rect 13460 -350 13860 -180
rect 13460 -430 13620 -350
rect 13700 -430 13860 -350
rect 13460 -580 13860 -430
rect 7160 -1050 7560 -880
rect 7160 -1130 7330 -1050
rect 7410 -1130 7560 -1050
rect 7160 -1280 7560 -1130
rect 7860 -1050 8260 -880
rect 7860 -1130 8020 -1050
rect 8100 -1130 8260 -1050
rect 7860 -1280 8260 -1130
rect 8560 -1050 8960 -880
rect 8560 -1130 8720 -1050
rect 8800 -1130 8960 -1050
rect 8560 -1280 8960 -1130
rect 9260 -1050 9660 -880
rect 9260 -1130 9420 -1050
rect 9500 -1130 9660 -1050
rect 9260 -1280 9660 -1130
rect 9960 -1050 10360 -880
rect 9960 -1130 10120 -1050
rect 10200 -1130 10360 -1050
rect 9960 -1280 10360 -1130
rect 10660 -1050 11060 -880
rect 10660 -1130 10820 -1050
rect 10900 -1130 11060 -1050
rect 10660 -1280 11060 -1130
rect 11360 -1050 11760 -880
rect 11360 -1130 11520 -1050
rect 11600 -1130 11760 -1050
rect 11360 -1280 11760 -1130
rect 12060 -1050 12460 -880
rect 12060 -1130 12220 -1050
rect 12300 -1130 12460 -1050
rect 12060 -1280 12460 -1130
rect 12760 -1050 13160 -880
rect 12760 -1130 12920 -1050
rect 13000 -1130 13160 -1050
rect 12760 -1280 13160 -1130
rect 13460 -1050 13860 -880
rect 13460 -1130 13620 -1050
rect 13700 -1130 13860 -1050
rect 13460 -1280 13860 -1130
rect 7160 -1750 7560 -1580
rect 7160 -1830 7330 -1750
rect 7410 -1830 7560 -1750
rect 7160 -1980 7560 -1830
rect 7860 -1750 8260 -1580
rect 7860 -1830 8020 -1750
rect 8100 -1830 8260 -1750
rect 7860 -1980 8260 -1830
rect 8560 -1750 8960 -1580
rect 8560 -1830 8720 -1750
rect 8800 -1830 8960 -1750
rect 8560 -1980 8960 -1830
rect 9260 -1750 9660 -1580
rect 9260 -1830 9420 -1750
rect 9500 -1830 9660 -1750
rect 9260 -1980 9660 -1830
rect 9960 -1750 10360 -1580
rect 9960 -1830 10120 -1750
rect 10200 -1830 10360 -1750
rect 9960 -1980 10360 -1830
rect 10660 -1750 11060 -1580
rect 10660 -1830 10820 -1750
rect 10900 -1830 11060 -1750
rect 10660 -1980 11060 -1830
rect 11360 -1750 11760 -1580
rect 11360 -1830 11520 -1750
rect 11600 -1830 11760 -1750
rect 11360 -1980 11760 -1830
rect 12060 -1750 12460 -1580
rect 12060 -1830 12220 -1750
rect 12300 -1830 12460 -1750
rect 12060 -1980 12460 -1830
rect 12760 -1750 13160 -1580
rect 12760 -1830 12920 -1750
rect 13000 -1830 13160 -1750
rect 12760 -1980 13160 -1830
rect 13460 -1750 13860 -1580
rect 13460 -1830 13620 -1750
rect 13700 -1830 13860 -1750
rect 13460 -1980 13860 -1830
rect 7160 -2450 7560 -2280
rect 7160 -2530 7330 -2450
rect 7410 -2530 7560 -2450
rect 7160 -2680 7560 -2530
rect 7860 -2450 8260 -2280
rect 7860 -2530 8020 -2450
rect 8100 -2530 8260 -2450
rect 7860 -2680 8260 -2530
rect 8560 -2450 8960 -2280
rect 8560 -2530 8720 -2450
rect 8800 -2530 8960 -2450
rect 8560 -2680 8960 -2530
rect 9260 -2450 9660 -2280
rect 9260 -2530 9420 -2450
rect 9500 -2530 9660 -2450
rect 9260 -2680 9660 -2530
rect 9960 -2450 10360 -2280
rect 9960 -2530 10120 -2450
rect 10200 -2530 10360 -2450
rect 9960 -2680 10360 -2530
rect 10660 -2450 11060 -2280
rect 10660 -2530 10820 -2450
rect 10900 -2530 11060 -2450
rect 10660 -2680 11060 -2530
rect 11360 -2450 11760 -2280
rect 11360 -2530 11520 -2450
rect 11600 -2530 11760 -2450
rect 11360 -2680 11760 -2530
rect 12060 -2450 12460 -2280
rect 12060 -2530 12220 -2450
rect 12300 -2530 12460 -2450
rect 12060 -2680 12460 -2530
rect 12760 -2450 13160 -2280
rect 12760 -2530 12920 -2450
rect 13000 -2530 13160 -2450
rect 12760 -2680 13160 -2530
rect 13460 -2450 13860 -2280
rect 13460 -2530 13620 -2450
rect 13700 -2530 13860 -2450
rect 13460 -2680 13860 -2530
rect -3040 -3770 10920 -3750
rect -3040 -3840 10830 -3770
rect 10900 -3840 10920 -3770
rect -3040 -15750 10920 -3840
rect 11310 -3770 14070 -3750
rect 11310 -3840 11330 -3770
rect 11400 -3840 14070 -3770
rect 11310 -15750 14070 -3840
<< mimcapcontact >>
rect 11150 9270 11220 9340
rect 11150 8740 11220 8810
rect 11850 5260 11920 5330
rect 11850 4750 11920 4820
rect 7330 970 7410 1050
rect 8020 970 8100 1050
rect 8720 970 8800 1050
rect 9420 970 9500 1050
rect 10120 970 10200 1050
rect 10820 970 10900 1050
rect 11520 970 11600 1050
rect 12220 970 12300 1050
rect 12920 970 13000 1050
rect 13620 970 13700 1050
rect 7330 270 7410 350
rect 8020 270 8100 350
rect 8720 270 8800 350
rect 9420 270 9500 350
rect 10120 270 10200 350
rect 10820 270 10900 350
rect 11520 270 11600 350
rect 12220 270 12300 350
rect 12920 270 13000 350
rect 13620 270 13700 350
rect 7330 -430 7410 -350
rect 8020 -430 8100 -350
rect 8720 -430 8800 -350
rect 9420 -430 9500 -350
rect 10120 -430 10200 -350
rect 10820 -430 10900 -350
rect 11520 -430 11600 -350
rect 12220 -430 12300 -350
rect 12920 -430 13000 -350
rect 13620 -430 13700 -350
rect 7330 -1130 7410 -1050
rect 8020 -1130 8100 -1050
rect 8720 -1130 8800 -1050
rect 9420 -1130 9500 -1050
rect 10120 -1130 10200 -1050
rect 10820 -1130 10900 -1050
rect 11520 -1130 11600 -1050
rect 12220 -1130 12300 -1050
rect 12920 -1130 13000 -1050
rect 13620 -1130 13700 -1050
rect 7330 -1830 7410 -1750
rect 8020 -1830 8100 -1750
rect 8720 -1830 8800 -1750
rect 9420 -1830 9500 -1750
rect 10120 -1830 10200 -1750
rect 10820 -1830 10900 -1750
rect 11520 -1830 11600 -1750
rect 12220 -1830 12300 -1750
rect 12920 -1830 13000 -1750
rect 13620 -1830 13700 -1750
rect 7330 -2530 7410 -2450
rect 8020 -2530 8100 -2450
rect 8720 -2530 8800 -2450
rect 9420 -2530 9500 -2450
rect 10120 -2530 10200 -2450
rect 10820 -2530 10900 -2450
rect 11520 -2530 11600 -2450
rect 12220 -2530 12300 -2450
rect 12920 -2530 13000 -2450
rect 13620 -2530 13700 -2450
rect 10830 -3840 10900 -3770
rect 11330 -3840 11400 -3770
<< metal4 >>
rect 10750 9340 11240 9360
rect 10750 9270 10770 9340
rect 10840 9270 11150 9340
rect 11220 9270 11240 9340
rect 10750 9250 11240 9270
rect 10750 8810 11240 8830
rect 10750 8740 10770 8810
rect 10840 8740 11150 8810
rect 11220 8740 11240 8810
rect 10750 8720 11240 8740
rect 11450 5330 11930 5350
rect 11450 5260 11470 5330
rect 11540 5260 11850 5330
rect 11920 5260 11930 5330
rect 11450 5240 11930 5260
rect 11450 4820 11930 4840
rect 11450 4750 11470 4820
rect 11540 4750 11850 4820
rect 11920 4750 11930 4820
rect 11450 4730 11930 4750
rect 6790 1050 13710 1060
rect 6790 970 6800 1050
rect 6880 970 7330 1050
rect 7410 970 8020 1050
rect 8100 970 8720 1050
rect 8800 970 9420 1050
rect 9500 970 10120 1050
rect 10200 970 10820 1050
rect 10900 970 11520 1050
rect 11600 970 12220 1050
rect 12300 970 12920 1050
rect 13000 970 13620 1050
rect 13700 970 13710 1050
rect 6790 960 13710 970
rect 13610 360 13710 960
rect 7320 350 13710 360
rect 7320 270 7330 350
rect 7410 270 8020 350
rect 8100 270 8720 350
rect 8800 270 9420 350
rect 9500 270 10120 350
rect 10200 270 10820 350
rect 10900 270 11520 350
rect 11600 270 12220 350
rect 12300 270 12920 350
rect 13000 270 13620 350
rect 13700 270 13710 350
rect 7320 260 13710 270
rect 6790 -350 13710 -340
rect 6790 -430 6800 -350
rect 6880 -430 7330 -350
rect 7410 -430 8020 -350
rect 8100 -430 8720 -350
rect 8800 -430 9420 -350
rect 9500 -430 10120 -350
rect 10200 -430 10820 -350
rect 10900 -430 11520 -350
rect 11600 -430 12220 -350
rect 12300 -430 12920 -350
rect 13000 -430 13620 -350
rect 13700 -430 13710 -350
rect 6790 -440 13710 -430
rect 13610 -1040 13710 -440
rect 7320 -1050 13710 -1040
rect 7320 -1130 7330 -1050
rect 7410 -1130 8020 -1050
rect 8100 -1130 8720 -1050
rect 8800 -1130 9420 -1050
rect 9500 -1130 10120 -1050
rect 10200 -1130 10820 -1050
rect 10900 -1130 11520 -1050
rect 11600 -1130 12220 -1050
rect 12300 -1130 12920 -1050
rect 13000 -1130 13620 -1050
rect 13700 -1130 13710 -1050
rect 7320 -1140 13710 -1130
rect 6650 -1750 13710 -1740
rect 6650 -1830 6660 -1750
rect 6740 -1830 7330 -1750
rect 7410 -1830 8020 -1750
rect 8100 -1830 8720 -1750
rect 8800 -1830 9420 -1750
rect 9500 -1830 10120 -1750
rect 10200 -1830 10820 -1750
rect 10900 -1830 11520 -1750
rect 11600 -1830 12220 -1750
rect 12300 -1830 12920 -1750
rect 13000 -1830 13620 -1750
rect 13700 -1830 13710 -1750
rect 6650 -1840 13710 -1830
rect 13610 -2440 13710 -1840
rect 7320 -2450 13710 -2440
rect 7320 -2530 7330 -2450
rect 7410 -2530 8020 -2450
rect 8100 -2530 8720 -2450
rect 8800 -2530 9420 -2450
rect 9500 -2530 10120 -2450
rect 10200 -2530 10820 -2450
rect 10900 -2530 11520 -2450
rect 11600 -2530 12220 -2450
rect 12300 -2530 12920 -2450
rect 13000 -2530 13620 -2450
rect 13700 -2530 13710 -2450
rect 7320 -2540 13710 -2530
rect 10810 -3390 10920 -3370
rect 10810 -3460 10830 -3390
rect 10900 -3460 10920 -3390
rect 10810 -3770 10920 -3460
rect 10810 -3840 10830 -3770
rect 10900 -3840 10920 -3770
rect 10810 -3850 10920 -3840
rect 11310 -3390 11420 -3370
rect 11310 -3460 11330 -3390
rect 11400 -3460 11420 -3390
rect 11310 -3770 11420 -3460
rect 11310 -3840 11330 -3770
rect 11400 -3840 11420 -3770
rect 11310 -3850 11420 -3840
<< end >>
