magic
tech sky130A
timestamp 1756512595
<< via1 >>
rect 13280 10055 13310 10085
<< metal2 >>
rect 11685 16840 11725 16845
rect 11685 16811 11690 16840
rect 11720 16811 11725 16840
rect 11685 16799 11725 16811
rect 11685 16770 11690 16799
rect 11720 16770 11725 16799
rect 11685 16765 11725 16770
rect 13275 10085 13315 10090
rect 13275 10055 13280 10085
rect 13310 10055 13315 10085
rect 13275 9765 13315 10055
rect 13255 9755 13335 9765
rect 13255 9725 13280 9755
rect 13310 9725 13335 9755
rect 13255 9715 13335 9725
<< via2 >>
rect 11690 16811 11720 16840
rect 11690 16770 11720 16799
rect 13280 9725 13310 9755
<< metal3 >>
rect 100 18210 11505 18215
rect 100 18170 105 18210
rect 145 18170 155 18210
rect 195 18170 205 18210
rect 245 18170 255 18210
rect 295 18170 11460 18210
rect 11500 18170 11505 18210
rect 100 18160 11505 18170
rect 100 18120 105 18160
rect 145 18120 155 18160
rect 195 18120 205 18160
rect 245 18120 255 18160
rect 295 18120 11460 18160
rect 11500 18120 11505 18160
rect 100 18110 11505 18120
rect 100 18070 105 18110
rect 145 18070 155 18110
rect 195 18070 205 18110
rect 245 18070 255 18110
rect 295 18070 11460 18110
rect 11500 18070 11505 18110
rect 100 18060 11505 18070
rect 100 18020 105 18060
rect 145 18020 155 18060
rect 195 18020 205 18060
rect 245 18020 255 18060
rect 295 18020 11460 18060
rect 11500 18020 11505 18060
rect 100 18015 11505 18020
rect 400 17795 12090 17800
rect 400 17755 405 17795
rect 445 17755 455 17795
rect 495 17755 505 17795
rect 545 17755 555 17795
rect 595 17755 12045 17795
rect 12085 17755 12090 17795
rect 400 17745 12090 17755
rect 400 17705 405 17745
rect 445 17705 455 17745
rect 495 17705 505 17745
rect 545 17705 555 17745
rect 595 17705 12045 17745
rect 12085 17705 12090 17745
rect 400 17695 12090 17705
rect 400 17655 405 17695
rect 445 17655 455 17695
rect 495 17655 505 17695
rect 545 17655 555 17695
rect 595 17655 12045 17695
rect 12085 17655 12090 17695
rect 400 17645 12090 17655
rect 400 17605 405 17645
rect 445 17605 455 17645
rect 495 17605 505 17645
rect 545 17605 555 17645
rect 595 17605 12045 17645
rect 12085 17605 12090 17645
rect 400 17600 12090 17605
rect 11685 16840 15265 16845
rect 11685 16811 11690 16840
rect 11720 16825 15265 16840
rect 11720 16811 15205 16825
rect 11685 16799 15205 16811
rect 11685 16770 11690 16799
rect 11720 16785 15205 16799
rect 15245 16785 15265 16825
rect 11720 16770 15265 16785
rect 11685 16765 15265 16770
rect 13255 9760 13335 9765
rect 13255 9720 13275 9760
rect 13315 9720 13335 9760
rect 13255 9715 13335 9720
<< via3 >>
rect 105 18170 145 18210
rect 155 18170 195 18210
rect 205 18170 245 18210
rect 255 18170 295 18210
rect 11460 18170 11500 18210
rect 105 18120 145 18160
rect 155 18120 195 18160
rect 205 18120 245 18160
rect 255 18120 295 18160
rect 11460 18120 11500 18160
rect 105 18070 145 18110
rect 155 18070 195 18110
rect 205 18070 245 18110
rect 255 18070 295 18110
rect 11460 18070 11500 18110
rect 105 18020 145 18060
rect 155 18020 195 18060
rect 205 18020 245 18060
rect 255 18020 295 18060
rect 11460 18020 11500 18060
rect 405 17755 445 17795
rect 455 17755 495 17795
rect 505 17755 545 17795
rect 555 17755 595 17795
rect 12045 17755 12085 17795
rect 405 17705 445 17745
rect 455 17705 495 17745
rect 505 17705 545 17745
rect 555 17705 595 17745
rect 12045 17705 12085 17745
rect 405 17655 445 17695
rect 455 17655 495 17695
rect 505 17655 545 17695
rect 555 17655 595 17695
rect 12045 17655 12085 17695
rect 405 17605 445 17645
rect 455 17605 495 17645
rect 505 17605 545 17645
rect 555 17605 595 17645
rect 12045 17605 12085 17645
rect 15205 16785 15245 16825
rect 13275 9755 13315 9760
rect 13275 9725 13280 9755
rect 13280 9725 13310 9755
rect 13310 9725 13315 9755
rect 13275 9720 13315 9725
<< metal4 >>
rect 3067 22476 3097 22576
rect 3343 22476 3373 22576
rect 3619 22476 3649 22576
rect 3895 22476 3925 22576
rect 4171 22476 4201 22576
rect 4447 22476 4477 22576
rect 4723 22476 4753 22576
rect 4999 22476 5029 22576
rect 5275 22476 5305 22576
rect 5551 22476 5581 22576
rect 5827 22476 5857 22576
rect 6103 22476 6133 22576
rect 6379 22476 6409 22576
rect 6655 22476 6685 22576
rect 6931 22476 6961 22576
rect 7207 22476 7237 22576
rect 7483 22476 7513 22576
rect 7759 22476 7789 22576
rect 8035 22476 8065 22576
rect 8311 22476 8341 22576
rect 8587 22476 8617 22576
rect 8863 22476 8893 22576
rect 9139 22476 9169 22576
rect 9415 22476 9445 22576
rect 9691 22476 9721 22576
rect 9967 22476 9997 22576
rect 10243 22476 10273 22576
rect 10519 22476 10549 22576
rect 10795 22476 10825 22576
rect 11071 22476 11101 22576
rect 11347 22476 11377 22576
rect 11623 22476 11653 22576
rect 11899 22476 11929 22576
rect 12175 22476 12205 22576
rect 12451 22476 12481 22576
rect 12727 22476 12757 22576
rect 13003 22476 13033 22576
rect 13279 22476 13309 22576
rect 13555 22476 13585 22576
rect 13831 22476 13861 22576
rect 14107 22476 14137 22576
rect 14383 22476 14413 22576
rect 14659 22476 14689 22576
rect 100 18210 300 22076
rect 100 18170 105 18210
rect 145 18170 155 18210
rect 195 18170 205 18210
rect 245 18170 255 18210
rect 295 18170 300 18210
rect 100 18160 300 18170
rect 100 18120 105 18160
rect 145 18120 155 18160
rect 195 18120 205 18160
rect 245 18120 255 18160
rect 295 18120 300 18160
rect 100 18110 300 18120
rect 100 18070 105 18110
rect 145 18070 155 18110
rect 195 18070 205 18110
rect 245 18070 255 18110
rect 295 18070 300 18110
rect 100 18060 300 18070
rect 100 18020 105 18060
rect 145 18020 155 18060
rect 195 18020 205 18060
rect 245 18020 255 18060
rect 295 18020 300 18060
rect 100 500 300 18020
rect 400 17795 600 22076
rect 400 17755 405 17795
rect 445 17755 455 17795
rect 495 17755 505 17795
rect 545 17755 555 17795
rect 595 17755 600 17795
rect 400 17745 600 17755
rect 400 17705 405 17745
rect 445 17705 455 17745
rect 495 17705 505 17745
rect 545 17705 555 17745
rect 595 17705 600 17745
rect 400 17695 600 17705
rect 400 17655 405 17695
rect 445 17655 455 17695
rect 495 17655 505 17695
rect 545 17655 555 17695
rect 595 17655 600 17695
rect 400 17645 600 17655
rect 400 17605 405 17645
rect 445 17605 455 17645
rect 495 17605 505 17645
rect 545 17605 555 17645
rect 595 17605 600 17645
rect 400 500 600 17605
rect 11455 18210 11505 18215
rect 11455 18170 11460 18210
rect 11500 18170 11505 18210
rect 11455 18160 11505 18170
rect 11455 18120 11460 18160
rect 11500 18120 11505 18160
rect 11455 18110 11505 18120
rect 11455 18070 11460 18110
rect 11500 18070 11505 18110
rect 11455 18060 11505 18070
rect 11455 18020 11460 18060
rect 11500 18020 11505 18060
rect 11455 16260 11505 18020
rect 12040 17795 12090 17800
rect 12040 17755 12045 17795
rect 12085 17755 12090 17795
rect 12040 17745 12090 17755
rect 12040 17705 12045 17745
rect 12085 17705 12090 17745
rect 12040 17695 12090 17705
rect 12040 17655 12045 17695
rect 12085 17655 12090 17695
rect 12040 17645 12090 17655
rect 12040 17605 12045 17645
rect 12085 17605 12090 17645
rect 12040 16410 12090 17605
rect 15185 16825 15265 16845
rect 15185 16785 15205 16825
rect 15245 16785 15265 16825
rect 13255 9760 13335 9765
rect 13255 9720 13275 9760
rect 13315 9720 13335 9760
rect 13255 100 13335 9720
rect 15185 100 15265 16785
rect 1657 0 1747 100
rect 3589 0 3679 100
rect 5521 0 5611 100
rect 7453 0 7543 100
rect 9385 0 9475 100
rect 11317 0 11407 100
rect 13249 0 13339 100
rect 15181 0 15271 100
use pll_bgr_magic_flat  pll_bgr_magic_flat_0
timestamp 1756511854
transform 0 -1 13930 -1 0 17120
box 0 0 15790 7605
<< labels >>
flabel metal4 s 14383 22476 14413 22576 0 FreeSans 240 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 14659 22476 14689 22576 0 FreeSans 240 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 14107 22476 14137 22576 0 FreeSans 240 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 15181 0 15271 100 0 FreeSans 480 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 13249 0 13339 100 0 FreeSans 480 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 11317 0 11407 100 0 FreeSans 480 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 9385 0 9475 100 0 FreeSans 480 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 7453 0 7543 100 0 FreeSans 480 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 5521 0 5611 100 0 FreeSans 480 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 3589 0 3679 100 0 FreeSans 480 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 1657 0 1747 100 0 FreeSans 480 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 13831 22476 13861 22576 0 FreeSans 240 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 13555 22476 13585 22576 0 FreeSans 240 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 13279 22476 13309 22576 0 FreeSans 240 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 13003 22476 13033 22576 0 FreeSans 240 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 12727 22476 12757 22576 0 FreeSans 240 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 12451 22476 12481 22576 0 FreeSans 240 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 12175 22476 12205 22576 0 FreeSans 240 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 11899 22476 11929 22576 0 FreeSans 240 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 11623 22476 11653 22576 0 FreeSans 240 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 11347 22476 11377 22576 0 FreeSans 240 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 11071 22476 11101 22576 0 FreeSans 240 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 10795 22476 10825 22576 0 FreeSans 240 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 10519 22476 10549 22576 0 FreeSans 240 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 10243 22476 10273 22576 0 FreeSans 240 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 9967 22476 9997 22576 0 FreeSans 240 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 9691 22476 9721 22576 0 FreeSans 240 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 4999 22476 5029 22576 0 FreeSans 240 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 4723 22476 4753 22576 0 FreeSans 240 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4447 22476 4477 22576 0 FreeSans 240 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 4171 22476 4201 22576 0 FreeSans 240 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3895 22476 3925 22576 0 FreeSans 240 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 3619 22476 3649 22576 0 FreeSans 240 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3343 22476 3373 22576 0 FreeSans 240 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3067 22476 3097 22576 0 FreeSans 240 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 7207 22476 7237 22576 0 FreeSans 240 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 6931 22476 6961 22576 0 FreeSans 240 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 6655 22476 6685 22576 0 FreeSans 240 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 6379 22476 6409 22576 0 FreeSans 240 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 6103 22476 6133 22576 0 FreeSans 240 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 5827 22476 5857 22576 0 FreeSans 240 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 5551 22476 5581 22576 0 FreeSans 240 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 5275 22476 5305 22576 0 FreeSans 240 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 9415 22476 9445 22576 0 FreeSans 240 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 9139 22476 9169 22576 0 FreeSans 240 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 8863 22476 8893 22576 0 FreeSans 240 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 8587 22476 8617 22576 0 FreeSans 240 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 8311 22476 8341 22576 0 FreeSans 240 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 8035 22476 8065 22576 0 FreeSans 240 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 7759 22476 7789 22576 0 FreeSans 240 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 7483 22476 7513 22576 0 FreeSans 240 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 100 500 300 22076 1 FreeSans 200 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 400 500 600 22076 1 FreeSans 200 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16100 22576
<< end >>
